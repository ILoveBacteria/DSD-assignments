module NeuralNetwork (
    input clk,
    input rst,
    input start,
    input [783:0] in_features, // 784 input features
    output reg [3:0] prediction, // 10 output classes (ArgMax index)
    output reg done
);

    // register to hold the input features
    reg [783:0] features;

    // state machine
    localparam IDLE = 0, COMPUTE = 1;
    reg state;
    reg [2:0] count_clocks; 

    // Define the parameters for layer sizes
    parameter INPUT_SIZE = 784;
    parameter HIDDEN1_SIZE = 64;
    parameter HIDDEN2_SIZE = 32;
    parameter OUTPUT_SIZE = 10;
    
    // Define memory for weights and biases (assumed preloaded)
    wire signed [15:0] weights1 [0:HIDDEN1_SIZE-1][0:INPUT_SIZE-1];
    wire signed [15:0] biases1 [0:HIDDEN1_SIZE-1];
    
    wire signed [15:0] weights2 [0:HIDDEN2_SIZE-1][0:HIDDEN1_SIZE-1];
    wire signed [15:0] biases2 [0:HIDDEN2_SIZE-1];
    
    wire signed [15:0] weights3 [0:OUTPUT_SIZE-1][0:HIDDEN2_SIZE-1];
    wire signed [15:0] biases3 [0:OUTPUT_SIZE-1];
    
    // Layer Outputs
    reg signed [15:0] hidden1 [0:HIDDEN1_SIZE-1];
    reg signed [15:0] hidden2 [0:HIDDEN2_SIZE-1];
    reg signed [15:0] output_layer [0:OUTPUT_SIZE-1];
    
    integer i, j;
    
    // ReLU activation function
    function signed [15:0] relu;
        input signed [15:0] x;
        begin
            relu = (x > 0) ? x : 0;
        end
    endfunction


    // ============================================
    // combinational Computation of the neurons
    // ============================================

    // layer 1
    reg signed [15:0] new_hidden1 [0:HIDDEN1_SIZE-1];
    always @(*) begin
        for (i = 0; i < HIDDEN1_SIZE; i = i + 1) begin
            new_hidden1[i] = biases1[i];
            for (j = 0; j < INPUT_SIZE; j = j + 1) begin
                new_hidden1[i] = new_hidden1[i] + (features[j] == 1 ? weights1[i][j] : 0); 
            end
            new_hidden1[i] = relu(new_hidden1[i]); 
        end
    end

    // layer 2
    reg signed [15:0] new_hidden2 [0:HIDDEN2_SIZE-1];
    reg signed [15:0] multiplier_out2 [0:HIDDEN2_SIZE-1][0:HIDDEN1_SIZE-1];
    reg signed [15:0] shift_out2 [0:HIDDEN2_SIZE-1][0:HIDDEN1_SIZE-1];
    always @(*) begin
        for (i = 0; i < HIDDEN2_SIZE; i = i + 1) begin
            new_hidden2[i] = biases2[i];
            for (j = 0; j < HIDDEN1_SIZE; j = j + 1) begin
                multiplier_out2[i][j] = hidden1[j] * weights2[i][j];
                shift_out2[i][j] = multiplier_out2[i][j] >> 8;
                new_hidden2[i] = new_hidden2[i] + shift_out2[i][j];
            end
            new_hidden2[i] = relu(new_hidden2[i]);
        end
    end

    // Output Layer computation
    reg signed [15:0] new_output_layer [0:OUTPUT_SIZE-1];
    reg signed [15:0] multiplier_out3 [0:OUTPUT_SIZE-1][0:HIDDEN2_SIZE-1];
    reg signed [15:0] shift_out3 [0:OUTPUT_SIZE-1][0:HIDDEN2_SIZE-1];
    always @(*) begin
        for (i = 0; i < OUTPUT_SIZE; i = i + 1) begin
            new_output_layer[i] = biases3[i];
            for (j = 0; j < HIDDEN2_SIZE; j = j + 1) begin
                multiplier_out3[i][j] = hidden2[j] * weights3[i][j];
                shift_out3[i][j] = multiplier_out3[i][j] >> 8;
                new_output_layer[i] = new_output_layer[i] + shift_out3[i][j];
            end
        end
    end

    // ArgMax operation
    reg [3:0] new_prediction;
    always @(*) begin
        new_prediction = 0;
        for (i = 1; i < OUTPUT_SIZE; i = i + 1) begin
            if (output_layer[i] > output_layer[new_prediction]) begin
                new_prediction = i;
            end
        end
    end
    

    // ============================================
    // Sequential update of the neurons
    // ============================================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            done <= 0;
            count_clocks <= 0;
            prediction <= 0;
            for (i = 0; i < INPUT_SIZE; i = i + 1) begin
                features[i] <= 0;
            end
        end 
        else if (state == IDLE) begin
            if (start) begin
                // Load the input features
                for (i = 0; i < INPUT_SIZE; i = i + 1) begin
                    features[i] <= in_features[i];
                end
                state <= COMPUTE;
                done <= 0;
                count_clocks <= 0;
            end
        end 
        else begin
            // Layer 1 computation
            for (i = 0; i < HIDDEN1_SIZE; i = i + 1) begin
                hidden1[i] <= new_hidden1[i];
            end

            // Layer 2 computation
            for (i = 0; i < HIDDEN2_SIZE; i = i + 1) begin
                hidden2[i] <= new_hidden2[i];
            end

            // Output Layer computation
            for (i = 0; i < OUTPUT_SIZE; i = i + 1) begin
                output_layer[i] <= new_output_layer[i];
            end

            // ArgMax operation
            prediction <= new_prediction;

            // Update state or increment the clock counter
            if (count_clocks >= 3) begin
                state <= IDLE;
                done <= 1;
            end
            else begin
                count_clocks <= count_clocks + 1;
            end
        end
    end

    // ============================================
    // Initialize the weights and biases
    // ============================================
    assign weights1[0][0] = 16'b0000000000000000;
    assign weights1[0][1] = 16'b0000000000000000;
    assign weights1[0][2] = 16'b0000000000000000;
    assign weights1[0][3] = 16'b0000000000000000;
    assign weights1[0][4] = 16'b0000000000001100;
    assign weights1[0][5] = 16'b0000000000011010;
    assign weights1[0][6] = 16'b0000000000100111;
    assign weights1[0][7] = 16'b0000000000101010;
    assign weights1[0][8] = 16'b0000000000111110;
    assign weights1[0][9] = 16'b0000000001001001;
    assign weights1[0][10] = 16'b0000000000111111;
    assign weights1[0][11] = 16'b0000000001000001;
    assign weights1[0][12] = 16'b0000000000110011;
    assign weights1[0][13] = 16'b0000000000100101;
    assign weights1[0][14] = 16'b0000000000100000;
    assign weights1[0][15] = 16'b0000000000011110;
    assign weights1[0][16] = 16'b0000000000000110;
    assign weights1[0][17] = 16'b0000000000000101;
    assign weights1[0][18] = 16'b0000000000011001;
    assign weights1[0][19] = 16'b1111111111110101;
    assign weights1[0][20] = 16'b0000000000000011;
    assign weights1[0][21] = 16'b0000000000000011;
    assign weights1[0][22] = 16'b0000000000001111;
    assign weights1[0][23] = 16'b1111111111110101;
    assign weights1[0][24] = 16'b1111111111101011;
    assign weights1[0][25] = 16'b1111111111101100;
    assign weights1[0][26] = 16'b1111111111110100;
    assign weights1[0][27] = 16'b1111111111111010;
    assign weights1[0][28] = 16'b0000000000000000;
    assign weights1[0][29] = 16'b0000000000000000;
    assign weights1[0][30] = 16'b0000000000000000;
    assign weights1[0][31] = 16'b0000000000001010;
    assign weights1[0][32] = 16'b0000000000010101;
    assign weights1[0][33] = 16'b0000000000100100;
    assign weights1[0][34] = 16'b0000000000101010;
    assign weights1[0][35] = 16'b0000000001000010;
    assign weights1[0][36] = 16'b0000000001010011;
    assign weights1[0][37] = 16'b0000000001000111;
    assign weights1[0][38] = 16'b0000000001010010;
    assign weights1[0][39] = 16'b0000000001011010;
    assign weights1[0][40] = 16'b0000000001001000;
    assign weights1[0][41] = 16'b0000000000101000;
    assign weights1[0][42] = 16'b0000000000100111;
    assign weights1[0][43] = 16'b0000000000011010;
    assign weights1[0][44] = 16'b0000000000011110;
    assign weights1[0][45] = 16'b0000000000011100;
    assign weights1[0][46] = 16'b0000000000000010;
    assign weights1[0][47] = 16'b0000000000000110;
    assign weights1[0][48] = 16'b1111111111110111;
    assign weights1[0][49] = 16'b0000000000010000;
    assign weights1[0][50] = 16'b0000000000001010;
    assign weights1[0][51] = 16'b0000000000000110;
    assign weights1[0][52] = 16'b1111111111111001;
    assign weights1[0][53] = 16'b1111111111111010;
    assign weights1[0][54] = 16'b1111111111110000;
    assign weights1[0][55] = 16'b1111111111101110;
    assign weights1[0][56] = 16'b0000000000000000;
    assign weights1[0][57] = 16'b0000000000000000;
    assign weights1[0][58] = 16'b0000000000000111;
    assign weights1[0][59] = 16'b0000000000001110;
    assign weights1[0][60] = 16'b0000000000011000;
    assign weights1[0][61] = 16'b0000000000011101;
    assign weights1[0][62] = 16'b0000000000100100;
    assign weights1[0][63] = 16'b0000000000110001;
    assign weights1[0][64] = 16'b0000000000111101;
    assign weights1[0][65] = 16'b0000000001000101;
    assign weights1[0][66] = 16'b0000000001001001;
    assign weights1[0][67] = 16'b0000000001000110;
    assign weights1[0][68] = 16'b0000000001001101;
    assign weights1[0][69] = 16'b0000000001000010;
    assign weights1[0][70] = 16'b0000000000101111;
    assign weights1[0][71] = 16'b0000000000011111;
    assign weights1[0][72] = 16'b0000000000101100;
    assign weights1[0][73] = 16'b0000000000100100;
    assign weights1[0][74] = 16'b0000000000001111;
    assign weights1[0][75] = 16'b0000000000001000;
    assign weights1[0][76] = 16'b0000000000010000;
    assign weights1[0][77] = 16'b0000000000011110;
    assign weights1[0][78] = 16'b0000000000000100;
    assign weights1[0][79] = 16'b0000000000000110;
    assign weights1[0][80] = 16'b0000000000001111;
    assign weights1[0][81] = 16'b1111111111110010;
    assign weights1[0][82] = 16'b1111111111110110;
    assign weights1[0][83] = 16'b1111111111110010;
    assign weights1[0][84] = 16'b0000000000000000;
    assign weights1[0][85] = 16'b0000000000000011;
    assign weights1[0][86] = 16'b0000000000001001;
    assign weights1[0][87] = 16'b0000000000010000;
    assign weights1[0][88] = 16'b0000000000011000;
    assign weights1[0][89] = 16'b0000000000010111;
    assign weights1[0][90] = 16'b0000000000010111;
    assign weights1[0][91] = 16'b0000000000101100;
    assign weights1[0][92] = 16'b0000000000110001;
    assign weights1[0][93] = 16'b0000000000111101;
    assign weights1[0][94] = 16'b0000000000111111;
    assign weights1[0][95] = 16'b0000000001000101;
    assign weights1[0][96] = 16'b0000000001010111;
    assign weights1[0][97] = 16'b0000000001010101;
    assign weights1[0][98] = 16'b0000000001001001;
    assign weights1[0][99] = 16'b0000000000110110;
    assign weights1[0][100] = 16'b0000000000010010;
    assign weights1[0][101] = 16'b0000000000101000;
    assign weights1[0][102] = 16'b0000000000011111;
    assign weights1[0][103] = 16'b0000000000011110;
    assign weights1[0][104] = 16'b0000000000010100;
    assign weights1[0][105] = 16'b0000000000010000;
    assign weights1[0][106] = 16'b0000000000011001;
    assign weights1[0][107] = 16'b0000000000001001;
    assign weights1[0][108] = 16'b0000000000000110;
    assign weights1[0][109] = 16'b0000000000000100;
    assign weights1[0][110] = 16'b1111111111111000;
    assign weights1[0][111] = 16'b1111111111101010;
    assign weights1[0][112] = 16'b0000000000000011;
    assign weights1[0][113] = 16'b0000000000000101;
    assign weights1[0][114] = 16'b1111111111111101;
    assign weights1[0][115] = 16'b1111111111110111;
    assign weights1[0][116] = 16'b1111111111110100;
    assign weights1[0][117] = 16'b1111111111110100;
    assign weights1[0][118] = 16'b1111111111111101;
    assign weights1[0][119] = 16'b0000000000000111;
    assign weights1[0][120] = 16'b0000000000100010;
    assign weights1[0][121] = 16'b0000000000011101;
    assign weights1[0][122] = 16'b0000000000101010;
    assign weights1[0][123] = 16'b0000000001000011;
    assign weights1[0][124] = 16'b0000000000110111;
    assign weights1[0][125] = 16'b0000000001100100;
    assign weights1[0][126] = 16'b0000000001100000;
    assign weights1[0][127] = 16'b0000000001001000;
    assign weights1[0][128] = 16'b0000000000110101;
    assign weights1[0][129] = 16'b0000000000100110;
    assign weights1[0][130] = 16'b0000000000011101;
    assign weights1[0][131] = 16'b0000000000010110;
    assign weights1[0][132] = 16'b0000000000010101;
    assign weights1[0][133] = 16'b0000000000001110;
    assign weights1[0][134] = 16'b0000000000010001;
    assign weights1[0][135] = 16'b0000000000010001;
    assign weights1[0][136] = 16'b0000000000001001;
    assign weights1[0][137] = 16'b0000000000000100;
    assign weights1[0][138] = 16'b0000000000001011;
    assign weights1[0][139] = 16'b1111111111110111;
    assign weights1[0][140] = 16'b1111111111111110;
    assign weights1[0][141] = 16'b1111111111110011;
    assign weights1[0][142] = 16'b1111111111101111;
    assign weights1[0][143] = 16'b1111111111100000;
    assign weights1[0][144] = 16'b1111111111010010;
    assign weights1[0][145] = 16'b1111111111001110;
    assign weights1[0][146] = 16'b1111111111010011;
    assign weights1[0][147] = 16'b1111111111100001;
    assign weights1[0][148] = 16'b1111111111010101;
    assign weights1[0][149] = 16'b1111111111001011;
    assign weights1[0][150] = 16'b1111111111101000;
    assign weights1[0][151] = 16'b1111111111101011;
    assign weights1[0][152] = 16'b0000000000010001;
    assign weights1[0][153] = 16'b0000000000110111;
    assign weights1[0][154] = 16'b0000000001000111;
    assign weights1[0][155] = 16'b0000000001010110;
    assign weights1[0][156] = 16'b0000000001010001;
    assign weights1[0][157] = 16'b0000000001000100;
    assign weights1[0][158] = 16'b0000000000100011;
    assign weights1[0][159] = 16'b0000000000010011;
    assign weights1[0][160] = 16'b0000000000101100;
    assign weights1[0][161] = 16'b0000000000100010;
    assign weights1[0][162] = 16'b0000000000011100;
    assign weights1[0][163] = 16'b0000000000011011;
    assign weights1[0][164] = 16'b0000000000010010;
    assign weights1[0][165] = 16'b0000000000010001;
    assign weights1[0][166] = 16'b0000000000010010;
    assign weights1[0][167] = 16'b1111111111111101;
    assign weights1[0][168] = 16'b1111111111111000;
    assign weights1[0][169] = 16'b1111111111100110;
    assign weights1[0][170] = 16'b1111111111001101;
    assign weights1[0][171] = 16'b1111111110111011;
    assign weights1[0][172] = 16'b1111111110100110;
    assign weights1[0][173] = 16'b1111111110011111;
    assign weights1[0][174] = 16'b1111111110100100;
    assign weights1[0][175] = 16'b1111111110101001;
    assign weights1[0][176] = 16'b1111111110011100;
    assign weights1[0][177] = 16'b1111111110011100;
    assign weights1[0][178] = 16'b1111111110011011;
    assign weights1[0][179] = 16'b1111111110111111;
    assign weights1[0][180] = 16'b1111111110100111;
    assign weights1[0][181] = 16'b1111111111000111;
    assign weights1[0][182] = 16'b1111111111101011;
    assign weights1[0][183] = 16'b0000000000100111;
    assign weights1[0][184] = 16'b0000000000111101;
    assign weights1[0][185] = 16'b0000000001000101;
    assign weights1[0][186] = 16'b0000000000101111;
    assign weights1[0][187] = 16'b0000000000101010;
    assign weights1[0][188] = 16'b0000000000011100;
    assign weights1[0][189] = 16'b0000000000010110;
    assign weights1[0][190] = 16'b0000000000100100;
    assign weights1[0][191] = 16'b0000000000001001;
    assign weights1[0][192] = 16'b0000000000010110;
    assign weights1[0][193] = 16'b0000000000011101;
    assign weights1[0][194] = 16'b0000000000001011;
    assign weights1[0][195] = 16'b0000000000001110;
    assign weights1[0][196] = 16'b1111111111110110;
    assign weights1[0][197] = 16'b1111111111001110;
    assign weights1[0][198] = 16'b1111111110110101;
    assign weights1[0][199] = 16'b1111111110011010;
    assign weights1[0][200] = 16'b1111111101110101;
    assign weights1[0][201] = 16'b1111111101110010;
    assign weights1[0][202] = 16'b1111111110000001;
    assign weights1[0][203] = 16'b1111111110000011;
    assign weights1[0][204] = 16'b1111111101101011;
    assign weights1[0][205] = 16'b1111111101110101;
    assign weights1[0][206] = 16'b1111111101101110;
    assign weights1[0][207] = 16'b1111111110010001;
    assign weights1[0][208] = 16'b1111111110001010;
    assign weights1[0][209] = 16'b1111111110001111;
    assign weights1[0][210] = 16'b1111111110100011;
    assign weights1[0][211] = 16'b1111111111001001;
    assign weights1[0][212] = 16'b1111111111111110;
    assign weights1[0][213] = 16'b0000000000101100;
    assign weights1[0][214] = 16'b0000000000101111;
    assign weights1[0][215] = 16'b0000000000101100;
    assign weights1[0][216] = 16'b0000000000101010;
    assign weights1[0][217] = 16'b0000000000101110;
    assign weights1[0][218] = 16'b0000000000100000;
    assign weights1[0][219] = 16'b0000000000100111;
    assign weights1[0][220] = 16'b0000000000101011;
    assign weights1[0][221] = 16'b0000000000010110;
    assign weights1[0][222] = 16'b0000000000001001;
    assign weights1[0][223] = 16'b0000000000010101;
    assign weights1[0][224] = 16'b1111111111101001;
    assign weights1[0][225] = 16'b1111111111000010;
    assign weights1[0][226] = 16'b1111111110100101;
    assign weights1[0][227] = 16'b1111111110010100;
    assign weights1[0][228] = 16'b1111111101111001;
    assign weights1[0][229] = 16'b1111111101110111;
    assign weights1[0][230] = 16'b1111111101111100;
    assign weights1[0][231] = 16'b1111111110001101;
    assign weights1[0][232] = 16'b1111111101111111;
    assign weights1[0][233] = 16'b1111111110000110;
    assign weights1[0][234] = 16'b1111111110110010;
    assign weights1[0][235] = 16'b1111111110101101;
    assign weights1[0][236] = 16'b1111111111001010;
    assign weights1[0][237] = 16'b1111111110111001;
    assign weights1[0][238] = 16'b1111111111001001;
    assign weights1[0][239] = 16'b1111111110111011;
    assign weights1[0][240] = 16'b1111111111001101;
    assign weights1[0][241] = 16'b1111111111111110;
    assign weights1[0][242] = 16'b0000000000011001;
    assign weights1[0][243] = 16'b0000000000101111;
    assign weights1[0][244] = 16'b0000000000000011;
    assign weights1[0][245] = 16'b0000000000110010;
    assign weights1[0][246] = 16'b0000000000010110;
    assign weights1[0][247] = 16'b0000000000011010;
    assign weights1[0][248] = 16'b0000000000010100;
    assign weights1[0][249] = 16'b0000000000000011;
    assign weights1[0][250] = 16'b0000000000100000;
    assign weights1[0][251] = 16'b0000000000001111;
    assign weights1[0][252] = 16'b1111111111101000;
    assign weights1[0][253] = 16'b1111111111000111;
    assign weights1[0][254] = 16'b1111111110101101;
    assign weights1[0][255] = 16'b1111111110011111;
    assign weights1[0][256] = 16'b1111111110100010;
    assign weights1[0][257] = 16'b1111111110100000;
    assign weights1[0][258] = 16'b1111111110110010;
    assign weights1[0][259] = 16'b1111111110110011;
    assign weights1[0][260] = 16'b1111111110100101;
    assign weights1[0][261] = 16'b1111111111100101;
    assign weights1[0][262] = 16'b1111111111011010;
    assign weights1[0][263] = 16'b1111111111101110;
    assign weights1[0][264] = 16'b1111111111101000;
    assign weights1[0][265] = 16'b1111111111100011;
    assign weights1[0][266] = 16'b1111111111001011;
    assign weights1[0][267] = 16'b1111111111001000;
    assign weights1[0][268] = 16'b1111111111001101;
    assign weights1[0][269] = 16'b1111111111100100;
    assign weights1[0][270] = 16'b1111111111101010;
    assign weights1[0][271] = 16'b0000000000000010;
    assign weights1[0][272] = 16'b0000000000000001;
    assign weights1[0][273] = 16'b0000000000011001;
    assign weights1[0][274] = 16'b0000000000100100;
    assign weights1[0][275] = 16'b0000000000011101;
    assign weights1[0][276] = 16'b0000000000010000;
    assign weights1[0][277] = 16'b0000000000010001;
    assign weights1[0][278] = 16'b0000000000010100;
    assign weights1[0][279] = 16'b0000000000010010;
    assign weights1[0][280] = 16'b1111111111111100;
    assign weights1[0][281] = 16'b1111111111101010;
    assign weights1[0][282] = 16'b1111111111011001;
    assign weights1[0][283] = 16'b1111111111100010;
    assign weights1[0][284] = 16'b1111111111110000;
    assign weights1[0][285] = 16'b0000000000000010;
    assign weights1[0][286] = 16'b0000000000000101;
    assign weights1[0][287] = 16'b0000000000000000;
    assign weights1[0][288] = 16'b0000000000010010;
    assign weights1[0][289] = 16'b0000000000011001;
    assign weights1[0][290] = 16'b1111111111111101;
    assign weights1[0][291] = 16'b1111111111101111;
    assign weights1[0][292] = 16'b1111111111110011;
    assign weights1[0][293] = 16'b1111111111101111;
    assign weights1[0][294] = 16'b1111111111100110;
    assign weights1[0][295] = 16'b1111111111110001;
    assign weights1[0][296] = 16'b1111111111011010;
    assign weights1[0][297] = 16'b1111111111011101;
    assign weights1[0][298] = 16'b1111111111011101;
    assign weights1[0][299] = 16'b1111111111100111;
    assign weights1[0][300] = 16'b1111111111101100;
    assign weights1[0][301] = 16'b0000000000000101;
    assign weights1[0][302] = 16'b0000000000011001;
    assign weights1[0][303] = 16'b0000000000011100;
    assign weights1[0][304] = 16'b0000000000011001;
    assign weights1[0][305] = 16'b0000000000011000;
    assign weights1[0][306] = 16'b0000000000011010;
    assign weights1[0][307] = 16'b0000000000011100;
    assign weights1[0][308] = 16'b0000000000001000;
    assign weights1[0][309] = 16'b0000000000010011;
    assign weights1[0][310] = 16'b0000000000100010;
    assign weights1[0][311] = 16'b0000000000101011;
    assign weights1[0][312] = 16'b0000000000110011;
    assign weights1[0][313] = 16'b0000000000111001;
    assign weights1[0][314] = 16'b0000000001000100;
    assign weights1[0][315] = 16'b0000000000101111;
    assign weights1[0][316] = 16'b0000000000011111;
    assign weights1[0][317] = 16'b0000000000010101;
    assign weights1[0][318] = 16'b0000000000001010;
    assign weights1[0][319] = 16'b1111111111111011;
    assign weights1[0][320] = 16'b1111111111101111;
    assign weights1[0][321] = 16'b1111111111111000;
    assign weights1[0][322] = 16'b1111111111100000;
    assign weights1[0][323] = 16'b1111111111100101;
    assign weights1[0][324] = 16'b1111111111111010;
    assign weights1[0][325] = 16'b1111111111110011;
    assign weights1[0][326] = 16'b1111111111100001;
    assign weights1[0][327] = 16'b1111111111110000;
    assign weights1[0][328] = 16'b1111111111101010;
    assign weights1[0][329] = 16'b0000000000000001;
    assign weights1[0][330] = 16'b0000000000010000;
    assign weights1[0][331] = 16'b0000000000001001;
    assign weights1[0][332] = 16'b0000000000001101;
    assign weights1[0][333] = 16'b0000000000011100;
    assign weights1[0][334] = 16'b0000000000011101;
    assign weights1[0][335] = 16'b0000000000001100;
    assign weights1[0][336] = 16'b0000000000011011;
    assign weights1[0][337] = 16'b0000000000101001;
    assign weights1[0][338] = 16'b0000000000110111;
    assign weights1[0][339] = 16'b0000000000111101;
    assign weights1[0][340] = 16'b0000000000111010;
    assign weights1[0][341] = 16'b0000000000100001;
    assign weights1[0][342] = 16'b0000000000010100;
    assign weights1[0][343] = 16'b1111111111101110;
    assign weights1[0][344] = 16'b0000000000001110;
    assign weights1[0][345] = 16'b0000000000000000;
    assign weights1[0][346] = 16'b1111111111110000;
    assign weights1[0][347] = 16'b0000000000000001;
    assign weights1[0][348] = 16'b1111111111110111;
    assign weights1[0][349] = 16'b1111111111110000;
    assign weights1[0][350] = 16'b1111111111101011;
    assign weights1[0][351] = 16'b1111111111110111;
    assign weights1[0][352] = 16'b1111111111101010;
    assign weights1[0][353] = 16'b1111111111110101;
    assign weights1[0][354] = 16'b1111111111101011;
    assign weights1[0][355] = 16'b1111111111101100;
    assign weights1[0][356] = 16'b1111111111111000;
    assign weights1[0][357] = 16'b1111111111110010;
    assign weights1[0][358] = 16'b0000000000000010;
    assign weights1[0][359] = 16'b0000000000001100;
    assign weights1[0][360] = 16'b0000000000010100;
    assign weights1[0][361] = 16'b0000000000000111;
    assign weights1[0][362] = 16'b0000000000010100;
    assign weights1[0][363] = 16'b0000000000010011;
    assign weights1[0][364] = 16'b0000000000101101;
    assign weights1[0][365] = 16'b0000000000101011;
    assign weights1[0][366] = 16'b0000000000110110;
    assign weights1[0][367] = 16'b0000000000111000;
    assign weights1[0][368] = 16'b0000000000101100;
    assign weights1[0][369] = 16'b0000000000001110;
    assign weights1[0][370] = 16'b0000000000000111;
    assign weights1[0][371] = 16'b0000000000000001;
    assign weights1[0][372] = 16'b0000000000001011;
    assign weights1[0][373] = 16'b1111111111110111;
    assign weights1[0][374] = 16'b0000000000011010;
    assign weights1[0][375] = 16'b1111111111111010;
    assign weights1[0][376] = 16'b1111111111110010;
    assign weights1[0][377] = 16'b1111111111101110;
    assign weights1[0][378] = 16'b1111111111011000;
    assign weights1[0][379] = 16'b1111111111110101;
    assign weights1[0][380] = 16'b1111111111101000;
    assign weights1[0][381] = 16'b1111111111110000;
    assign weights1[0][382] = 16'b1111111111100110;
    assign weights1[0][383] = 16'b1111111111111111;
    assign weights1[0][384] = 16'b1111111111110000;
    assign weights1[0][385] = 16'b1111111111101111;
    assign weights1[0][386] = 16'b0000000000001010;
    assign weights1[0][387] = 16'b1111111111110111;
    assign weights1[0][388] = 16'b1111111111111101;
    assign weights1[0][389] = 16'b0000000000001110;
    assign weights1[0][390] = 16'b0000000000000101;
    assign weights1[0][391] = 16'b0000000000010011;
    assign weights1[0][392] = 16'b0000000000110010;
    assign weights1[0][393] = 16'b0000000000010010;
    assign weights1[0][394] = 16'b0000000000011110;
    assign weights1[0][395] = 16'b0000000000010011;
    assign weights1[0][396] = 16'b0000000000001000;
    assign weights1[0][397] = 16'b0000000000010000;
    assign weights1[0][398] = 16'b0000000000000011;
    assign weights1[0][399] = 16'b0000000000010010;
    assign weights1[0][400] = 16'b1111111111111000;
    assign weights1[0][401] = 16'b0000000000000111;
    assign weights1[0][402] = 16'b0000000000000010;
    assign weights1[0][403] = 16'b0000000000001111;
    assign weights1[0][404] = 16'b0000000000000101;
    assign weights1[0][405] = 16'b1111111111111111;
    assign weights1[0][406] = 16'b0000000000000011;
    assign weights1[0][407] = 16'b1111111111100110;
    assign weights1[0][408] = 16'b1111111111111011;
    assign weights1[0][409] = 16'b1111111111111100;
    assign weights1[0][410] = 16'b1111111111100100;
    assign weights1[0][411] = 16'b1111111111111000;
    assign weights1[0][412] = 16'b1111111111101011;
    assign weights1[0][413] = 16'b1111111111110110;
    assign weights1[0][414] = 16'b0000000000000001;
    assign weights1[0][415] = 16'b0000000000010000;
    assign weights1[0][416] = 16'b1111111111111110;
    assign weights1[0][417] = 16'b1111111111101000;
    assign weights1[0][418] = 16'b1111111111111101;
    assign weights1[0][419] = 16'b0000000000011011;
    assign weights1[0][420] = 16'b0000000000010001;
    assign weights1[0][421] = 16'b0000000000010101;
    assign weights1[0][422] = 16'b1111111111111111;
    assign weights1[0][423] = 16'b0000000000010100;
    assign weights1[0][424] = 16'b1111111111110110;
    assign weights1[0][425] = 16'b0000000000000001;
    assign weights1[0][426] = 16'b0000000000001101;
    assign weights1[0][427] = 16'b1111111111110011;
    assign weights1[0][428] = 16'b0000000000010011;
    assign weights1[0][429] = 16'b1111111111111100;
    assign weights1[0][430] = 16'b0000000000001000;
    assign weights1[0][431] = 16'b0000000000000111;
    assign weights1[0][432] = 16'b0000000000000001;
    assign weights1[0][433] = 16'b0000000000000000;
    assign weights1[0][434] = 16'b1111111111110001;
    assign weights1[0][435] = 16'b1111111111101110;
    assign weights1[0][436] = 16'b1111111111111100;
    assign weights1[0][437] = 16'b1111111111101101;
    assign weights1[0][438] = 16'b1111111111101111;
    assign weights1[0][439] = 16'b1111111111110010;
    assign weights1[0][440] = 16'b1111111111111100;
    assign weights1[0][441] = 16'b0000000000001001;
    assign weights1[0][442] = 16'b1111111111111111;
    assign weights1[0][443] = 16'b1111111111111010;
    assign weights1[0][444] = 16'b0000000000001111;
    assign weights1[0][445] = 16'b0000000000001001;
    assign weights1[0][446] = 16'b0000000000000110;
    assign weights1[0][447] = 16'b0000000000100111;
    assign weights1[0][448] = 16'b0000000000010001;
    assign weights1[0][449] = 16'b0000000000001100;
    assign weights1[0][450] = 16'b1111111111110001;
    assign weights1[0][451] = 16'b0000000000000001;
    assign weights1[0][452] = 16'b1111111111111011;
    assign weights1[0][453] = 16'b0000000000010110;
    assign weights1[0][454] = 16'b1111111111111100;
    assign weights1[0][455] = 16'b0000000000010000;
    assign weights1[0][456] = 16'b0000000000000101;
    assign weights1[0][457] = 16'b0000000000001110;
    assign weights1[0][458] = 16'b0000000000000001;
    assign weights1[0][459] = 16'b0000000000001001;
    assign weights1[0][460] = 16'b0000000000000011;
    assign weights1[0][461] = 16'b0000000000000101;
    assign weights1[0][462] = 16'b1111111111111111;
    assign weights1[0][463] = 16'b0000000000001101;
    assign weights1[0][464] = 16'b1111111111100100;
    assign weights1[0][465] = 16'b0000000000000100;
    assign weights1[0][466] = 16'b1111111111101101;
    assign weights1[0][467] = 16'b1111111111101111;
    assign weights1[0][468] = 16'b1111111111110001;
    assign weights1[0][469] = 16'b1111111111110110;
    assign weights1[0][470] = 16'b1111111111111001;
    assign weights1[0][471] = 16'b1111111111110010;
    assign weights1[0][472] = 16'b1111111111101000;
    assign weights1[0][473] = 16'b0000000000000100;
    assign weights1[0][474] = 16'b0000000000000110;
    assign weights1[0][475] = 16'b0000000000100101;
    assign weights1[0][476] = 16'b0000000000000101;
    assign weights1[0][477] = 16'b0000000000010001;
    assign weights1[0][478] = 16'b0000000000001110;
    assign weights1[0][479] = 16'b1111111111110000;
    assign weights1[0][480] = 16'b0000000000001000;
    assign weights1[0][481] = 16'b0000000000000011;
    assign weights1[0][482] = 16'b0000000000010000;
    assign weights1[0][483] = 16'b0000000000001001;
    assign weights1[0][484] = 16'b0000000000011001;
    assign weights1[0][485] = 16'b0000000000000000;
    assign weights1[0][486] = 16'b0000000000000111;
    assign weights1[0][487] = 16'b0000000000001101;
    assign weights1[0][488] = 16'b1111111111110110;
    assign weights1[0][489] = 16'b0000000000000111;
    assign weights1[0][490] = 16'b1111111111111100;
    assign weights1[0][491] = 16'b1111111111110110;
    assign weights1[0][492] = 16'b1111111111111001;
    assign weights1[0][493] = 16'b1111111111101101;
    assign weights1[0][494] = 16'b1111111111111011;
    assign weights1[0][495] = 16'b1111111111111001;
    assign weights1[0][496] = 16'b1111111111101100;
    assign weights1[0][497] = 16'b1111111111110010;
    assign weights1[0][498] = 16'b1111111111101101;
    assign weights1[0][499] = 16'b1111111111110001;
    assign weights1[0][500] = 16'b1111111111111010;
    assign weights1[0][501] = 16'b0000000000001100;
    assign weights1[0][502] = 16'b0000000000010110;
    assign weights1[0][503] = 16'b0000000000011110;
    assign weights1[0][504] = 16'b0000000000001100;
    assign weights1[0][505] = 16'b0000000000010001;
    assign weights1[0][506] = 16'b0000000000000001;
    assign weights1[0][507] = 16'b1111111111111111;
    assign weights1[0][508] = 16'b1111111111111010;
    assign weights1[0][509] = 16'b0000000000010101;
    assign weights1[0][510] = 16'b0000000000000101;
    assign weights1[0][511] = 16'b1111111111101001;
    assign weights1[0][512] = 16'b0000000000011100;
    assign weights1[0][513] = 16'b0000000000000001;
    assign weights1[0][514] = 16'b1111111111111001;
    assign weights1[0][515] = 16'b0000000000001001;
    assign weights1[0][516] = 16'b0000000000001111;
    assign weights1[0][517] = 16'b1111111111110101;
    assign weights1[0][518] = 16'b1111111111110010;
    assign weights1[0][519] = 16'b1111111111100100;
    assign weights1[0][520] = 16'b1111111111110110;
    assign weights1[0][521] = 16'b1111111111110111;
    assign weights1[0][522] = 16'b1111111111110011;
    assign weights1[0][523] = 16'b1111111111111000;
    assign weights1[0][524] = 16'b1111111111100110;
    assign weights1[0][525] = 16'b0000000000000101;
    assign weights1[0][526] = 16'b1111111111111101;
    assign weights1[0][527] = 16'b0000000000011100;
    assign weights1[0][528] = 16'b0000000000010101;
    assign weights1[0][529] = 16'b1111111111111100;
    assign weights1[0][530] = 16'b0000000000000001;
    assign weights1[0][531] = 16'b0000000000010011;
    assign weights1[0][532] = 16'b0000000000010001;
    assign weights1[0][533] = 16'b0000000000010001;
    assign weights1[0][534] = 16'b0000000000001100;
    assign weights1[0][535] = 16'b1111111111110101;
    assign weights1[0][536] = 16'b0000000000000001;
    assign weights1[0][537] = 16'b0000000000010101;
    assign weights1[0][538] = 16'b0000000000001011;
    assign weights1[0][539] = 16'b0000000000000100;
    assign weights1[0][540] = 16'b0000000000001110;
    assign weights1[0][541] = 16'b0000000000000100;
    assign weights1[0][542] = 16'b0000000000000001;
    assign weights1[0][543] = 16'b0000000000000100;
    assign weights1[0][544] = 16'b0000000000001010;
    assign weights1[0][545] = 16'b0000000000001011;
    assign weights1[0][546] = 16'b1111111111101110;
    assign weights1[0][547] = 16'b0000000000000100;
    assign weights1[0][548] = 16'b1111111111110101;
    assign weights1[0][549] = 16'b1111111111110010;
    assign weights1[0][550] = 16'b1111111111111111;
    assign weights1[0][551] = 16'b0000000000000100;
    assign weights1[0][552] = 16'b1111111111111110;
    assign weights1[0][553] = 16'b1111111111101101;
    assign weights1[0][554] = 16'b0000000000000000;
    assign weights1[0][555] = 16'b1111111111100111;
    assign weights1[0][556] = 16'b0000000000000000;
    assign weights1[0][557] = 16'b1111111111110001;
    assign weights1[0][558] = 16'b0000000000001000;
    assign weights1[0][559] = 16'b0000000000001110;
    assign weights1[0][560] = 16'b0000000000000101;
    assign weights1[0][561] = 16'b0000000000001100;
    assign weights1[0][562] = 16'b0000000000001010;
    assign weights1[0][563] = 16'b0000000000001100;
    assign weights1[0][564] = 16'b0000000000000011;
    assign weights1[0][565] = 16'b0000000000001000;
    assign weights1[0][566] = 16'b0000000000001011;
    assign weights1[0][567] = 16'b0000000000001100;
    assign weights1[0][568] = 16'b1111111111111110;
    assign weights1[0][569] = 16'b0000000000001101;
    assign weights1[0][570] = 16'b1111111111111011;
    assign weights1[0][571] = 16'b0000000000000001;
    assign weights1[0][572] = 16'b1111111111111110;
    assign weights1[0][573] = 16'b0000000000000100;
    assign weights1[0][574] = 16'b1111111111110000;
    assign weights1[0][575] = 16'b0000000000000010;
    assign weights1[0][576] = 16'b1111111111111101;
    assign weights1[0][577] = 16'b1111111111101101;
    assign weights1[0][578] = 16'b1111111111111110;
    assign weights1[0][579] = 16'b1111111111111100;
    assign weights1[0][580] = 16'b1111111111101110;
    assign weights1[0][581] = 16'b0000000000001100;
    assign weights1[0][582] = 16'b1111111111100010;
    assign weights1[0][583] = 16'b1111111111101000;
    assign weights1[0][584] = 16'b1111111111110000;
    assign weights1[0][585] = 16'b1111111111101111;
    assign weights1[0][586] = 16'b1111111111111011;
    assign weights1[0][587] = 16'b0000000000000011;
    assign weights1[0][588] = 16'b0000000000000010;
    assign weights1[0][589] = 16'b0000000000001010;
    assign weights1[0][590] = 16'b0000000000000100;
    assign weights1[0][591] = 16'b0000000000001011;
    assign weights1[0][592] = 16'b1111111111111010;
    assign weights1[0][593] = 16'b1111111111111000;
    assign weights1[0][594] = 16'b0000000000000010;
    assign weights1[0][595] = 16'b1111111111110100;
    assign weights1[0][596] = 16'b1111111111111110;
    assign weights1[0][597] = 16'b0000000000001001;
    assign weights1[0][598] = 16'b0000000000000011;
    assign weights1[0][599] = 16'b1111111111101110;
    assign weights1[0][600] = 16'b1111111111110011;
    assign weights1[0][601] = 16'b1111111111111100;
    assign weights1[0][602] = 16'b0000000000000011;
    assign weights1[0][603] = 16'b1111111111110101;
    assign weights1[0][604] = 16'b1111111111111111;
    assign weights1[0][605] = 16'b1111111111111001;
    assign weights1[0][606] = 16'b1111111111110111;
    assign weights1[0][607] = 16'b0000000000000100;
    assign weights1[0][608] = 16'b1111111111111110;
    assign weights1[0][609] = 16'b0000000000010001;
    assign weights1[0][610] = 16'b1111111111111110;
    assign weights1[0][611] = 16'b1111111111111100;
    assign weights1[0][612] = 16'b1111111111110011;
    assign weights1[0][613] = 16'b1111111111110011;
    assign weights1[0][614] = 16'b1111111111111000;
    assign weights1[0][615] = 16'b0000000000000001;
    assign weights1[0][616] = 16'b1111111111111110;
    assign weights1[0][617] = 16'b0000000000000100;
    assign weights1[0][618] = 16'b0000000000000101;
    assign weights1[0][619] = 16'b0000000000000111;
    assign weights1[0][620] = 16'b0000000000001000;
    assign weights1[0][621] = 16'b1111111111111100;
    assign weights1[0][622] = 16'b0000000000000101;
    assign weights1[0][623] = 16'b0000000000100001;
    assign weights1[0][624] = 16'b1111111111110001;
    assign weights1[0][625] = 16'b0000000000000011;
    assign weights1[0][626] = 16'b1111111111110001;
    assign weights1[0][627] = 16'b1111111111111101;
    assign weights1[0][628] = 16'b1111111111111100;
    assign weights1[0][629] = 16'b1111111111101111;
    assign weights1[0][630] = 16'b0000000000000010;
    assign weights1[0][631] = 16'b1111111111100010;
    assign weights1[0][632] = 16'b0000000000000110;
    assign weights1[0][633] = 16'b0000000000001011;
    assign weights1[0][634] = 16'b0000000000001000;
    assign weights1[0][635] = 16'b1111111111111011;
    assign weights1[0][636] = 16'b1111111111111110;
    assign weights1[0][637] = 16'b0000000000001000;
    assign weights1[0][638] = 16'b0000000000000000;
    assign weights1[0][639] = 16'b0000000000000000;
    assign weights1[0][640] = 16'b1111111111110100;
    assign weights1[0][641] = 16'b1111111111111100;
    assign weights1[0][642] = 16'b1111111111111100;
    assign weights1[0][643] = 16'b1111111111110110;
    assign weights1[0][644] = 16'b0000000000000010;
    assign weights1[0][645] = 16'b0000000000000001;
    assign weights1[0][646] = 16'b1111111111111101;
    assign weights1[0][647] = 16'b1111111111110110;
    assign weights1[0][648] = 16'b1111111111111001;
    assign weights1[0][649] = 16'b0000000000000001;
    assign weights1[0][650] = 16'b1111111111111010;
    assign weights1[0][651] = 16'b1111111111110101;
    assign weights1[0][652] = 16'b1111111111111100;
    assign weights1[0][653] = 16'b1111111111110001;
    assign weights1[0][654] = 16'b0000000000000101;
    assign weights1[0][655] = 16'b1111111111111000;
    assign weights1[0][656] = 16'b0000000000000101;
    assign weights1[0][657] = 16'b1111111111100010;
    assign weights1[0][658] = 16'b1111111111011100;
    assign weights1[0][659] = 16'b0000000000000101;
    assign weights1[0][660] = 16'b1111111111111011;
    assign weights1[0][661] = 16'b1111111111110110;
    assign weights1[0][662] = 16'b1111111111111111;
    assign weights1[0][663] = 16'b0000000000010101;
    assign weights1[0][664] = 16'b1111111111110001;
    assign weights1[0][665] = 16'b0000000000000010;
    assign weights1[0][666] = 16'b0000000000000101;
    assign weights1[0][667] = 16'b1111111111111101;
    assign weights1[0][668] = 16'b1111111111110010;
    assign weights1[0][669] = 16'b1111111111110101;
    assign weights1[0][670] = 16'b1111111111110100;
    assign weights1[0][671] = 16'b1111111111111001;
    assign weights1[0][672] = 16'b1111111111111011;
    assign weights1[0][673] = 16'b1111111111111101;
    assign weights1[0][674] = 16'b1111111111111011;
    assign weights1[0][675] = 16'b1111111111111010;
    assign weights1[0][676] = 16'b1111111111110001;
    assign weights1[0][677] = 16'b1111111111110110;
    assign weights1[0][678] = 16'b1111111111101000;
    assign weights1[0][679] = 16'b1111111111011100;
    assign weights1[0][680] = 16'b0000000000001110;
    assign weights1[0][681] = 16'b1111111111011001;
    assign weights1[0][682] = 16'b1111111111111101;
    assign weights1[0][683] = 16'b1111111111111010;
    assign weights1[0][684] = 16'b0000000000000011;
    assign weights1[0][685] = 16'b0000000000010000;
    assign weights1[0][686] = 16'b1111111111111101;
    assign weights1[0][687] = 16'b1111111111111111;
    assign weights1[0][688] = 16'b1111111111111111;
    assign weights1[0][689] = 16'b1111111111110011;
    assign weights1[0][690] = 16'b0000000000000111;
    assign weights1[0][691] = 16'b0000000000000100;
    assign weights1[0][692] = 16'b1111111111111010;
    assign weights1[0][693] = 16'b0000000000000011;
    assign weights1[0][694] = 16'b0000000000000110;
    assign weights1[0][695] = 16'b0000000000000011;
    assign weights1[0][696] = 16'b1111111111110110;
    assign weights1[0][697] = 16'b1111111111111001;
    assign weights1[0][698] = 16'b1111111111111101;
    assign weights1[0][699] = 16'b0000000000000000;
    assign weights1[0][700] = 16'b1111111111111110;
    assign weights1[0][701] = 16'b0000000000000000;
    assign weights1[0][702] = 16'b0000000000000100;
    assign weights1[0][703] = 16'b1111111111111101;
    assign weights1[0][704] = 16'b1111111111111010;
    assign weights1[0][705] = 16'b1111111111101101;
    assign weights1[0][706] = 16'b1111111111101111;
    assign weights1[0][707] = 16'b1111111111110101;
    assign weights1[0][708] = 16'b1111111111110111;
    assign weights1[0][709] = 16'b0000000000000000;
    assign weights1[0][710] = 16'b0000000000000001;
    assign weights1[0][711] = 16'b0000000000010000;
    assign weights1[0][712] = 16'b0000000000000101;
    assign weights1[0][713] = 16'b1111111111111001;
    assign weights1[0][714] = 16'b0000000000001010;
    assign weights1[0][715] = 16'b1111111111111001;
    assign weights1[0][716] = 16'b1111111111110100;
    assign weights1[0][717] = 16'b1111111111011010;
    assign weights1[0][718] = 16'b1111111111110011;
    assign weights1[0][719] = 16'b0000000000000001;
    assign weights1[0][720] = 16'b1111111111111111;
    assign weights1[0][721] = 16'b1111111111110111;
    assign weights1[0][722] = 16'b1111111111111110;
    assign weights1[0][723] = 16'b0000000000000000;
    assign weights1[0][724] = 16'b0000000000000100;
    assign weights1[0][725] = 16'b1111111111111111;
    assign weights1[0][726] = 16'b1111111111111111;
    assign weights1[0][727] = 16'b0000000000000100;
    assign weights1[0][728] = 16'b0000000000000000;
    assign weights1[0][729] = 16'b0000000000000010;
    assign weights1[0][730] = 16'b0000000000000001;
    assign weights1[0][731] = 16'b1111111111111100;
    assign weights1[0][732] = 16'b1111111111111010;
    assign weights1[0][733] = 16'b1111111111110110;
    assign weights1[0][734] = 16'b0000000000000110;
    assign weights1[0][735] = 16'b1111111111111001;
    assign weights1[0][736] = 16'b0000000000000011;
    assign weights1[0][737] = 16'b0000000000000001;
    assign weights1[0][738] = 16'b0000000000000110;
    assign weights1[0][739] = 16'b1111111111110100;
    assign weights1[0][740] = 16'b0000000000000011;
    assign weights1[0][741] = 16'b0000000000000001;
    assign weights1[0][742] = 16'b0000000000000100;
    assign weights1[0][743] = 16'b1111111111111010;
    assign weights1[0][744] = 16'b1111111111110111;
    assign weights1[0][745] = 16'b1111111111110000;
    assign weights1[0][746] = 16'b1111111111101011;
    assign weights1[0][747] = 16'b1111111111110010;
    assign weights1[0][748] = 16'b1111111111111110;
    assign weights1[0][749] = 16'b1111111111111001;
    assign weights1[0][750] = 16'b1111111111110001;
    assign weights1[0][751] = 16'b1111111111110111;
    assign weights1[0][752] = 16'b1111111111111011;
    assign weights1[0][753] = 16'b1111111111111010;
    assign weights1[0][754] = 16'b1111111111111100;
    assign weights1[0][755] = 16'b0000000000000001;
    assign weights1[0][756] = 16'b0000000000000000;
    assign weights1[0][757] = 16'b0000000000000000;
    assign weights1[0][758] = 16'b1111111111111101;
    assign weights1[0][759] = 16'b1111111111111111;
    assign weights1[0][760] = 16'b1111111111111010;
    assign weights1[0][761] = 16'b1111111111111000;
    assign weights1[0][762] = 16'b1111111111111111;
    assign weights1[0][763] = 16'b1111111111111110;
    assign weights1[0][764] = 16'b0000000000001001;
    assign weights1[0][765] = 16'b1111111111110111;
    assign weights1[0][766] = 16'b1111111111111110;
    assign weights1[0][767] = 16'b0000000000000111;
    assign weights1[0][768] = 16'b0000000000000100;
    assign weights1[0][769] = 16'b1111111111110100;
    assign weights1[0][770] = 16'b0000000000000011;
    assign weights1[0][771] = 16'b1111111111111101;
    assign weights1[0][772] = 16'b1111111111111001;
    assign weights1[0][773] = 16'b1111111111111000;
    assign weights1[0][774] = 16'b1111111111101001;
    assign weights1[0][775] = 16'b1111111111110101;
    assign weights1[0][776] = 16'b1111111111101110;
    assign weights1[0][777] = 16'b1111111111111001;
    assign weights1[0][778] = 16'b1111111111111011;
    assign weights1[0][779] = 16'b1111111111111100;
    assign weights1[0][780] = 16'b1111111111111011;
    assign weights1[0][781] = 16'b1111111111111110;
    assign weights1[0][782] = 16'b1111111111111111;
    assign weights1[0][783] = 16'b0000000000000000;
    assign weights1[1][0] = 16'b0000000000000000;
    assign weights1[1][1] = 16'b0000000000000000;
    assign weights1[1][2] = 16'b1111111111111110;
    assign weights1[1][3] = 16'b1111111111111111;
    assign weights1[1][4] = 16'b0000000000000000;
    assign weights1[1][5] = 16'b1111111111111110;
    assign weights1[1][6] = 16'b0000000000000001;
    assign weights1[1][7] = 16'b1111111111111000;
    assign weights1[1][8] = 16'b0000000000000000;
    assign weights1[1][9] = 16'b1111111111110110;
    assign weights1[1][10] = 16'b1111111111110001;
    assign weights1[1][11] = 16'b1111111111101100;
    assign weights1[1][12] = 16'b1111111111101010;
    assign weights1[1][13] = 16'b1111111111101101;
    assign weights1[1][14] = 16'b1111111111111010;
    assign weights1[1][15] = 16'b1111111111110101;
    assign weights1[1][16] = 16'b1111111111110000;
    assign weights1[1][17] = 16'b1111111111101100;
    assign weights1[1][18] = 16'b1111111111110101;
    assign weights1[1][19] = 16'b1111111111111001;
    assign weights1[1][20] = 16'b0000000000000011;
    assign weights1[1][21] = 16'b0000000000000010;
    assign weights1[1][22] = 16'b0000000000000011;
    assign weights1[1][23] = 16'b0000000000000011;
    assign weights1[1][24] = 16'b1111111111111111;
    assign weights1[1][25] = 16'b0000000000000000;
    assign weights1[1][26] = 16'b1111111111111110;
    assign weights1[1][27] = 16'b0000000000000000;
    assign weights1[1][28] = 16'b0000000000000000;
    assign weights1[1][29] = 16'b0000000000000000;
    assign weights1[1][30] = 16'b0000000000000010;
    assign weights1[1][31] = 16'b0000000000000001;
    assign weights1[1][32] = 16'b0000000000000100;
    assign weights1[1][33] = 16'b0000000000000110;
    assign weights1[1][34] = 16'b0000000000000110;
    assign weights1[1][35] = 16'b1111111111111110;
    assign weights1[1][36] = 16'b0000000000001011;
    assign weights1[1][37] = 16'b1111111111111011;
    assign weights1[1][38] = 16'b1111111111111000;
    assign weights1[1][39] = 16'b0000000000000001;
    assign weights1[1][40] = 16'b1111111111111000;
    assign weights1[1][41] = 16'b1111111111111011;
    assign weights1[1][42] = 16'b1111111111111100;
    assign weights1[1][43] = 16'b0000000000000100;
    assign weights1[1][44] = 16'b1111111111101100;
    assign weights1[1][45] = 16'b1111111111111000;
    assign weights1[1][46] = 16'b1111111111101111;
    assign weights1[1][47] = 16'b0000000000000011;
    assign weights1[1][48] = 16'b1111111111111101;
    assign weights1[1][49] = 16'b1111111111111110;
    assign weights1[1][50] = 16'b0000000000001101;
    assign weights1[1][51] = 16'b0000000000001001;
    assign weights1[1][52] = 16'b1111111111111111;
    assign weights1[1][53] = 16'b1111111111110011;
    assign weights1[1][54] = 16'b1111111111111100;
    assign weights1[1][55] = 16'b0000000000000000;
    assign weights1[1][56] = 16'b0000000000000000;
    assign weights1[1][57] = 16'b1111111111111111;
    assign weights1[1][58] = 16'b0000000000000011;
    assign weights1[1][59] = 16'b1111111111111011;
    assign weights1[1][60] = 16'b0000000000000111;
    assign weights1[1][61] = 16'b0000000000000011;
    assign weights1[1][62] = 16'b1111111111111011;
    assign weights1[1][63] = 16'b0000000000001000;
    assign weights1[1][64] = 16'b1111111111110110;
    assign weights1[1][65] = 16'b1111111111111100;
    assign weights1[1][66] = 16'b1111111111111111;
    assign weights1[1][67] = 16'b1111111111111111;
    assign weights1[1][68] = 16'b0000000000010111;
    assign weights1[1][69] = 16'b0000000000001011;
    assign weights1[1][70] = 16'b0000000000000010;
    assign weights1[1][71] = 16'b0000000000000001;
    assign weights1[1][72] = 16'b0000000000001000;
    assign weights1[1][73] = 16'b1111111111101010;
    assign weights1[1][74] = 16'b0000000000001010;
    assign weights1[1][75] = 16'b1111111111111101;
    assign weights1[1][76] = 16'b0000000000001010;
    assign weights1[1][77] = 16'b0000000000000000;
    assign weights1[1][78] = 16'b0000000000000000;
    assign weights1[1][79] = 16'b0000000000000010;
    assign weights1[1][80] = 16'b0000000000000011;
    assign weights1[1][81] = 16'b1111111111111010;
    assign weights1[1][82] = 16'b1111111111111001;
    assign weights1[1][83] = 16'b0000000000000000;
    assign weights1[1][84] = 16'b0000000000000000;
    assign weights1[1][85] = 16'b0000000000000001;
    assign weights1[1][86] = 16'b1111111111111010;
    assign weights1[1][87] = 16'b1111111111111011;
    assign weights1[1][88] = 16'b1111111111111110;
    assign weights1[1][89] = 16'b0000000000000100;
    assign weights1[1][90] = 16'b0000000000000000;
    assign weights1[1][91] = 16'b0000000000000111;
    assign weights1[1][92] = 16'b1111111111111001;
    assign weights1[1][93] = 16'b0000000000000011;
    assign weights1[1][94] = 16'b1111111111111011;
    assign weights1[1][95] = 16'b1111111111111110;
    assign weights1[1][96] = 16'b1111111111110111;
    assign weights1[1][97] = 16'b0000000000001011;
    assign weights1[1][98] = 16'b0000000000000110;
    assign weights1[1][99] = 16'b1111111111111001;
    assign weights1[1][100] = 16'b0000000000000010;
    assign weights1[1][101] = 16'b0000000000010010;
    assign weights1[1][102] = 16'b1111111111111111;
    assign weights1[1][103] = 16'b1111111111111011;
    assign weights1[1][104] = 16'b1111111111111011;
    assign weights1[1][105] = 16'b1111111111110111;
    assign weights1[1][106] = 16'b0000000000000110;
    assign weights1[1][107] = 16'b1111111111110111;
    assign weights1[1][108] = 16'b1111111111110101;
    assign weights1[1][109] = 16'b0000000000000001;
    assign weights1[1][110] = 16'b0000000000001011;
    assign weights1[1][111] = 16'b0000000000000111;
    assign weights1[1][112] = 16'b1111111111111110;
    assign weights1[1][113] = 16'b1111111111110111;
    assign weights1[1][114] = 16'b1111111111111001;
    assign weights1[1][115] = 16'b1111111111110101;
    assign weights1[1][116] = 16'b1111111111111101;
    assign weights1[1][117] = 16'b1111111111111000;
    assign weights1[1][118] = 16'b0000000000000100;
    assign weights1[1][119] = 16'b0000000000010101;
    assign weights1[1][120] = 16'b0000000000000101;
    assign weights1[1][121] = 16'b0000000000010000;
    assign weights1[1][122] = 16'b0000000000001100;
    assign weights1[1][123] = 16'b0000000000000011;
    assign weights1[1][124] = 16'b0000000000010110;
    assign weights1[1][125] = 16'b1111111111110011;
    assign weights1[1][126] = 16'b1111111111111100;
    assign weights1[1][127] = 16'b0000000000001100;
    assign weights1[1][128] = 16'b1111111111110101;
    assign weights1[1][129] = 16'b0000000000001010;
    assign weights1[1][130] = 16'b1111111111101100;
    assign weights1[1][131] = 16'b1111111111111110;
    assign weights1[1][132] = 16'b0000000000010000;
    assign weights1[1][133] = 16'b1111111111110000;
    assign weights1[1][134] = 16'b1111111111110010;
    assign weights1[1][135] = 16'b1111111111110101;
    assign weights1[1][136] = 16'b1111111111111010;
    assign weights1[1][137] = 16'b0000000000000101;
    assign weights1[1][138] = 16'b0000000000001000;
    assign weights1[1][139] = 16'b0000000000000100;
    assign weights1[1][140] = 16'b1111111111111100;
    assign weights1[1][141] = 16'b1111111111111101;
    assign weights1[1][142] = 16'b1111111111111010;
    assign weights1[1][143] = 16'b1111111111111010;
    assign weights1[1][144] = 16'b1111111111111010;
    assign weights1[1][145] = 16'b1111111111111100;
    assign weights1[1][146] = 16'b0000000000011010;
    assign weights1[1][147] = 16'b0000000000010000;
    assign weights1[1][148] = 16'b0000000000000101;
    assign weights1[1][149] = 16'b0000000000001011;
    assign weights1[1][150] = 16'b1111111111111000;
    assign weights1[1][151] = 16'b0000000000001001;
    assign weights1[1][152] = 16'b1111111111111111;
    assign weights1[1][153] = 16'b0000000000000111;
    assign weights1[1][154] = 16'b0000000000001101;
    assign weights1[1][155] = 16'b1111111111110101;
    assign weights1[1][156] = 16'b1111111111111111;
    assign weights1[1][157] = 16'b0000000000000110;
    assign weights1[1][158] = 16'b0000000000001000;
    assign weights1[1][159] = 16'b0000000000001000;
    assign weights1[1][160] = 16'b0000000000001011;
    assign weights1[1][161] = 16'b0000000000000110;
    assign weights1[1][162] = 16'b1111111111111111;
    assign weights1[1][163] = 16'b0000000000000000;
    assign weights1[1][164] = 16'b0000000000001111;
    assign weights1[1][165] = 16'b1111111111111101;
    assign weights1[1][166] = 16'b0000000000010111;
    assign weights1[1][167] = 16'b0000000000001001;
    assign weights1[1][168] = 16'b0000000000000001;
    assign weights1[1][169] = 16'b0000000000001101;
    assign weights1[1][170] = 16'b0000000000010111;
    assign weights1[1][171] = 16'b0000000000001001;
    assign weights1[1][172] = 16'b0000000000000011;
    assign weights1[1][173] = 16'b1111111111111001;
    assign weights1[1][174] = 16'b1111111111110101;
    assign weights1[1][175] = 16'b0000000000000001;
    assign weights1[1][176] = 16'b0000000000001101;
    assign weights1[1][177] = 16'b0000000000000010;
    assign weights1[1][178] = 16'b0000000000001001;
    assign weights1[1][179] = 16'b0000000000001000;
    assign weights1[1][180] = 16'b0000000000000100;
    assign weights1[1][181] = 16'b1111111111111010;
    assign weights1[1][182] = 16'b0000000000000111;
    assign weights1[1][183] = 16'b0000000000000101;
    assign weights1[1][184] = 16'b0000000000010000;
    assign weights1[1][185] = 16'b1111111111111000;
    assign weights1[1][186] = 16'b0000000000001011;
    assign weights1[1][187] = 16'b1111111111100101;
    assign weights1[1][188] = 16'b0000000000010000;
    assign weights1[1][189] = 16'b1111111111101101;
    assign weights1[1][190] = 16'b0000000000011010;
    assign weights1[1][191] = 16'b0000000000001110;
    assign weights1[1][192] = 16'b0000000000001100;
    assign weights1[1][193] = 16'b0000000000000001;
    assign weights1[1][194] = 16'b1111111111111001;
    assign weights1[1][195] = 16'b0000000000001001;
    assign weights1[1][196] = 16'b0000000000001000;
    assign weights1[1][197] = 16'b1111111111111101;
    assign weights1[1][198] = 16'b1111111111111001;
    assign weights1[1][199] = 16'b1111111111111011;
    assign weights1[1][200] = 16'b0000000000000011;
    assign weights1[1][201] = 16'b1111111111111111;
    assign weights1[1][202] = 16'b0000000000010100;
    assign weights1[1][203] = 16'b0000000000000101;
    assign weights1[1][204] = 16'b0000000000010001;
    assign weights1[1][205] = 16'b1111111111111101;
    assign weights1[1][206] = 16'b0000000000000000;
    assign weights1[1][207] = 16'b1111111111111111;
    assign weights1[1][208] = 16'b0000000000000100;
    assign weights1[1][209] = 16'b0000000000010101;
    assign weights1[1][210] = 16'b0000000000001110;
    assign weights1[1][211] = 16'b1111111111111011;
    assign weights1[1][212] = 16'b0000000000000101;
    assign weights1[1][213] = 16'b1111111111111110;
    assign weights1[1][214] = 16'b1111111111111110;
    assign weights1[1][215] = 16'b0000000000000011;
    assign weights1[1][216] = 16'b0000000000001011;
    assign weights1[1][217] = 16'b0000000000001110;
    assign weights1[1][218] = 16'b0000000000000110;
    assign weights1[1][219] = 16'b1111111111111011;
    assign weights1[1][220] = 16'b1111111111110100;
    assign weights1[1][221] = 16'b0000000000000000;
    assign weights1[1][222] = 16'b0000000000000011;
    assign weights1[1][223] = 16'b0000000000000011;
    assign weights1[1][224] = 16'b0000000000000100;
    assign weights1[1][225] = 16'b0000000000000110;
    assign weights1[1][226] = 16'b1111111111111101;
    assign weights1[1][227] = 16'b0000000000000000;
    assign weights1[1][228] = 16'b1111111111111110;
    assign weights1[1][229] = 16'b0000000000001000;
    assign weights1[1][230] = 16'b1111111111110100;
    assign weights1[1][231] = 16'b0000000000000000;
    assign weights1[1][232] = 16'b0000000000000100;
    assign weights1[1][233] = 16'b0000000000001000;
    assign weights1[1][234] = 16'b1111111111111101;
    assign weights1[1][235] = 16'b0000000000001111;
    assign weights1[1][236] = 16'b1111111111111100;
    assign weights1[1][237] = 16'b0000000000000011;
    assign weights1[1][238] = 16'b0000000000000001;
    assign weights1[1][239] = 16'b1111111111111011;
    assign weights1[1][240] = 16'b0000000000001101;
    assign weights1[1][241] = 16'b0000000000010000;
    assign weights1[1][242] = 16'b0000000000010111;
    assign weights1[1][243] = 16'b0000000000000110;
    assign weights1[1][244] = 16'b1111111111100110;
    assign weights1[1][245] = 16'b0000000000000100;
    assign weights1[1][246] = 16'b1111111111111001;
    assign weights1[1][247] = 16'b1111111111110011;
    assign weights1[1][248] = 16'b0000000000000100;
    assign weights1[1][249] = 16'b0000000000000011;
    assign weights1[1][250] = 16'b1111111111110110;
    assign weights1[1][251] = 16'b0000000000001110;
    assign weights1[1][252] = 16'b0000000000000001;
    assign weights1[1][253] = 16'b1111111111111111;
    assign weights1[1][254] = 16'b1111111111111010;
    assign weights1[1][255] = 16'b0000000000001100;
    assign weights1[1][256] = 16'b0000000000010110;
    assign weights1[1][257] = 16'b0000000000000010;
    assign weights1[1][258] = 16'b0000000000000100;
    assign weights1[1][259] = 16'b0000000000010001;
    assign weights1[1][260] = 16'b1111111111101001;
    assign weights1[1][261] = 16'b1111111111111000;
    assign weights1[1][262] = 16'b0000000000000111;
    assign weights1[1][263] = 16'b0000000000001111;
    assign weights1[1][264] = 16'b0000000000010000;
    assign weights1[1][265] = 16'b0000000000010011;
    assign weights1[1][266] = 16'b0000000000000110;
    assign weights1[1][267] = 16'b0000000000001101;
    assign weights1[1][268] = 16'b1111111111110101;
    assign weights1[1][269] = 16'b1111111111111110;
    assign weights1[1][270] = 16'b0000000000000111;
    assign weights1[1][271] = 16'b0000000000001011;
    assign weights1[1][272] = 16'b0000000000000000;
    assign weights1[1][273] = 16'b1111111111110100;
    assign weights1[1][274] = 16'b1111111111111110;
    assign weights1[1][275] = 16'b1111111111111101;
    assign weights1[1][276] = 16'b1111111111101011;
    assign weights1[1][277] = 16'b1111111111111101;
    assign weights1[1][278] = 16'b0000000000000100;
    assign weights1[1][279] = 16'b1111111111110111;
    assign weights1[1][280] = 16'b0000000000001000;
    assign weights1[1][281] = 16'b0000000000011101;
    assign weights1[1][282] = 16'b0000000000001001;
    assign weights1[1][283] = 16'b0000000000011000;
    assign weights1[1][284] = 16'b1111111111111100;
    assign weights1[1][285] = 16'b1111111111111111;
    assign weights1[1][286] = 16'b0000000000000001;
    assign weights1[1][287] = 16'b0000000000000100;
    assign weights1[1][288] = 16'b0000000000001010;
    assign weights1[1][289] = 16'b1111111111110111;
    assign weights1[1][290] = 16'b1111111111111111;
    assign weights1[1][291] = 16'b0000000000000001;
    assign weights1[1][292] = 16'b0000000000001110;
    assign weights1[1][293] = 16'b1111111111110000;
    assign weights1[1][294] = 16'b0000000000000000;
    assign weights1[1][295] = 16'b0000000000000000;
    assign weights1[1][296] = 16'b1111111111111001;
    assign weights1[1][297] = 16'b1111111111111011;
    assign weights1[1][298] = 16'b1111111111111100;
    assign weights1[1][299] = 16'b1111111111110011;
    assign weights1[1][300] = 16'b0000000000010010;
    assign weights1[1][301] = 16'b1111111111111111;
    assign weights1[1][302] = 16'b1111111111110100;
    assign weights1[1][303] = 16'b1111111111111101;
    assign weights1[1][304] = 16'b0000000000000001;
    assign weights1[1][305] = 16'b0000000000000100;
    assign weights1[1][306] = 16'b0000000000000010;
    assign weights1[1][307] = 16'b0000000000001010;
    assign weights1[1][308] = 16'b1111111111111011;
    assign weights1[1][309] = 16'b0000000000001000;
    assign weights1[1][310] = 16'b1111111111110111;
    assign weights1[1][311] = 16'b1111111111111111;
    assign weights1[1][312] = 16'b0000000000010010;
    assign weights1[1][313] = 16'b1111111111111010;
    assign weights1[1][314] = 16'b1111111111111001;
    assign weights1[1][315] = 16'b1111111111111001;
    assign weights1[1][316] = 16'b1111111111111000;
    assign weights1[1][317] = 16'b0000000000000001;
    assign weights1[1][318] = 16'b0000000000010001;
    assign weights1[1][319] = 16'b1111111111101100;
    assign weights1[1][320] = 16'b1111111111111110;
    assign weights1[1][321] = 16'b0000000000000011;
    assign weights1[1][322] = 16'b1111111111110111;
    assign weights1[1][323] = 16'b1111111111111010;
    assign weights1[1][324] = 16'b1111111111110100;
    assign weights1[1][325] = 16'b1111111111111000;
    assign weights1[1][326] = 16'b0000000000001001;
    assign weights1[1][327] = 16'b0000000000000111;
    assign weights1[1][328] = 16'b1111111111111000;
    assign weights1[1][329] = 16'b1111111111111100;
    assign weights1[1][330] = 16'b0000000000010011;
    assign weights1[1][331] = 16'b1111111111111011;
    assign weights1[1][332] = 16'b1111111111110000;
    assign weights1[1][333] = 16'b1111111111111100;
    assign weights1[1][334] = 16'b0000000000000001;
    assign weights1[1][335] = 16'b0000000000000110;
    assign weights1[1][336] = 16'b1111111111110000;
    assign weights1[1][337] = 16'b1111111111111010;
    assign weights1[1][338] = 16'b1111111111111101;
    assign weights1[1][339] = 16'b0000000000000000;
    assign weights1[1][340] = 16'b0000000000000100;
    assign weights1[1][341] = 16'b1111111111111011;
    assign weights1[1][342] = 16'b1111111111111110;
    assign weights1[1][343] = 16'b1111111111101111;
    assign weights1[1][344] = 16'b1111111111110001;
    assign weights1[1][345] = 16'b1111111111111000;
    assign weights1[1][346] = 16'b1111111111101110;
    assign weights1[1][347] = 16'b1111111111111101;
    assign weights1[1][348] = 16'b1111111111110110;
    assign weights1[1][349] = 16'b0000000000000011;
    assign weights1[1][350] = 16'b1111111111111110;
    assign weights1[1][351] = 16'b1111111111111110;
    assign weights1[1][352] = 16'b1111111111111100;
    assign weights1[1][353] = 16'b0000000000000000;
    assign weights1[1][354] = 16'b1111111111110100;
    assign weights1[1][355] = 16'b1111111111100101;
    assign weights1[1][356] = 16'b1111111111111001;
    assign weights1[1][357] = 16'b1111111111111101;
    assign weights1[1][358] = 16'b0000000000000010;
    assign weights1[1][359] = 16'b1111111111111110;
    assign weights1[1][360] = 16'b0000000000000010;
    assign weights1[1][361] = 16'b1111111111110000;
    assign weights1[1][362] = 16'b1111111111111100;
    assign weights1[1][363] = 16'b1111111111111011;
    assign weights1[1][364] = 16'b1111111111100100;
    assign weights1[1][365] = 16'b1111111111100110;
    assign weights1[1][366] = 16'b1111111111101110;
    assign weights1[1][367] = 16'b1111111111111111;
    assign weights1[1][368] = 16'b0000000000001011;
    assign weights1[1][369] = 16'b0000000000001110;
    assign weights1[1][370] = 16'b1111111111111101;
    assign weights1[1][371] = 16'b1111111111110001;
    assign weights1[1][372] = 16'b1111111111110110;
    assign weights1[1][373] = 16'b0000000000010110;
    assign weights1[1][374] = 16'b1111111111110001;
    assign weights1[1][375] = 16'b0000000000001010;
    assign weights1[1][376] = 16'b0000000000011110;
    assign weights1[1][377] = 16'b0000000000011000;
    assign weights1[1][378] = 16'b0000000000010110;
    assign weights1[1][379] = 16'b0000000000001100;
    assign weights1[1][380] = 16'b0000000000001001;
    assign weights1[1][381] = 16'b0000000000001001;
    assign weights1[1][382] = 16'b1111111111111101;
    assign weights1[1][383] = 16'b1111111111111101;
    assign weights1[1][384] = 16'b1111111111111001;
    assign weights1[1][385] = 16'b1111111111100010;
    assign weights1[1][386] = 16'b1111111111111100;
    assign weights1[1][387] = 16'b1111111111110011;
    assign weights1[1][388] = 16'b0000000000000111;
    assign weights1[1][389] = 16'b0000000000000111;
    assign weights1[1][390] = 16'b1111111111110110;
    assign weights1[1][391] = 16'b1111111111111010;
    assign weights1[1][392] = 16'b1111111111011001;
    assign weights1[1][393] = 16'b1111111110111111;
    assign weights1[1][394] = 16'b1111111111010001;
    assign weights1[1][395] = 16'b1111111111100000;
    assign weights1[1][396] = 16'b0000000000000111;
    assign weights1[1][397] = 16'b0000000000010001;
    assign weights1[1][398] = 16'b0000000000011101;
    assign weights1[1][399] = 16'b0000000000010110;
    assign weights1[1][400] = 16'b0000000000100010;
    assign weights1[1][401] = 16'b0000000000010000;
    assign weights1[1][402] = 16'b0000000000000000;
    assign weights1[1][403] = 16'b0000000000001011;
    assign weights1[1][404] = 16'b0000000000011001;
    assign weights1[1][405] = 16'b0000000000010101;
    assign weights1[1][406] = 16'b0000000000001011;
    assign weights1[1][407] = 16'b0000000000010010;
    assign weights1[1][408] = 16'b0000000000000001;
    assign weights1[1][409] = 16'b1111111111101001;
    assign weights1[1][410] = 16'b0000000000000101;
    assign weights1[1][411] = 16'b0000000000000010;
    assign weights1[1][412] = 16'b1111111111111101;
    assign weights1[1][413] = 16'b0000000000001011;
    assign weights1[1][414] = 16'b1111111111100111;
    assign weights1[1][415] = 16'b1111111111110010;
    assign weights1[1][416] = 16'b0000000000001110;
    assign weights1[1][417] = 16'b1111111111111010;
    assign weights1[1][418] = 16'b1111111111110100;
    assign weights1[1][419] = 16'b0000000000001000;
    assign weights1[1][420] = 16'b1111111111001000;
    assign weights1[1][421] = 16'b1111111110100110;
    assign weights1[1][422] = 16'b1111111110101010;
    assign weights1[1][423] = 16'b1111111110110001;
    assign weights1[1][424] = 16'b1111111111001010;
    assign weights1[1][425] = 16'b1111111111110010;
    assign weights1[1][426] = 16'b0000000000101101;
    assign weights1[1][427] = 16'b0000000000100010;
    assign weights1[1][428] = 16'b0000000000001001;
    assign weights1[1][429] = 16'b0000000000001111;
    assign weights1[1][430] = 16'b0000000000011101;
    assign weights1[1][431] = 16'b0000000000011001;
    assign weights1[1][432] = 16'b0000000000001110;
    assign weights1[1][433] = 16'b0000000000000000;
    assign weights1[1][434] = 16'b1111111111110111;
    assign weights1[1][435] = 16'b0000000000000111;
    assign weights1[1][436] = 16'b1111111111110110;
    assign weights1[1][437] = 16'b0000000000001001;
    assign weights1[1][438] = 16'b0000000000001011;
    assign weights1[1][439] = 16'b1111111111101001;
    assign weights1[1][440] = 16'b1111111111111101;
    assign weights1[1][441] = 16'b1111111111111000;
    assign weights1[1][442] = 16'b1111111111011100;
    assign weights1[1][443] = 16'b0000000000001011;
    assign weights1[1][444] = 16'b0000000000000000;
    assign weights1[1][445] = 16'b1111111111111011;
    assign weights1[1][446] = 16'b0000000000010000;
    assign weights1[1][447] = 16'b0000000000000001;
    assign weights1[1][448] = 16'b1111111111001010;
    assign weights1[1][449] = 16'b1111111110111000;
    assign weights1[1][450] = 16'b1111111110100110;
    assign weights1[1][451] = 16'b1111111101111101;
    assign weights1[1][452] = 16'b1111111101001001;
    assign weights1[1][453] = 16'b1111111101110000;
    assign weights1[1][454] = 16'b1111111110110001;
    assign weights1[1][455] = 16'b1111111111010100;
    assign weights1[1][456] = 16'b0000000000000100;
    assign weights1[1][457] = 16'b0000000000010010;
    assign weights1[1][458] = 16'b0000000000000100;
    assign weights1[1][459] = 16'b0000000001000000;
    assign weights1[1][460] = 16'b0000000000100110;
    assign weights1[1][461] = 16'b0000000000100010;
    assign weights1[1][462] = 16'b0000000000001001;
    assign weights1[1][463] = 16'b1111111111111111;
    assign weights1[1][464] = 16'b0000000000000010;
    assign weights1[1][465] = 16'b0000000000000001;
    assign weights1[1][466] = 16'b1111111111101100;
    assign weights1[1][467] = 16'b0000000000000010;
    assign weights1[1][468] = 16'b1111111111110010;
    assign weights1[1][469] = 16'b1111111111110100;
    assign weights1[1][470] = 16'b1111111111111101;
    assign weights1[1][471] = 16'b1111111111110000;
    assign weights1[1][472] = 16'b1111111111111011;
    assign weights1[1][473] = 16'b0000000000001101;
    assign weights1[1][474] = 16'b0000000000010011;
    assign weights1[1][475] = 16'b0000000000000101;
    assign weights1[1][476] = 16'b1111111111010001;
    assign weights1[1][477] = 16'b1111111110110100;
    assign weights1[1][478] = 16'b1111111110110111;
    assign weights1[1][479] = 16'b1111111110000010;
    assign weights1[1][480] = 16'b1111111101011001;
    assign weights1[1][481] = 16'b1111111100101010;
    assign weights1[1][482] = 16'b1111111011101011;
    assign weights1[1][483] = 16'b1111111100011111;
    assign weights1[1][484] = 16'b1111111101101101;
    assign weights1[1][485] = 16'b1111111110111100;
    assign weights1[1][486] = 16'b1111111111100010;
    assign weights1[1][487] = 16'b0000000000000100;
    assign weights1[1][488] = 16'b0000000000010100;
    assign weights1[1][489] = 16'b0000000000001101;
    assign weights1[1][490] = 16'b0000000000000101;
    assign weights1[1][491] = 16'b1111111111110011;
    assign weights1[1][492] = 16'b1111111111101100;
    assign weights1[1][493] = 16'b1111111111100000;
    assign weights1[1][494] = 16'b1111111111111000;
    assign weights1[1][495] = 16'b1111111111101100;
    assign weights1[1][496] = 16'b1111111111111000;
    assign weights1[1][497] = 16'b1111111111110010;
    assign weights1[1][498] = 16'b1111111111110100;
    assign weights1[1][499] = 16'b0000000000001001;
    assign weights1[1][500] = 16'b1111111111111011;
    assign weights1[1][501] = 16'b0000000000000101;
    assign weights1[1][502] = 16'b0000000000000010;
    assign weights1[1][503] = 16'b0000000000001010;
    assign weights1[1][504] = 16'b1111111111011010;
    assign weights1[1][505] = 16'b1111111111001011;
    assign weights1[1][506] = 16'b1111111111001010;
    assign weights1[1][507] = 16'b1111111110111001;
    assign weights1[1][508] = 16'b1111111110011011;
    assign weights1[1][509] = 16'b1111111101101101;
    assign weights1[1][510] = 16'b1111111101000001;
    assign weights1[1][511] = 16'b1111111100000110;
    assign weights1[1][512] = 16'b1111111010111000;
    assign weights1[1][513] = 16'b1111111010101000;
    assign weights1[1][514] = 16'b1111111010110000;
    assign weights1[1][515] = 16'b1111111011101101;
    assign weights1[1][516] = 16'b1111111101000000;
    assign weights1[1][517] = 16'b1111111101111010;
    assign weights1[1][518] = 16'b1111111110010111;
    assign weights1[1][519] = 16'b1111111111001100;
    assign weights1[1][520] = 16'b1111111111001011;
    assign weights1[1][521] = 16'b1111111111100101;
    assign weights1[1][522] = 16'b1111111111110110;
    assign weights1[1][523] = 16'b1111111111111001;
    assign weights1[1][524] = 16'b1111111111111000;
    assign weights1[1][525] = 16'b1111111111111010;
    assign weights1[1][526] = 16'b0000000000000010;
    assign weights1[1][527] = 16'b0000000000010010;
    assign weights1[1][528] = 16'b1111111111111011;
    assign weights1[1][529] = 16'b0000000000001011;
    assign weights1[1][530] = 16'b0000000000000011;
    assign weights1[1][531] = 16'b0000000000001010;
    assign weights1[1][532] = 16'b1111111111110110;
    assign weights1[1][533] = 16'b1111111111101111;
    assign weights1[1][534] = 16'b1111111111110000;
    assign weights1[1][535] = 16'b1111111111101111;
    assign weights1[1][536] = 16'b1111111111011010;
    assign weights1[1][537] = 16'b1111111111100101;
    assign weights1[1][538] = 16'b1111111111010101;
    assign weights1[1][539] = 16'b1111111110101110;
    assign weights1[1][540] = 16'b1111111101010110;
    assign weights1[1][541] = 16'b1111111100100110;
    assign weights1[1][542] = 16'b1111111100011100;
    assign weights1[1][543] = 16'b1111111101000011;
    assign weights1[1][544] = 16'b1111111101100010;
    assign weights1[1][545] = 16'b1111111110101010;
    assign weights1[1][546] = 16'b1111111110110110;
    assign weights1[1][547] = 16'b1111111110111010;
    assign weights1[1][548] = 16'b1111111111110010;
    assign weights1[1][549] = 16'b1111111111110100;
    assign weights1[1][550] = 16'b1111111111110111;
    assign weights1[1][551] = 16'b1111111111111100;
    assign weights1[1][552] = 16'b0000000000011000;
    assign weights1[1][553] = 16'b1111111111111000;
    assign weights1[1][554] = 16'b0000000000001010;
    assign weights1[1][555] = 16'b1111111111111010;
    assign weights1[1][556] = 16'b0000000000010110;
    assign weights1[1][557] = 16'b0000000000001000;
    assign weights1[1][558] = 16'b0000000000010010;
    assign weights1[1][559] = 16'b0000000000000110;
    assign weights1[1][560] = 16'b0000000000000010;
    assign weights1[1][561] = 16'b0000000000000110;
    assign weights1[1][562] = 16'b0000000000010000;
    assign weights1[1][563] = 16'b0000000000001110;
    assign weights1[1][564] = 16'b0000000000010100;
    assign weights1[1][565] = 16'b0000000000001110;
    assign weights1[1][566] = 16'b0000000000011000;
    assign weights1[1][567] = 16'b0000000000010011;
    assign weights1[1][568] = 16'b0000000000111110;
    assign weights1[1][569] = 16'b0000000000111010;
    assign weights1[1][570] = 16'b0000000000101000;
    assign weights1[1][571] = 16'b0000000000101001;
    assign weights1[1][572] = 16'b1111111111111001;
    assign weights1[1][573] = 16'b1111111111110010;
    assign weights1[1][574] = 16'b0000000000000101;
    assign weights1[1][575] = 16'b1111111111111011;
    assign weights1[1][576] = 16'b1111111111111100;
    assign weights1[1][577] = 16'b0000000000000101;
    assign weights1[1][578] = 16'b0000000000001011;
    assign weights1[1][579] = 16'b0000000000001111;
    assign weights1[1][580] = 16'b0000000000000011;
    assign weights1[1][581] = 16'b0000000000001001;
    assign weights1[1][582] = 16'b0000000000010011;
    assign weights1[1][583] = 16'b0000000000000001;
    assign weights1[1][584] = 16'b1111111111111110;
    assign weights1[1][585] = 16'b0000000000001001;
    assign weights1[1][586] = 16'b0000000000001111;
    assign weights1[1][587] = 16'b0000000000001011;
    assign weights1[1][588] = 16'b0000000000010101;
    assign weights1[1][589] = 16'b0000000000010011;
    assign weights1[1][590] = 16'b0000000000011100;
    assign weights1[1][591] = 16'b0000000000011111;
    assign weights1[1][592] = 16'b0000000000110010;
    assign weights1[1][593] = 16'b0000000001000101;
    assign weights1[1][594] = 16'b0000000001011010;
    assign weights1[1][595] = 16'b0000000001001111;
    assign weights1[1][596] = 16'b0000000001101100;
    assign weights1[1][597] = 16'b0000000001011101;
    assign weights1[1][598] = 16'b0000000001000011;
    assign weights1[1][599] = 16'b0000000000111111;
    assign weights1[1][600] = 16'b0000000000101000;
    assign weights1[1][601] = 16'b0000000000100101;
    assign weights1[1][602] = 16'b0000000000000111;
    assign weights1[1][603] = 16'b0000000000001000;
    assign weights1[1][604] = 16'b0000000000011010;
    assign weights1[1][605] = 16'b1111111111110111;
    assign weights1[1][606] = 16'b1111111111110110;
    assign weights1[1][607] = 16'b0000000000001101;
    assign weights1[1][608] = 16'b1111111111111000;
    assign weights1[1][609] = 16'b0000000000000010;
    assign weights1[1][610] = 16'b1111111111111000;
    assign weights1[1][611] = 16'b0000000000001010;
    assign weights1[1][612] = 16'b0000000000000111;
    assign weights1[1][613] = 16'b0000000000000011;
    assign weights1[1][614] = 16'b0000000000000101;
    assign weights1[1][615] = 16'b1111111111111100;
    assign weights1[1][616] = 16'b0000000000000111;
    assign weights1[1][617] = 16'b0000000000000111;
    assign weights1[1][618] = 16'b0000000000100001;
    assign weights1[1][619] = 16'b0000000000100001;
    assign weights1[1][620] = 16'b0000000000101011;
    assign weights1[1][621] = 16'b0000000000101010;
    assign weights1[1][622] = 16'b0000000000011010;
    assign weights1[1][623] = 16'b0000000001000101;
    assign weights1[1][624] = 16'b0000000000111011;
    assign weights1[1][625] = 16'b0000000000111000;
    assign weights1[1][626] = 16'b0000000000100110;
    assign weights1[1][627] = 16'b0000000000111100;
    assign weights1[1][628] = 16'b0000000000011011;
    assign weights1[1][629] = 16'b0000000000001110;
    assign weights1[1][630] = 16'b0000000000101100;
    assign weights1[1][631] = 16'b0000000000000101;
    assign weights1[1][632] = 16'b0000000000000101;
    assign weights1[1][633] = 16'b1111111111111000;
    assign weights1[1][634] = 16'b0000000000000110;
    assign weights1[1][635] = 16'b1111111111111101;
    assign weights1[1][636] = 16'b1111111111111011;
    assign weights1[1][637] = 16'b0000000000000000;
    assign weights1[1][638] = 16'b0000000000001101;
    assign weights1[1][639] = 16'b1111111111110110;
    assign weights1[1][640] = 16'b0000000000000100;
    assign weights1[1][641] = 16'b1111111111110101;
    assign weights1[1][642] = 16'b0000000000000100;
    assign weights1[1][643] = 16'b0000000000000010;
    assign weights1[1][644] = 16'b0000000000001001;
    assign weights1[1][645] = 16'b0000000000000101;
    assign weights1[1][646] = 16'b0000000000010001;
    assign weights1[1][647] = 16'b0000000000100001;
    assign weights1[1][648] = 16'b0000000000100011;
    assign weights1[1][649] = 16'b0000000001000001;
    assign weights1[1][650] = 16'b0000000000101111;
    assign weights1[1][651] = 16'b0000000000000100;
    assign weights1[1][652] = 16'b1111111111110111;
    assign weights1[1][653] = 16'b0000000000100000;
    assign weights1[1][654] = 16'b0000000000011011;
    assign weights1[1][655] = 16'b0000000000001000;
    assign weights1[1][656] = 16'b0000000000001100;
    assign weights1[1][657] = 16'b0000000000100011;
    assign weights1[1][658] = 16'b1111111111111011;
    assign weights1[1][659] = 16'b0000000000010011;
    assign weights1[1][660] = 16'b0000000000000101;
    assign weights1[1][661] = 16'b0000000000001011;
    assign weights1[1][662] = 16'b0000000000000111;
    assign weights1[1][663] = 16'b0000000000000011;
    assign weights1[1][664] = 16'b0000000000010010;
    assign weights1[1][665] = 16'b1111111111111010;
    assign weights1[1][666] = 16'b0000000000001000;
    assign weights1[1][667] = 16'b0000000000001110;
    assign weights1[1][668] = 16'b0000000000001011;
    assign weights1[1][669] = 16'b1111111111110110;
    assign weights1[1][670] = 16'b1111111111111011;
    assign weights1[1][671] = 16'b1111111111111110;
    assign weights1[1][672] = 16'b0000000000000000;
    assign weights1[1][673] = 16'b1111111111111100;
    assign weights1[1][674] = 16'b1111111111110010;
    assign weights1[1][675] = 16'b0000000000010111;
    assign weights1[1][676] = 16'b0000000000001011;
    assign weights1[1][677] = 16'b0000000000010010;
    assign weights1[1][678] = 16'b0000000000101000;
    assign weights1[1][679] = 16'b0000000000110110;
    assign weights1[1][680] = 16'b0000000000010100;
    assign weights1[1][681] = 16'b0000000000100000;
    assign weights1[1][682] = 16'b0000000000001100;
    assign weights1[1][683] = 16'b0000000000100010;
    assign weights1[1][684] = 16'b0000000000000001;
    assign weights1[1][685] = 16'b0000000000000011;
    assign weights1[1][686] = 16'b0000000000011011;
    assign weights1[1][687] = 16'b1111111111111110;
    assign weights1[1][688] = 16'b0000000000000000;
    assign weights1[1][689] = 16'b0000000000001110;
    assign weights1[1][690] = 16'b1111111111111110;
    assign weights1[1][691] = 16'b1111111111110110;
    assign weights1[1][692] = 16'b0000000000000101;
    assign weights1[1][693] = 16'b1111111111111001;
    assign weights1[1][694] = 16'b0000000000000001;
    assign weights1[1][695] = 16'b1111111111110110;
    assign weights1[1][696] = 16'b1111111111101110;
    assign weights1[1][697] = 16'b1111111111110111;
    assign weights1[1][698] = 16'b1111111111111110;
    assign weights1[1][699] = 16'b1111111111111100;
    assign weights1[1][700] = 16'b1111111111111100;
    assign weights1[1][701] = 16'b1111111111111110;
    assign weights1[1][702] = 16'b1111111111110110;
    assign weights1[1][703] = 16'b1111111111110001;
    assign weights1[1][704] = 16'b1111111111111010;
    assign weights1[1][705] = 16'b1111111111111010;
    assign weights1[1][706] = 16'b1111111111110010;
    assign weights1[1][707] = 16'b0000000000010010;
    assign weights1[1][708] = 16'b0000000000000010;
    assign weights1[1][709] = 16'b0000000000001111;
    assign weights1[1][710] = 16'b0000000000000111;
    assign weights1[1][711] = 16'b0000000000001011;
    assign weights1[1][712] = 16'b0000000000011000;
    assign weights1[1][713] = 16'b0000000000010010;
    assign weights1[1][714] = 16'b1111111111111100;
    assign weights1[1][715] = 16'b0000000000010100;
    assign weights1[1][716] = 16'b0000000000000001;
    assign weights1[1][717] = 16'b0000000000000101;
    assign weights1[1][718] = 16'b0000000000000011;
    assign weights1[1][719] = 16'b0000000000001001;
    assign weights1[1][720] = 16'b1111111111111111;
    assign weights1[1][721] = 16'b0000000000000001;
    assign weights1[1][722] = 16'b1111111111111110;
    assign weights1[1][723] = 16'b0000000000000000;
    assign weights1[1][724] = 16'b1111111111111100;
    assign weights1[1][725] = 16'b1111111111110011;
    assign weights1[1][726] = 16'b1111111111111111;
    assign weights1[1][727] = 16'b1111111111111100;
    assign weights1[1][728] = 16'b1111111111111101;
    assign weights1[1][729] = 16'b1111111111111101;
    assign weights1[1][730] = 16'b1111111111111100;
    assign weights1[1][731] = 16'b1111111111101111;
    assign weights1[1][732] = 16'b1111111111011110;
    assign weights1[1][733] = 16'b1111111111011101;
    assign weights1[1][734] = 16'b1111111111010111;
    assign weights1[1][735] = 16'b1111111111001111;
    assign weights1[1][736] = 16'b1111111111100000;
    assign weights1[1][737] = 16'b1111111111110101;
    assign weights1[1][738] = 16'b1111111111111011;
    assign weights1[1][739] = 16'b1111111111101001;
    assign weights1[1][740] = 16'b1111111111100111;
    assign weights1[1][741] = 16'b0000000000000011;
    assign weights1[1][742] = 16'b0000000000001011;
    assign weights1[1][743] = 16'b1111111111101111;
    assign weights1[1][744] = 16'b0000000000011010;
    assign weights1[1][745] = 16'b1111111111110100;
    assign weights1[1][746] = 16'b1111111111111010;
    assign weights1[1][747] = 16'b0000000000000110;
    assign weights1[1][748] = 16'b0000000000000111;
    assign weights1[1][749] = 16'b0000000000000000;
    assign weights1[1][750] = 16'b1111111111101110;
    assign weights1[1][751] = 16'b1111111111111011;
    assign weights1[1][752] = 16'b1111111111111010;
    assign weights1[1][753] = 16'b1111111111111110;
    assign weights1[1][754] = 16'b1111111111111100;
    assign weights1[1][755] = 16'b0000000000000000;
    assign weights1[1][756] = 16'b0000000000000000;
    assign weights1[1][757] = 16'b1111111111111111;
    assign weights1[1][758] = 16'b1111111111111001;
    assign weights1[1][759] = 16'b1111111111101110;
    assign weights1[1][760] = 16'b1111111111100101;
    assign weights1[1][761] = 16'b1111111111100001;
    assign weights1[1][762] = 16'b1111111111100110;
    assign weights1[1][763] = 16'b1111111111010010;
    assign weights1[1][764] = 16'b1111111111010000;
    assign weights1[1][765] = 16'b1111111111011011;
    assign weights1[1][766] = 16'b1111111111101111;
    assign weights1[1][767] = 16'b1111111111101010;
    assign weights1[1][768] = 16'b1111111111111100;
    assign weights1[1][769] = 16'b1111111111111000;
    assign weights1[1][770] = 16'b1111111111100001;
    assign weights1[1][771] = 16'b1111111111100110;
    assign weights1[1][772] = 16'b1111111111011111;
    assign weights1[1][773] = 16'b1111111111100101;
    assign weights1[1][774] = 16'b1111111111110000;
    assign weights1[1][775] = 16'b1111111111100010;
    assign weights1[1][776] = 16'b1111111111110001;
    assign weights1[1][777] = 16'b1111111111101101;
    assign weights1[1][778] = 16'b1111111111111000;
    assign weights1[1][779] = 16'b0000000000000011;
    assign weights1[1][780] = 16'b1111111111111111;
    assign weights1[1][781] = 16'b0000000000000001;
    assign weights1[1][782] = 16'b1111111111111101;
    assign weights1[1][783] = 16'b0000000000000000;
    assign weights1[2][0] = 16'b0000000000000000;
    assign weights1[2][1] = 16'b0000000000000000;
    assign weights1[2][2] = 16'b0000000000000000;
    assign weights1[2][3] = 16'b0000000000000000;
    assign weights1[2][4] = 16'b1111111111111110;
    assign weights1[2][5] = 16'b1111111111111111;
    assign weights1[2][6] = 16'b1111111111111000;
    assign weights1[2][7] = 16'b1111111111110101;
    assign weights1[2][8] = 16'b1111111111111001;
    assign weights1[2][9] = 16'b0000000000000110;
    assign weights1[2][10] = 16'b0000000000000100;
    assign weights1[2][11] = 16'b0000000000001101;
    assign weights1[2][12] = 16'b0000000000010000;
    assign weights1[2][13] = 16'b1111111111110101;
    assign weights1[2][14] = 16'b1111111111111111;
    assign weights1[2][15] = 16'b0000000000001100;
    assign weights1[2][16] = 16'b0000000000000010;
    assign weights1[2][17] = 16'b0000000000000010;
    assign weights1[2][18] = 16'b0000000000000010;
    assign weights1[2][19] = 16'b0000000000001000;
    assign weights1[2][20] = 16'b0000000000000001;
    assign weights1[2][21] = 16'b1111111111111101;
    assign weights1[2][22] = 16'b1111111111111100;
    assign weights1[2][23] = 16'b1111111111111111;
    assign weights1[2][24] = 16'b0000000000000000;
    assign weights1[2][25] = 16'b0000000000000001;
    assign weights1[2][26] = 16'b0000000000000000;
    assign weights1[2][27] = 16'b0000000000000000;
    assign weights1[2][28] = 16'b0000000000000000;
    assign weights1[2][29] = 16'b0000000000000000;
    assign weights1[2][30] = 16'b0000000000000000;
    assign weights1[2][31] = 16'b1111111111111111;
    assign weights1[2][32] = 16'b1111111111111001;
    assign weights1[2][33] = 16'b1111111111110101;
    assign weights1[2][34] = 16'b1111111111110101;
    assign weights1[2][35] = 16'b1111111111110000;
    assign weights1[2][36] = 16'b1111111111110110;
    assign weights1[2][37] = 16'b0000000000000101;
    assign weights1[2][38] = 16'b0000000000010000;
    assign weights1[2][39] = 16'b0000000000000111;
    assign weights1[2][40] = 16'b0000000000000010;
    assign weights1[2][41] = 16'b1111111111101100;
    assign weights1[2][42] = 16'b1111111111111001;
    assign weights1[2][43] = 16'b0000000000001101;
    assign weights1[2][44] = 16'b0000000000000010;
    assign weights1[2][45] = 16'b1111111111111101;
    assign weights1[2][46] = 16'b0000000000000101;
    assign weights1[2][47] = 16'b0000000000000011;
    assign weights1[2][48] = 16'b0000000000000011;
    assign weights1[2][49] = 16'b1111111111111000;
    assign weights1[2][50] = 16'b1111111111111001;
    assign weights1[2][51] = 16'b1111111111110111;
    assign weights1[2][52] = 16'b1111111111111011;
    assign weights1[2][53] = 16'b1111111111111101;
    assign weights1[2][54] = 16'b1111111111111110;
    assign weights1[2][55] = 16'b1111111111111111;
    assign weights1[2][56] = 16'b0000000000000000;
    assign weights1[2][57] = 16'b0000000000000000;
    assign weights1[2][58] = 16'b1111111111111111;
    assign weights1[2][59] = 16'b1111111111111010;
    assign weights1[2][60] = 16'b1111111111110100;
    assign weights1[2][61] = 16'b1111111111101101;
    assign weights1[2][62] = 16'b1111111111101001;
    assign weights1[2][63] = 16'b1111111111101010;
    assign weights1[2][64] = 16'b1111111111110110;
    assign weights1[2][65] = 16'b0000000000000100;
    assign weights1[2][66] = 16'b0000000000010111;
    assign weights1[2][67] = 16'b0000000000010000;
    assign weights1[2][68] = 16'b1111111111110100;
    assign weights1[2][69] = 16'b0000000000001100;
    assign weights1[2][70] = 16'b1111111111101111;
    assign weights1[2][71] = 16'b0000000000000010;
    assign weights1[2][72] = 16'b0000000000000011;
    assign weights1[2][73] = 16'b1111111111111011;
    assign weights1[2][74] = 16'b0000000000000010;
    assign weights1[2][75] = 16'b0000000000011101;
    assign weights1[2][76] = 16'b1111111111111100;
    assign weights1[2][77] = 16'b1111111111111001;
    assign weights1[2][78] = 16'b1111111111110111;
    assign weights1[2][79] = 16'b1111111111110101;
    assign weights1[2][80] = 16'b1111111111110100;
    assign weights1[2][81] = 16'b1111111111111101;
    assign weights1[2][82] = 16'b1111111111111111;
    assign weights1[2][83] = 16'b0000000000000000;
    assign weights1[2][84] = 16'b0000000000000000;
    assign weights1[2][85] = 16'b0000000000000000;
    assign weights1[2][86] = 16'b1111111111111001;
    assign weights1[2][87] = 16'b1111111111110100;
    assign weights1[2][88] = 16'b1111111111110010;
    assign weights1[2][89] = 16'b1111111111100110;
    assign weights1[2][90] = 16'b1111111111011100;
    assign weights1[2][91] = 16'b1111111111011100;
    assign weights1[2][92] = 16'b1111111111101001;
    assign weights1[2][93] = 16'b0000000000001010;
    assign weights1[2][94] = 16'b0000000000001100;
    assign weights1[2][95] = 16'b0000000000000101;
    assign weights1[2][96] = 16'b1111111111111011;
    assign weights1[2][97] = 16'b1111111111101101;
    assign weights1[2][98] = 16'b1111111111111110;
    assign weights1[2][99] = 16'b1111111111111100;
    assign weights1[2][100] = 16'b1111111111111010;
    assign weights1[2][101] = 16'b0000000000000100;
    assign weights1[2][102] = 16'b0000000000001110;
    assign weights1[2][103] = 16'b0000000000000000;
    assign weights1[2][104] = 16'b0000000000000101;
    assign weights1[2][105] = 16'b1111111111110011;
    assign weights1[2][106] = 16'b1111111111110010;
    assign weights1[2][107] = 16'b1111111111110100;
    assign weights1[2][108] = 16'b1111111111110101;
    assign weights1[2][109] = 16'b1111111111111101;
    assign weights1[2][110] = 16'b1111111111111111;
    assign weights1[2][111] = 16'b0000000000000000;
    assign weights1[2][112] = 16'b1111111111111110;
    assign weights1[2][113] = 16'b1111111111111100;
    assign weights1[2][114] = 16'b0000000000000000;
    assign weights1[2][115] = 16'b1111111111110001;
    assign weights1[2][116] = 16'b1111111111101100;
    assign weights1[2][117] = 16'b1111111111101000;
    assign weights1[2][118] = 16'b1111111111011001;
    assign weights1[2][119] = 16'b1111111111011001;
    assign weights1[2][120] = 16'b1111111111100101;
    assign weights1[2][121] = 16'b0000000000000101;
    assign weights1[2][122] = 16'b0000000000001001;
    assign weights1[2][123] = 16'b0000000000100111;
    assign weights1[2][124] = 16'b1111111111110101;
    assign weights1[2][125] = 16'b0000000000001001;
    assign weights1[2][126] = 16'b1111111111111100;
    assign weights1[2][127] = 16'b0000000000001000;
    assign weights1[2][128] = 16'b1111111111110011;
    assign weights1[2][129] = 16'b0000000000001010;
    assign weights1[2][130] = 16'b0000000000001000;
    assign weights1[2][131] = 16'b1111111111101000;
    assign weights1[2][132] = 16'b1111111111111101;
    assign weights1[2][133] = 16'b1111111111101111;
    assign weights1[2][134] = 16'b1111111111010111;
    assign weights1[2][135] = 16'b1111111111101111;
    assign weights1[2][136] = 16'b1111111111110101;
    assign weights1[2][137] = 16'b1111111111111011;
    assign weights1[2][138] = 16'b1111111111111111;
    assign weights1[2][139] = 16'b1111111111111111;
    assign weights1[2][140] = 16'b0000000000000000;
    assign weights1[2][141] = 16'b1111111111111100;
    assign weights1[2][142] = 16'b1111111111111100;
    assign weights1[2][143] = 16'b1111111111111110;
    assign weights1[2][144] = 16'b1111111111111101;
    assign weights1[2][145] = 16'b1111111111110111;
    assign weights1[2][146] = 16'b1111111111011101;
    assign weights1[2][147] = 16'b1111111111110010;
    assign weights1[2][148] = 16'b1111111111100000;
    assign weights1[2][149] = 16'b1111111111111110;
    assign weights1[2][150] = 16'b0000000000000101;
    assign weights1[2][151] = 16'b0000000000000111;
    assign weights1[2][152] = 16'b1111111111101001;
    assign weights1[2][153] = 16'b1111111111111101;
    assign weights1[2][154] = 16'b1111111111011100;
    assign weights1[2][155] = 16'b1111111111110100;
    assign weights1[2][156] = 16'b1111111111111001;
    assign weights1[2][157] = 16'b1111111111010000;
    assign weights1[2][158] = 16'b1111111111100111;
    assign weights1[2][159] = 16'b1111111111101011;
    assign weights1[2][160] = 16'b1111111111101110;
    assign weights1[2][161] = 16'b1111111111011001;
    assign weights1[2][162] = 16'b1111111111010000;
    assign weights1[2][163] = 16'b1111111111011100;
    assign weights1[2][164] = 16'b1111111111110100;
    assign weights1[2][165] = 16'b1111111111111011;
    assign weights1[2][166] = 16'b0000000000000100;
    assign weights1[2][167] = 16'b0000000000000010;
    assign weights1[2][168] = 16'b0000000000000011;
    assign weights1[2][169] = 16'b1111111111111110;
    assign weights1[2][170] = 16'b1111111111111110;
    assign weights1[2][171] = 16'b1111111111111100;
    assign weights1[2][172] = 16'b1111111111110010;
    assign weights1[2][173] = 16'b1111111111101111;
    assign weights1[2][174] = 16'b1111111111101000;
    assign weights1[2][175] = 16'b1111111111101000;
    assign weights1[2][176] = 16'b1111111111011111;
    assign weights1[2][177] = 16'b1111111111010001;
    assign weights1[2][178] = 16'b1111111111110010;
    assign weights1[2][179] = 16'b0000000000010001;
    assign weights1[2][180] = 16'b0000000000000101;
    assign weights1[2][181] = 16'b1111111111111110;
    assign weights1[2][182] = 16'b1111111111101001;
    assign weights1[2][183] = 16'b1111111111110010;
    assign weights1[2][184] = 16'b1111111111111000;
    assign weights1[2][185] = 16'b1111111111110001;
    assign weights1[2][186] = 16'b1111111111110000;
    assign weights1[2][187] = 16'b1111111111001100;
    assign weights1[2][188] = 16'b1111111111011111;
    assign weights1[2][189] = 16'b1111111111000111;
    assign weights1[2][190] = 16'b1111111111011100;
    assign weights1[2][191] = 16'b1111111111101011;
    assign weights1[2][192] = 16'b1111111111110001;
    assign weights1[2][193] = 16'b1111111111110001;
    assign weights1[2][194] = 16'b0000000000000001;
    assign weights1[2][195] = 16'b0000000000000001;
    assign weights1[2][196] = 16'b0000000000000100;
    assign weights1[2][197] = 16'b0000000000001001;
    assign weights1[2][198] = 16'b0000000000000101;
    assign weights1[2][199] = 16'b0000000000001000;
    assign weights1[2][200] = 16'b0000000000000001;
    assign weights1[2][201] = 16'b0000000000000000;
    assign weights1[2][202] = 16'b0000000000000000;
    assign weights1[2][203] = 16'b1111111111101000;
    assign weights1[2][204] = 16'b1111111111101010;
    assign weights1[2][205] = 16'b1111111111010110;
    assign weights1[2][206] = 16'b1111111111101000;
    assign weights1[2][207] = 16'b0000000000010010;
    assign weights1[2][208] = 16'b0000000000010011;
    assign weights1[2][209] = 16'b1111111111111110;
    assign weights1[2][210] = 16'b1111111111111110;
    assign weights1[2][211] = 16'b1111111111101011;
    assign weights1[2][212] = 16'b1111111111110101;
    assign weights1[2][213] = 16'b0000000000001100;
    assign weights1[2][214] = 16'b1111111111010110;
    assign weights1[2][215] = 16'b1111111111101011;
    assign weights1[2][216] = 16'b1111111111001011;
    assign weights1[2][217] = 16'b1111111111000110;
    assign weights1[2][218] = 16'b1111111111100110;
    assign weights1[2][219] = 16'b1111111111101110;
    assign weights1[2][220] = 16'b1111111111101000;
    assign weights1[2][221] = 16'b1111111111110010;
    assign weights1[2][222] = 16'b0000000000000001;
    assign weights1[2][223] = 16'b0000000000000010;
    assign weights1[2][224] = 16'b0000000000001011;
    assign weights1[2][225] = 16'b0000000000001001;
    assign weights1[2][226] = 16'b0000000000001000;
    assign weights1[2][227] = 16'b0000000000001101;
    assign weights1[2][228] = 16'b0000000000001000;
    assign weights1[2][229] = 16'b0000000000000101;
    assign weights1[2][230] = 16'b0000000000010001;
    assign weights1[2][231] = 16'b1111111111111010;
    assign weights1[2][232] = 16'b1111111111011110;
    assign weights1[2][233] = 16'b1111111111101001;
    assign weights1[2][234] = 16'b1111111111100111;
    assign weights1[2][235] = 16'b1111111111110110;
    assign weights1[2][236] = 16'b1111111111110111;
    assign weights1[2][237] = 16'b0000000000010000;
    assign weights1[2][238] = 16'b0000000000011010;
    assign weights1[2][239] = 16'b0000000000001101;
    assign weights1[2][240] = 16'b1111111111110110;
    assign weights1[2][241] = 16'b1111111111101001;
    assign weights1[2][242] = 16'b1111111110111000;
    assign weights1[2][243] = 16'b1111111111011111;
    assign weights1[2][244] = 16'b1111111110111011;
    assign weights1[2][245] = 16'b1111111110111010;
    assign weights1[2][246] = 16'b1111111111011111;
    assign weights1[2][247] = 16'b1111111111100010;
    assign weights1[2][248] = 16'b1111111111100111;
    assign weights1[2][249] = 16'b1111111111101101;
    assign weights1[2][250] = 16'b0000000000000001;
    assign weights1[2][251] = 16'b0000000000000101;
    assign weights1[2][252] = 16'b0000000000001001;
    assign weights1[2][253] = 16'b0000000000010000;
    assign weights1[2][254] = 16'b0000000000001101;
    assign weights1[2][255] = 16'b0000000000000111;
    assign weights1[2][256] = 16'b1111111111101110;
    assign weights1[2][257] = 16'b1111111111111111;
    assign weights1[2][258] = 16'b0000000000001010;
    assign weights1[2][259] = 16'b0000000000000100;
    assign weights1[2][260] = 16'b1111111111110001;
    assign weights1[2][261] = 16'b1111111111010101;
    assign weights1[2][262] = 16'b1111111111101001;
    assign weights1[2][263] = 16'b1111111111110100;
    assign weights1[2][264] = 16'b1111111111110000;
    assign weights1[2][265] = 16'b0000000000000001;
    assign weights1[2][266] = 16'b0000000000101100;
    assign weights1[2][267] = 16'b0000000000010111;
    assign weights1[2][268] = 16'b1111111111111110;
    assign weights1[2][269] = 16'b1111111111100100;
    assign weights1[2][270] = 16'b1111111111011010;
    assign weights1[2][271] = 16'b1111111111000011;
    assign weights1[2][272] = 16'b1111111110101110;
    assign weights1[2][273] = 16'b1111111111001100;
    assign weights1[2][274] = 16'b1111111111011001;
    assign weights1[2][275] = 16'b1111111111100011;
    assign weights1[2][276] = 16'b1111111111101000;
    assign weights1[2][277] = 16'b1111111111110011;
    assign weights1[2][278] = 16'b1111111111111101;
    assign weights1[2][279] = 16'b1111111111111111;
    assign weights1[2][280] = 16'b0000000000000111;
    assign weights1[2][281] = 16'b0000000000000111;
    assign weights1[2][282] = 16'b0000000000001001;
    assign weights1[2][283] = 16'b0000000000000100;
    assign weights1[2][284] = 16'b1111111111111101;
    assign weights1[2][285] = 16'b1111111111110010;
    assign weights1[2][286] = 16'b1111111111110010;
    assign weights1[2][287] = 16'b1111111111110111;
    assign weights1[2][288] = 16'b0000000000001001;
    assign weights1[2][289] = 16'b1111111111010110;
    assign weights1[2][290] = 16'b1111111111100000;
    assign weights1[2][291] = 16'b1111111111100101;
    assign weights1[2][292] = 16'b0000000000000000;
    assign weights1[2][293] = 16'b0000000000010101;
    assign weights1[2][294] = 16'b0000000000100101;
    assign weights1[2][295] = 16'b0000000001010010;
    assign weights1[2][296] = 16'b0000000000000111;
    assign weights1[2][297] = 16'b1111111111101111;
    assign weights1[2][298] = 16'b1111111111001001;
    assign weights1[2][299] = 16'b1111111110010110;
    assign weights1[2][300] = 16'b1111111110111011;
    assign weights1[2][301] = 16'b1111111111010001;
    assign weights1[2][302] = 16'b1111111111100100;
    assign weights1[2][303] = 16'b1111111111100001;
    assign weights1[2][304] = 16'b1111111111110100;
    assign weights1[2][305] = 16'b1111111111110110;
    assign weights1[2][306] = 16'b1111111111111000;
    assign weights1[2][307] = 16'b1111111111111111;
    assign weights1[2][308] = 16'b0000000000001100;
    assign weights1[2][309] = 16'b0000000000000010;
    assign weights1[2][310] = 16'b0000000000001001;
    assign weights1[2][311] = 16'b1111111111110110;
    assign weights1[2][312] = 16'b0000000000000011;
    assign weights1[2][313] = 16'b0000000000001111;
    assign weights1[2][314] = 16'b1111111111110011;
    assign weights1[2][315] = 16'b1111111111101111;
    assign weights1[2][316] = 16'b0000000000010010;
    assign weights1[2][317] = 16'b1111111111100000;
    assign weights1[2][318] = 16'b1111111111001111;
    assign weights1[2][319] = 16'b1111111111010000;
    assign weights1[2][320] = 16'b1111111111100110;
    assign weights1[2][321] = 16'b0000000000010011;
    assign weights1[2][322] = 16'b0000000000111010;
    assign weights1[2][323] = 16'b0000000000011010;
    assign weights1[2][324] = 16'b0000000000010010;
    assign weights1[2][325] = 16'b0000000000000101;
    assign weights1[2][326] = 16'b1111111110011001;
    assign weights1[2][327] = 16'b1111111110101111;
    assign weights1[2][328] = 16'b1111111110111110;
    assign weights1[2][329] = 16'b1111111111010100;
    assign weights1[2][330] = 16'b1111111111011011;
    assign weights1[2][331] = 16'b1111111111101010;
    assign weights1[2][332] = 16'b1111111111101101;
    assign weights1[2][333] = 16'b1111111111110001;
    assign weights1[2][334] = 16'b1111111111110101;
    assign weights1[2][335] = 16'b1111111111111100;
    assign weights1[2][336] = 16'b0000000000001001;
    assign weights1[2][337] = 16'b0000000000000110;
    assign weights1[2][338] = 16'b0000000000000110;
    assign weights1[2][339] = 16'b0000000000001010;
    assign weights1[2][340] = 16'b0000000000001101;
    assign weights1[2][341] = 16'b0000000000011000;
    assign weights1[2][342] = 16'b1111111111111110;
    assign weights1[2][343] = 16'b1111111111100010;
    assign weights1[2][344] = 16'b1111111111101110;
    assign weights1[2][345] = 16'b1111111111110110;
    assign weights1[2][346] = 16'b1111111111001010;
    assign weights1[2][347] = 16'b1111111111010110;
    assign weights1[2][348] = 16'b0000000000011000;
    assign weights1[2][349] = 16'b0000000000011010;
    assign weights1[2][350] = 16'b0000000000101110;
    assign weights1[2][351] = 16'b0000000000010000;
    assign weights1[2][352] = 16'b0000000000011000;
    assign weights1[2][353] = 16'b0000000000000001;
    assign weights1[2][354] = 16'b1111111110111110;
    assign weights1[2][355] = 16'b1111111110011001;
    assign weights1[2][356] = 16'b1111111110110111;
    assign weights1[2][357] = 16'b1111111111011010;
    assign weights1[2][358] = 16'b1111111111011101;
    assign weights1[2][359] = 16'b1111111111110001;
    assign weights1[2][360] = 16'b1111111111100100;
    assign weights1[2][361] = 16'b1111111111101111;
    assign weights1[2][362] = 16'b0000000000000000;
    assign weights1[2][363] = 16'b1111111111111111;
    assign weights1[2][364] = 16'b1111111111111111;
    assign weights1[2][365] = 16'b0000000000000100;
    assign weights1[2][366] = 16'b0000000000000100;
    assign weights1[2][367] = 16'b1111111111110110;
    assign weights1[2][368] = 16'b0000000000000000;
    assign weights1[2][369] = 16'b1111111111111110;
    assign weights1[2][370] = 16'b1111111111101110;
    assign weights1[2][371] = 16'b1111111111100101;
    assign weights1[2][372] = 16'b1111111111011111;
    assign weights1[2][373] = 16'b1111111111000000;
    assign weights1[2][374] = 16'b1111111110101010;
    assign weights1[2][375] = 16'b1111111111001110;
    assign weights1[2][376] = 16'b0000000000100011;
    assign weights1[2][377] = 16'b1111111111111000;
    assign weights1[2][378] = 16'b0000000000101010;
    assign weights1[2][379] = 16'b0000000000011010;
    assign weights1[2][380] = 16'b0000000000001101;
    assign weights1[2][381] = 16'b1111111111110000;
    assign weights1[2][382] = 16'b1111111110111001;
    assign weights1[2][383] = 16'b1111111110110100;
    assign weights1[2][384] = 16'b1111111110111111;
    assign weights1[2][385] = 16'b1111111111001111;
    assign weights1[2][386] = 16'b1111111111011110;
    assign weights1[2][387] = 16'b1111111111101011;
    assign weights1[2][388] = 16'b1111111111101011;
    assign weights1[2][389] = 16'b1111111111110011;
    assign weights1[2][390] = 16'b1111111111111110;
    assign weights1[2][391] = 16'b0000000000000001;
    assign weights1[2][392] = 16'b1111111111111010;
    assign weights1[2][393] = 16'b1111111111111000;
    assign weights1[2][394] = 16'b1111111111111101;
    assign weights1[2][395] = 16'b1111111111111010;
    assign weights1[2][396] = 16'b0000000000000101;
    assign weights1[2][397] = 16'b1111111111110110;
    assign weights1[2][398] = 16'b1111111111110010;
    assign weights1[2][399] = 16'b1111111111010100;
    assign weights1[2][400] = 16'b1111111110110110;
    assign weights1[2][401] = 16'b1111111110101111;
    assign weights1[2][402] = 16'b1111111111001101;
    assign weights1[2][403] = 16'b1111111111011000;
    assign weights1[2][404] = 16'b1111111111110101;
    assign weights1[2][405] = 16'b1111111111111111;
    assign weights1[2][406] = 16'b0000000000011110;
    assign weights1[2][407] = 16'b0000000000010100;
    assign weights1[2][408] = 16'b0000000000010110;
    assign weights1[2][409] = 16'b1111111111100110;
    assign weights1[2][410] = 16'b1111111111001111;
    assign weights1[2][411] = 16'b1111111110111101;
    assign weights1[2][412] = 16'b1111111110111001;
    assign weights1[2][413] = 16'b1111111111001010;
    assign weights1[2][414] = 16'b1111111111011011;
    assign weights1[2][415] = 16'b1111111111011011;
    assign weights1[2][416] = 16'b1111111111101101;
    assign weights1[2][417] = 16'b1111111111110111;
    assign weights1[2][418] = 16'b0000000000000110;
    assign weights1[2][419] = 16'b1111111111110111;
    assign weights1[2][420] = 16'b1111111111111101;
    assign weights1[2][421] = 16'b0000000000000001;
    assign weights1[2][422] = 16'b1111111111111100;
    assign weights1[2][423] = 16'b1111111111110110;
    assign weights1[2][424] = 16'b1111111111110111;
    assign weights1[2][425] = 16'b1111111111101101;
    assign weights1[2][426] = 16'b1111111111011100;
    assign weights1[2][427] = 16'b1111111111000110;
    assign weights1[2][428] = 16'b1111111110101111;
    assign weights1[2][429] = 16'b1111111111001000;
    assign weights1[2][430] = 16'b1111111110101100;
    assign weights1[2][431] = 16'b1111111111101100;
    assign weights1[2][432] = 16'b1111111111110101;
    assign weights1[2][433] = 16'b0000000000100010;
    assign weights1[2][434] = 16'b0000000000001101;
    assign weights1[2][435] = 16'b0000000000001001;
    assign weights1[2][436] = 16'b1111111111101001;
    assign weights1[2][437] = 16'b1111111111010110;
    assign weights1[2][438] = 16'b1111111111001011;
    assign weights1[2][439] = 16'b1111111110010100;
    assign weights1[2][440] = 16'b1111111110100101;
    assign weights1[2][441] = 16'b1111111111001011;
    assign weights1[2][442] = 16'b1111111111100010;
    assign weights1[2][443] = 16'b1111111111100011;
    assign weights1[2][444] = 16'b1111111111110011;
    assign weights1[2][445] = 16'b0000000000000010;
    assign weights1[2][446] = 16'b1111111111111001;
    assign weights1[2][447] = 16'b1111111111111000;
    assign weights1[2][448] = 16'b1111111111111010;
    assign weights1[2][449] = 16'b1111111111111000;
    assign weights1[2][450] = 16'b1111111111111001;
    assign weights1[2][451] = 16'b1111111111110001;
    assign weights1[2][452] = 16'b1111111111100000;
    assign weights1[2][453] = 16'b1111111111010100;
    assign weights1[2][454] = 16'b1111111111000010;
    assign weights1[2][455] = 16'b1111111111000101;
    assign weights1[2][456] = 16'b1111111111000100;
    assign weights1[2][457] = 16'b1111111111101100;
    assign weights1[2][458] = 16'b1111111111011011;
    assign weights1[2][459] = 16'b1111111111110100;
    assign weights1[2][460] = 16'b0000000000000110;
    assign weights1[2][461] = 16'b1111111111111000;
    assign weights1[2][462] = 16'b0000000000010011;
    assign weights1[2][463] = 16'b1111111111110001;
    assign weights1[2][464] = 16'b1111111111110011;
    assign weights1[2][465] = 16'b1111111111001001;
    assign weights1[2][466] = 16'b1111111111101100;
    assign weights1[2][467] = 16'b1111111110110011;
    assign weights1[2][468] = 16'b1111111110110010;
    assign weights1[2][469] = 16'b1111111111011001;
    assign weights1[2][470] = 16'b1111111111100000;
    assign weights1[2][471] = 16'b1111111111101110;
    assign weights1[2][472] = 16'b1111111111110100;
    assign weights1[2][473] = 16'b1111111111111001;
    assign weights1[2][474] = 16'b1111111111111111;
    assign weights1[2][475] = 16'b0000000000000001;
    assign weights1[2][476] = 16'b1111111111111101;
    assign weights1[2][477] = 16'b1111111111111011;
    assign weights1[2][478] = 16'b1111111111101111;
    assign weights1[2][479] = 16'b1111111111011001;
    assign weights1[2][480] = 16'b1111111111010101;
    assign weights1[2][481] = 16'b1111111111000111;
    assign weights1[2][482] = 16'b1111111111100010;
    assign weights1[2][483] = 16'b1111111111011100;
    assign weights1[2][484] = 16'b1111111111110011;
    assign weights1[2][485] = 16'b1111111111101100;
    assign weights1[2][486] = 16'b1111111111110110;
    assign weights1[2][487] = 16'b0000000000000101;
    assign weights1[2][488] = 16'b1111111111111000;
    assign weights1[2][489] = 16'b0000000000011101;
    assign weights1[2][490] = 16'b0000000000011001;
    assign weights1[2][491] = 16'b1111111111101011;
    assign weights1[2][492] = 16'b1111111111110110;
    assign weights1[2][493] = 16'b1111111111011010;
    assign weights1[2][494] = 16'b1111111110111111;
    assign weights1[2][495] = 16'b1111111110110011;
    assign weights1[2][496] = 16'b1111111111100011;
    assign weights1[2][497] = 16'b1111111111011111;
    assign weights1[2][498] = 16'b1111111111101101;
    assign weights1[2][499] = 16'b0000000000000001;
    assign weights1[2][500] = 16'b0000000000000001;
    assign weights1[2][501] = 16'b1111111111110000;
    assign weights1[2][502] = 16'b1111111111111101;
    assign weights1[2][503] = 16'b1111111111111011;
    assign weights1[2][504] = 16'b0000000000000001;
    assign weights1[2][505] = 16'b1111111111110010;
    assign weights1[2][506] = 16'b1111111111101001;
    assign weights1[2][507] = 16'b1111111111010010;
    assign weights1[2][508] = 16'b1111111111011010;
    assign weights1[2][509] = 16'b1111111111011111;
    assign weights1[2][510] = 16'b1111111111011111;
    assign weights1[2][511] = 16'b0000000000000010;
    assign weights1[2][512] = 16'b1111111111111010;
    assign weights1[2][513] = 16'b0000000000001111;
    assign weights1[2][514] = 16'b1111111111110000;
    assign weights1[2][515] = 16'b1111111111101100;
    assign weights1[2][516] = 16'b1111111111100110;
    assign weights1[2][517] = 16'b0000000000010100;
    assign weights1[2][518] = 16'b0000000000010100;
    assign weights1[2][519] = 16'b0000000000010010;
    assign weights1[2][520] = 16'b1111111111100000;
    assign weights1[2][521] = 16'b0000000000000010;
    assign weights1[2][522] = 16'b0000000000000011;
    assign weights1[2][523] = 16'b0000000000000001;
    assign weights1[2][524] = 16'b0000000000100100;
    assign weights1[2][525] = 16'b1111111111111010;
    assign weights1[2][526] = 16'b0000000000000101;
    assign weights1[2][527] = 16'b0000000000100011;
    assign weights1[2][528] = 16'b0000000000010110;
    assign weights1[2][529] = 16'b0000000000000001;
    assign weights1[2][530] = 16'b0000000000000001;
    assign weights1[2][531] = 16'b0000000000000110;
    assign weights1[2][532] = 16'b1111111111111100;
    assign weights1[2][533] = 16'b1111111111110100;
    assign weights1[2][534] = 16'b1111111111110000;
    assign weights1[2][535] = 16'b1111111111011000;
    assign weights1[2][536] = 16'b1111111111100100;
    assign weights1[2][537] = 16'b1111111111101011;
    assign weights1[2][538] = 16'b1111111111111101;
    assign weights1[2][539] = 16'b1111111111110111;
    assign weights1[2][540] = 16'b1111111111111100;
    assign weights1[2][541] = 16'b0000000000011100;
    assign weights1[2][542] = 16'b0000000000001110;
    assign weights1[2][543] = 16'b1111111111111101;
    assign weights1[2][544] = 16'b0000000000010000;
    assign weights1[2][545] = 16'b0000000000011101;
    assign weights1[2][546] = 16'b0000000000011101;
    assign weights1[2][547] = 16'b0000000000000111;
    assign weights1[2][548] = 16'b0000000000011011;
    assign weights1[2][549] = 16'b1111111111110111;
    assign weights1[2][550] = 16'b0000000000011101;
    assign weights1[2][551] = 16'b0000000000010101;
    assign weights1[2][552] = 16'b0000000000110000;
    assign weights1[2][553] = 16'b0000000000001001;
    assign weights1[2][554] = 16'b0000000000000001;
    assign weights1[2][555] = 16'b0000000000000001;
    assign weights1[2][556] = 16'b0000000000010001;
    assign weights1[2][557] = 16'b0000000000010111;
    assign weights1[2][558] = 16'b0000000000000111;
    assign weights1[2][559] = 16'b0000000000000110;
    assign weights1[2][560] = 16'b1111111111111001;
    assign weights1[2][561] = 16'b1111111111111000;
    assign weights1[2][562] = 16'b1111111111101100;
    assign weights1[2][563] = 16'b1111111111100010;
    assign weights1[2][564] = 16'b1111111111100000;
    assign weights1[2][565] = 16'b1111111111011010;
    assign weights1[2][566] = 16'b0000000000001001;
    assign weights1[2][567] = 16'b0000000000001101;
    assign weights1[2][568] = 16'b0000000000011111;
    assign weights1[2][569] = 16'b0000000000011001;
    assign weights1[2][570] = 16'b0000000000000100;
    assign weights1[2][571] = 16'b0000000000101001;
    assign weights1[2][572] = 16'b0000000000011101;
    assign weights1[2][573] = 16'b0000000000000011;
    assign weights1[2][574] = 16'b0000000000011110;
    assign weights1[2][575] = 16'b0000000000011100;
    assign weights1[2][576] = 16'b0000000000000110;
    assign weights1[2][577] = 16'b0000000000100100;
    assign weights1[2][578] = 16'b0000000001000010;
    assign weights1[2][579] = 16'b0000000000101010;
    assign weights1[2][580] = 16'b0000000000011101;
    assign weights1[2][581] = 16'b0000000000010101;
    assign weights1[2][582] = 16'b0000000000010000;
    assign weights1[2][583] = 16'b0000000000001110;
    assign weights1[2][584] = 16'b0000000000010110;
    assign weights1[2][585] = 16'b0000000000000110;
    assign weights1[2][586] = 16'b0000000000000111;
    assign weights1[2][587] = 16'b0000000000000010;
    assign weights1[2][588] = 16'b1111111111111000;
    assign weights1[2][589] = 16'b1111111111110001;
    assign weights1[2][590] = 16'b1111111111110001;
    assign weights1[2][591] = 16'b1111111111101001;
    assign weights1[2][592] = 16'b1111111111101011;
    assign weights1[2][593] = 16'b1111111111111001;
    assign weights1[2][594] = 16'b1111111111111100;
    assign weights1[2][595] = 16'b0000000000001100;
    assign weights1[2][596] = 16'b0000000000001011;
    assign weights1[2][597] = 16'b0000000000001111;
    assign weights1[2][598] = 16'b0000000000011000;
    assign weights1[2][599] = 16'b0000000000001011;
    assign weights1[2][600] = 16'b1111111111100110;
    assign weights1[2][601] = 16'b0000000000001000;
    assign weights1[2][602] = 16'b1111111111111111;
    assign weights1[2][603] = 16'b0000000000010111;
    assign weights1[2][604] = 16'b0000000000001101;
    assign weights1[2][605] = 16'b0000000000011101;
    assign weights1[2][606] = 16'b0000000000101001;
    assign weights1[2][607] = 16'b0000000000011001;
    assign weights1[2][608] = 16'b0000000000100001;
    assign weights1[2][609] = 16'b0000000000001001;
    assign weights1[2][610] = 16'b0000000000000101;
    assign weights1[2][611] = 16'b0000000000001111;
    assign weights1[2][612] = 16'b0000000000001000;
    assign weights1[2][613] = 16'b0000000000001000;
    assign weights1[2][614] = 16'b0000000000000101;
    assign weights1[2][615] = 16'b0000000000000100;
    assign weights1[2][616] = 16'b1111111111111100;
    assign weights1[2][617] = 16'b0000000000000000;
    assign weights1[2][618] = 16'b1111111111111100;
    assign weights1[2][619] = 16'b1111111111111010;
    assign weights1[2][620] = 16'b1111111111111111;
    assign weights1[2][621] = 16'b1111111111111111;
    assign weights1[2][622] = 16'b1111111111111001;
    assign weights1[2][623] = 16'b0000000000000111;
    assign weights1[2][624] = 16'b0000000000101001;
    assign weights1[2][625] = 16'b0000000000011001;
    assign weights1[2][626] = 16'b0000000000011000;
    assign weights1[2][627] = 16'b1111111111101000;
    assign weights1[2][628] = 16'b1111111111110000;
    assign weights1[2][629] = 16'b1111111111001101;
    assign weights1[2][630] = 16'b1111111111111101;
    assign weights1[2][631] = 16'b1111111111101110;
    assign weights1[2][632] = 16'b0000000000001011;
    assign weights1[2][633] = 16'b0000000000000111;
    assign weights1[2][634] = 16'b0000000000110000;
    assign weights1[2][635] = 16'b0000000000100011;
    assign weights1[2][636] = 16'b0000000000011110;
    assign weights1[2][637] = 16'b0000000000100001;
    assign weights1[2][638] = 16'b0000000000010101;
    assign weights1[2][639] = 16'b0000000000000010;
    assign weights1[2][640] = 16'b0000000000000110;
    assign weights1[2][641] = 16'b0000000000001001;
    assign weights1[2][642] = 16'b0000000000000101;
    assign weights1[2][643] = 16'b0000000000000011;
    assign weights1[2][644] = 16'b1111111111111110;
    assign weights1[2][645] = 16'b0000000000000111;
    assign weights1[2][646] = 16'b0000000000001000;
    assign weights1[2][647] = 16'b0000000000000110;
    assign weights1[2][648] = 16'b0000000000010101;
    assign weights1[2][649] = 16'b0000000000000101;
    assign weights1[2][650] = 16'b0000000000000101;
    assign weights1[2][651] = 16'b0000000000011101;
    assign weights1[2][652] = 16'b0000000000011110;
    assign weights1[2][653] = 16'b0000000000000000;
    assign weights1[2][654] = 16'b0000000000000010;
    assign weights1[2][655] = 16'b0000000000011110;
    assign weights1[2][656] = 16'b0000000000001010;
    assign weights1[2][657] = 16'b1111111111100011;
    assign weights1[2][658] = 16'b1111111111110101;
    assign weights1[2][659] = 16'b1111111111111110;
    assign weights1[2][660] = 16'b1111111111101110;
    assign weights1[2][661] = 16'b0000000000010010;
    assign weights1[2][662] = 16'b1111111111110111;
    assign weights1[2][663] = 16'b0000000000001000;
    assign weights1[2][664] = 16'b0000000000001110;
    assign weights1[2][665] = 16'b0000000000000111;
    assign weights1[2][666] = 16'b0000000000001111;
    assign weights1[2][667] = 16'b0000000000000101;
    assign weights1[2][668] = 16'b0000000000000111;
    assign weights1[2][669] = 16'b0000000000000101;
    assign weights1[2][670] = 16'b0000000000001000;
    assign weights1[2][671] = 16'b0000000000000100;
    assign weights1[2][672] = 16'b0000000000000000;
    assign weights1[2][673] = 16'b0000000000000001;
    assign weights1[2][674] = 16'b0000000000000110;
    assign weights1[2][675] = 16'b0000000000000101;
    assign weights1[2][676] = 16'b0000000000010010;
    assign weights1[2][677] = 16'b1111111111111111;
    assign weights1[2][678] = 16'b0000000000001111;
    assign weights1[2][679] = 16'b0000000000010001;
    assign weights1[2][680] = 16'b0000000000010010;
    assign weights1[2][681] = 16'b0000000000000111;
    assign weights1[2][682] = 16'b0000000000001110;
    assign weights1[2][683] = 16'b0000000000000011;
    assign weights1[2][684] = 16'b1111111111100111;
    assign weights1[2][685] = 16'b1111111111101000;
    assign weights1[2][686] = 16'b1111111111011001;
    assign weights1[2][687] = 16'b1111111111111101;
    assign weights1[2][688] = 16'b1111111111000100;
    assign weights1[2][689] = 16'b1111111111101101;
    assign weights1[2][690] = 16'b1111111111100011;
    assign weights1[2][691] = 16'b1111111111110101;
    assign weights1[2][692] = 16'b1111111111111100;
    assign weights1[2][693] = 16'b0000000000001000;
    assign weights1[2][694] = 16'b0000000000000110;
    assign weights1[2][695] = 16'b0000000000000100;
    assign weights1[2][696] = 16'b0000000000000100;
    assign weights1[2][697] = 16'b0000000000000001;
    assign weights1[2][698] = 16'b0000000000000011;
    assign weights1[2][699] = 16'b1111111111111111;
    assign weights1[2][700] = 16'b0000000000000100;
    assign weights1[2][701] = 16'b0000000000000101;
    assign weights1[2][702] = 16'b0000000000000100;
    assign weights1[2][703] = 16'b0000000000000010;
    assign weights1[2][704] = 16'b0000000000010111;
    assign weights1[2][705] = 16'b0000000000010001;
    assign weights1[2][706] = 16'b0000000000011100;
    assign weights1[2][707] = 16'b0000000000000111;
    assign weights1[2][708] = 16'b0000000000010001;
    assign weights1[2][709] = 16'b1111111111111011;
    assign weights1[2][710] = 16'b1111111111111001;
    assign weights1[2][711] = 16'b1111111111111100;
    assign weights1[2][712] = 16'b1111111111110101;
    assign weights1[2][713] = 16'b1111111111101111;
    assign weights1[2][714] = 16'b1111111111111000;
    assign weights1[2][715] = 16'b1111111111100001;
    assign weights1[2][716] = 16'b1111111111111110;
    assign weights1[2][717] = 16'b0000000000000011;
    assign weights1[2][718] = 16'b1111111111110110;
    assign weights1[2][719] = 16'b1111111111111001;
    assign weights1[2][720] = 16'b1111111111111000;
    assign weights1[2][721] = 16'b1111111111111110;
    assign weights1[2][722] = 16'b1111111111111101;
    assign weights1[2][723] = 16'b1111111111111100;
    assign weights1[2][724] = 16'b0000000000000010;
    assign weights1[2][725] = 16'b1111111111111111;
    assign weights1[2][726] = 16'b1111111111111111;
    assign weights1[2][727] = 16'b1111111111111111;
    assign weights1[2][728] = 16'b0000000000000100;
    assign weights1[2][729] = 16'b0000000000000110;
    assign weights1[2][730] = 16'b0000000000000011;
    assign weights1[2][731] = 16'b0000000000000000;
    assign weights1[2][732] = 16'b0000000000001010;
    assign weights1[2][733] = 16'b0000000000000111;
    assign weights1[2][734] = 16'b0000000000000010;
    assign weights1[2][735] = 16'b0000000000001110;
    assign weights1[2][736] = 16'b1111111111111100;
    assign weights1[2][737] = 16'b0000000000000001;
    assign weights1[2][738] = 16'b0000000000000010;
    assign weights1[2][739] = 16'b1111111111111110;
    assign weights1[2][740] = 16'b0000000000001110;
    assign weights1[2][741] = 16'b1111111111111011;
    assign weights1[2][742] = 16'b1111111111110100;
    assign weights1[2][743] = 16'b1111111111110010;
    assign weights1[2][744] = 16'b0000000000000010;
    assign weights1[2][745] = 16'b0000000000000001;
    assign weights1[2][746] = 16'b1111111111101100;
    assign weights1[2][747] = 16'b1111111111101000;
    assign weights1[2][748] = 16'b1111111111101110;
    assign weights1[2][749] = 16'b1111111111111000;
    assign weights1[2][750] = 16'b1111111111111111;
    assign weights1[2][751] = 16'b0000000000000000;
    assign weights1[2][752] = 16'b1111111111111110;
    assign weights1[2][753] = 16'b1111111111111110;
    assign weights1[2][754] = 16'b0000000000000000;
    assign weights1[2][755] = 16'b0000000000000000;
    assign weights1[2][756] = 16'b1111111111111111;
    assign weights1[2][757] = 16'b0000000000000001;
    assign weights1[2][758] = 16'b0000000000000001;
    assign weights1[2][759] = 16'b0000000000000001;
    assign weights1[2][760] = 16'b0000000000000111;
    assign weights1[2][761] = 16'b0000000000001101;
    assign weights1[2][762] = 16'b0000000000000100;
    assign weights1[2][763] = 16'b0000000000000100;
    assign weights1[2][764] = 16'b0000000000001100;
    assign weights1[2][765] = 16'b0000000000000000;
    assign weights1[2][766] = 16'b1111111111111000;
    assign weights1[2][767] = 16'b1111111111101001;
    assign weights1[2][768] = 16'b1111111111110001;
    assign weights1[2][769] = 16'b1111111111101111;
    assign weights1[2][770] = 16'b1111111111101010;
    assign weights1[2][771] = 16'b1111111111101010;
    assign weights1[2][772] = 16'b1111111111101101;
    assign weights1[2][773] = 16'b1111111111101011;
    assign weights1[2][774] = 16'b1111111111101010;
    assign weights1[2][775] = 16'b1111111111101110;
    assign weights1[2][776] = 16'b1111111111101001;
    assign weights1[2][777] = 16'b1111111111111011;
    assign weights1[2][778] = 16'b1111111111110111;
    assign weights1[2][779] = 16'b1111111111110110;
    assign weights1[2][780] = 16'b1111111111111111;
    assign weights1[2][781] = 16'b1111111111111101;
    assign weights1[2][782] = 16'b0000000000000000;
    assign weights1[2][783] = 16'b0000000000000000;
    assign weights1[3][0] = 16'b1111111111111111;
    assign weights1[3][1] = 16'b1111111111111111;
    assign weights1[3][2] = 16'b1111111111111111;
    assign weights1[3][3] = 16'b1111111111111111;
    assign weights1[3][4] = 16'b1111111111111111;
    assign weights1[3][5] = 16'b0000000000000000;
    assign weights1[3][6] = 16'b1111111111111010;
    assign weights1[3][7] = 16'b1111111111111110;
    assign weights1[3][8] = 16'b1111111111111111;
    assign weights1[3][9] = 16'b1111111111110100;
    assign weights1[3][10] = 16'b1111111111101011;
    assign weights1[3][11] = 16'b1111111111100110;
    assign weights1[3][12] = 16'b1111111111100001;
    assign weights1[3][13] = 16'b1111111111100010;
    assign weights1[3][14] = 16'b1111111111011111;
    assign weights1[3][15] = 16'b1111111111101011;
    assign weights1[3][16] = 16'b0000000000001101;
    assign weights1[3][17] = 16'b0000000000010101;
    assign weights1[3][18] = 16'b0000000000100110;
    assign weights1[3][19] = 16'b0000000000010100;
    assign weights1[3][20] = 16'b0000000000010011;
    assign weights1[3][21] = 16'b0000000000000110;
    assign weights1[3][22] = 16'b0000000000000011;
    assign weights1[3][23] = 16'b1111111111111101;
    assign weights1[3][24] = 16'b1111111111111010;
    assign weights1[3][25] = 16'b1111111111111100;
    assign weights1[3][26] = 16'b1111111111111111;
    assign weights1[3][27] = 16'b0000000000000000;
    assign weights1[3][28] = 16'b1111111111111111;
    assign weights1[3][29] = 16'b0000000000000000;
    assign weights1[3][30] = 16'b0000000000000000;
    assign weights1[3][31] = 16'b1111111111111111;
    assign weights1[3][32] = 16'b1111111111111011;
    assign weights1[3][33] = 16'b1111111111111011;
    assign weights1[3][34] = 16'b1111111111111111;
    assign weights1[3][35] = 16'b0000000000000011;
    assign weights1[3][36] = 16'b0000000000000110;
    assign weights1[3][37] = 16'b1111111111101110;
    assign weights1[3][38] = 16'b1111111111101110;
    assign weights1[3][39] = 16'b1111111111100000;
    assign weights1[3][40] = 16'b1111111111000111;
    assign weights1[3][41] = 16'b1111111111000000;
    assign weights1[3][42] = 16'b1111111111000011;
    assign weights1[3][43] = 16'b1111111111100001;
    assign weights1[3][44] = 16'b1111111111111011;
    assign weights1[3][45] = 16'b0000000000101111;
    assign weights1[3][46] = 16'b0000000000100101;
    assign weights1[3][47] = 16'b0000000000100001;
    assign weights1[3][48] = 16'b0000000000010011;
    assign weights1[3][49] = 16'b0000000000001100;
    assign weights1[3][50] = 16'b0000000000001101;
    assign weights1[3][51] = 16'b0000000000000010;
    assign weights1[3][52] = 16'b1111111111101101;
    assign weights1[3][53] = 16'b1111111111110111;
    assign weights1[3][54] = 16'b1111111111111011;
    assign weights1[3][55] = 16'b1111111111111110;
    assign weights1[3][56] = 16'b0000000000000000;
    assign weights1[3][57] = 16'b0000000000000000;
    assign weights1[3][58] = 16'b0000000000000001;
    assign weights1[3][59] = 16'b1111111111111011;
    assign weights1[3][60] = 16'b1111111111110110;
    assign weights1[3][61] = 16'b1111111111111010;
    assign weights1[3][62] = 16'b1111111111111011;
    assign weights1[3][63] = 16'b1111111111111001;
    assign weights1[3][64] = 16'b0000000000010011;
    assign weights1[3][65] = 16'b0000000000001001;
    assign weights1[3][66] = 16'b1111111111011110;
    assign weights1[3][67] = 16'b1111111111100101;
    assign weights1[3][68] = 16'b1111111110111111;
    assign weights1[3][69] = 16'b1111111110011001;
    assign weights1[3][70] = 16'b1111111110011000;
    assign weights1[3][71] = 16'b1111111111001111;
    assign weights1[3][72] = 16'b0000000000011110;
    assign weights1[3][73] = 16'b0000000000011101;
    assign weights1[3][74] = 16'b0000000000010010;
    assign weights1[3][75] = 16'b0000000000001010;
    assign weights1[3][76] = 16'b0000000000010011;
    assign weights1[3][77] = 16'b1111111111110111;
    assign weights1[3][78] = 16'b1111111111110100;
    assign weights1[3][79] = 16'b1111111111101000;
    assign weights1[3][80] = 16'b1111111111101011;
    assign weights1[3][81] = 16'b1111111111110011;
    assign weights1[3][82] = 16'b1111111111110001;
    assign weights1[3][83] = 16'b1111111111111000;
    assign weights1[3][84] = 16'b0000000000000001;
    assign weights1[3][85] = 16'b0000000000000001;
    assign weights1[3][86] = 16'b0000000000000011;
    assign weights1[3][87] = 16'b0000000000000000;
    assign weights1[3][88] = 16'b1111111111111000;
    assign weights1[3][89] = 16'b1111111111111111;
    assign weights1[3][90] = 16'b1111111111111010;
    assign weights1[3][91] = 16'b1111111111111100;
    assign weights1[3][92] = 16'b0000000000000110;
    assign weights1[3][93] = 16'b0000000000000011;
    assign weights1[3][94] = 16'b1111111111110111;
    assign weights1[3][95] = 16'b1111111111100100;
    assign weights1[3][96] = 16'b1111111111001000;
    assign weights1[3][97] = 16'b1111111101111111;
    assign weights1[3][98] = 16'b1111111110000101;
    assign weights1[3][99] = 16'b1111111111000011;
    assign weights1[3][100] = 16'b1111111111010111;
    assign weights1[3][101] = 16'b0000000000011001;
    assign weights1[3][102] = 16'b0000000000001100;
    assign weights1[3][103] = 16'b0000000000010100;
    assign weights1[3][104] = 16'b1111111111011110;
    assign weights1[3][105] = 16'b1111111111101000;
    assign weights1[3][106] = 16'b0000000000001010;
    assign weights1[3][107] = 16'b1111111111101001;
    assign weights1[3][108] = 16'b1111111111100110;
    assign weights1[3][109] = 16'b1111111111100100;
    assign weights1[3][110] = 16'b1111111111100110;
    assign weights1[3][111] = 16'b1111111111110111;
    assign weights1[3][112] = 16'b0000000000000100;
    assign weights1[3][113] = 16'b0000000000000100;
    assign weights1[3][114] = 16'b0000000000000000;
    assign weights1[3][115] = 16'b0000000000000001;
    assign weights1[3][116] = 16'b1111111111111001;
    assign weights1[3][117] = 16'b1111111111111011;
    assign weights1[3][118] = 16'b1111111111110110;
    assign weights1[3][119] = 16'b0000000000000001;
    assign weights1[3][120] = 16'b1111111111111111;
    assign weights1[3][121] = 16'b0000000000010000;
    assign weights1[3][122] = 16'b1111111111110111;
    assign weights1[3][123] = 16'b1111111111110100;
    assign weights1[3][124] = 16'b1111111111001111;
    assign weights1[3][125] = 16'b1111111101111001;
    assign weights1[3][126] = 16'b1111111101100101;
    assign weights1[3][127] = 16'b1111111110110000;
    assign weights1[3][128] = 16'b0000000000010001;
    assign weights1[3][129] = 16'b0000000000000111;
    assign weights1[3][130] = 16'b0000000000001010;
    assign weights1[3][131] = 16'b1111111111111001;
    assign weights1[3][132] = 16'b0000000000001110;
    assign weights1[3][133] = 16'b1111111111111110;
    assign weights1[3][134] = 16'b1111111111101010;
    assign weights1[3][135] = 16'b1111111111110111;
    assign weights1[3][136] = 16'b1111111111001110;
    assign weights1[3][137] = 16'b1111111111011111;
    assign weights1[3][138] = 16'b1111111111100101;
    assign weights1[3][139] = 16'b1111111111110010;
    assign weights1[3][140] = 16'b0000000000001000;
    assign weights1[3][141] = 16'b0000000000000001;
    assign weights1[3][142] = 16'b0000000000000000;
    assign weights1[3][143] = 16'b0000000000001010;
    assign weights1[3][144] = 16'b1111111111110011;
    assign weights1[3][145] = 16'b1111111111111101;
    assign weights1[3][146] = 16'b0000000000000100;
    assign weights1[3][147] = 16'b0000000000000001;
    assign weights1[3][148] = 16'b0000000000000001;
    assign weights1[3][149] = 16'b0000000000000001;
    assign weights1[3][150] = 16'b0000000000010001;
    assign weights1[3][151] = 16'b1111111111111101;
    assign weights1[3][152] = 16'b1111111111000001;
    assign weights1[3][153] = 16'b1111111101100000;
    assign weights1[3][154] = 16'b1111111101000110;
    assign weights1[3][155] = 16'b1111111110100000;
    assign weights1[3][156] = 16'b0000000000110001;
    assign weights1[3][157] = 16'b0000000000111100;
    assign weights1[3][158] = 16'b0000000000100111;
    assign weights1[3][159] = 16'b1111111111111110;
    assign weights1[3][160] = 16'b0000000000001001;
    assign weights1[3][161] = 16'b0000000000010010;
    assign weights1[3][162] = 16'b0000000000000001;
    assign weights1[3][163] = 16'b1111111111001000;
    assign weights1[3][164] = 16'b1111111111001010;
    assign weights1[3][165] = 16'b1111111111010110;
    assign weights1[3][166] = 16'b1111111111101010;
    assign weights1[3][167] = 16'b1111111111110100;
    assign weights1[3][168] = 16'b0000000000000100;
    assign weights1[3][169] = 16'b1111111111111101;
    assign weights1[3][170] = 16'b1111111111111111;
    assign weights1[3][171] = 16'b1111111111111011;
    assign weights1[3][172] = 16'b0000000000000000;
    assign weights1[3][173] = 16'b0000000000000010;
    assign weights1[3][174] = 16'b1111111111111111;
    assign weights1[3][175] = 16'b1111111111111000;
    assign weights1[3][176] = 16'b0000000000000011;
    assign weights1[3][177] = 16'b0000000000011011;
    assign weights1[3][178] = 16'b0000000000010100;
    assign weights1[3][179] = 16'b0000000000000110;
    assign weights1[3][180] = 16'b1111111111010100;
    assign weights1[3][181] = 16'b1111111101110001;
    assign weights1[3][182] = 16'b1111111100000100;
    assign weights1[3][183] = 16'b1111111111000111;
    assign weights1[3][184] = 16'b0000000000010111;
    assign weights1[3][185] = 16'b0000000000110011;
    assign weights1[3][186] = 16'b0000000000010011;
    assign weights1[3][187] = 16'b0000000000001010;
    assign weights1[3][188] = 16'b0000000000101111;
    assign weights1[3][189] = 16'b1111111111111111;
    assign weights1[3][190] = 16'b1111111111100101;
    assign weights1[3][191] = 16'b1111111111001000;
    assign weights1[3][192] = 16'b1111111111001011;
    assign weights1[3][193] = 16'b1111111111010000;
    assign weights1[3][194] = 16'b1111111111011110;
    assign weights1[3][195] = 16'b1111111111101101;
    assign weights1[3][196] = 16'b1111111111111110;
    assign weights1[3][197] = 16'b1111111111111011;
    assign weights1[3][198] = 16'b1111111111111100;
    assign weights1[3][199] = 16'b0000000000000111;
    assign weights1[3][200] = 16'b1111111111101001;
    assign weights1[3][201] = 16'b0000000000011000;
    assign weights1[3][202] = 16'b0000000000000110;
    assign weights1[3][203] = 16'b0000000000010101;
    assign weights1[3][204] = 16'b0000000000010100;
    assign weights1[3][205] = 16'b0000000000010010;
    assign weights1[3][206] = 16'b0000000000100011;
    assign weights1[3][207] = 16'b0000000000100000;
    assign weights1[3][208] = 16'b1111111111100101;
    assign weights1[3][209] = 16'b1111111101000010;
    assign weights1[3][210] = 16'b1111111011110010;
    assign weights1[3][211] = 16'b1111111111111111;
    assign weights1[3][212] = 16'b0000000000111100;
    assign weights1[3][213] = 16'b0000000000101100;
    assign weights1[3][214] = 16'b0000000000001001;
    assign weights1[3][215] = 16'b0000000000010111;
    assign weights1[3][216] = 16'b0000000000000011;
    assign weights1[3][217] = 16'b0000000000000111;
    assign weights1[3][218] = 16'b1111111111010100;
    assign weights1[3][219] = 16'b1111111110111001;
    assign weights1[3][220] = 16'b1111111110111111;
    assign weights1[3][221] = 16'b1111111111010011;
    assign weights1[3][222] = 16'b1111111111100001;
    assign weights1[3][223] = 16'b1111111111110101;
    assign weights1[3][224] = 16'b1111111111111111;
    assign weights1[3][225] = 16'b1111111111111100;
    assign weights1[3][226] = 16'b1111111111111101;
    assign weights1[3][227] = 16'b1111111111111110;
    assign weights1[3][228] = 16'b1111111111111101;
    assign weights1[3][229] = 16'b0000000000000110;
    assign weights1[3][230] = 16'b0000000000100010;
    assign weights1[3][231] = 16'b0000000000000111;
    assign weights1[3][232] = 16'b1111111111110011;
    assign weights1[3][233] = 16'b0000000000101001;
    assign weights1[3][234] = 16'b0000000000000010;
    assign weights1[3][235] = 16'b0000000000101101;
    assign weights1[3][236] = 16'b1111111111100100;
    assign weights1[3][237] = 16'b1111111101000010;
    assign weights1[3][238] = 16'b1111111101010010;
    assign weights1[3][239] = 16'b0000000000100011;
    assign weights1[3][240] = 16'b0000000000100010;
    assign weights1[3][241] = 16'b0000000000101001;
    assign weights1[3][242] = 16'b0000000000100101;
    assign weights1[3][243] = 16'b0000000000000010;
    assign weights1[3][244] = 16'b0000000000010111;
    assign weights1[3][245] = 16'b0000000000000010;
    assign weights1[3][246] = 16'b1111111110111101;
    assign weights1[3][247] = 16'b1111111110101111;
    assign weights1[3][248] = 16'b1111111110101111;
    assign weights1[3][249] = 16'b1111111111010100;
    assign weights1[3][250] = 16'b1111111111100111;
    assign weights1[3][251] = 16'b0000000000000000;
    assign weights1[3][252] = 16'b1111111111111101;
    assign weights1[3][253] = 16'b1111111111111100;
    assign weights1[3][254] = 16'b1111111111111100;
    assign weights1[3][255] = 16'b1111111111111111;
    assign weights1[3][256] = 16'b1111111111110110;
    assign weights1[3][257] = 16'b1111111111111110;
    assign weights1[3][258] = 16'b1111111111111010;
    assign weights1[3][259] = 16'b1111111111110110;
    assign weights1[3][260] = 16'b0000000000011010;
    assign weights1[3][261] = 16'b0000000000001111;
    assign weights1[3][262] = 16'b0000000000101101;
    assign weights1[3][263] = 16'b0000000000101010;
    assign weights1[3][264] = 16'b1111111111011001;
    assign weights1[3][265] = 16'b1111111101000101;
    assign weights1[3][266] = 16'b1111111110001101;
    assign weights1[3][267] = 16'b0000000000001110;
    assign weights1[3][268] = 16'b0000000000100011;
    assign weights1[3][269] = 16'b0000000000010100;
    assign weights1[3][270] = 16'b0000000000011100;
    assign weights1[3][271] = 16'b0000000000010101;
    assign weights1[3][272] = 16'b0000000000010001;
    assign weights1[3][273] = 16'b1111111111111000;
    assign weights1[3][274] = 16'b1111111110011101;
    assign weights1[3][275] = 16'b1111111111001101;
    assign weights1[3][276] = 16'b1111111111010011;
    assign weights1[3][277] = 16'b1111111111101111;
    assign weights1[3][278] = 16'b1111111111111111;
    assign weights1[3][279] = 16'b0000000000011000;
    assign weights1[3][280] = 16'b1111111111111110;
    assign weights1[3][281] = 16'b0000000000000101;
    assign weights1[3][282] = 16'b1111111111111000;
    assign weights1[3][283] = 16'b0000000000000000;
    assign weights1[3][284] = 16'b1111111111111000;
    assign weights1[3][285] = 16'b1111111111110100;
    assign weights1[3][286] = 16'b1111111111101110;
    assign weights1[3][287] = 16'b0000000000011011;
    assign weights1[3][288] = 16'b1111111111111101;
    assign weights1[3][289] = 16'b0000000000000000;
    assign weights1[3][290] = 16'b0000000000101010;
    assign weights1[3][291] = 16'b0000000000110110;
    assign weights1[3][292] = 16'b1111111111010100;
    assign weights1[3][293] = 16'b1111111101111000;
    assign weights1[3][294] = 16'b1111111111010100;
    assign weights1[3][295] = 16'b0000000000001101;
    assign weights1[3][296] = 16'b0000000000010111;
    assign weights1[3][297] = 16'b0000000000100001;
    assign weights1[3][298] = 16'b0000000000001110;
    assign weights1[3][299] = 16'b0000000000010001;
    assign weights1[3][300] = 16'b1111111111100110;
    assign weights1[3][301] = 16'b1111111110111111;
    assign weights1[3][302] = 16'b1111111110111011;
    assign weights1[3][303] = 16'b1111111111000011;
    assign weights1[3][304] = 16'b1111111111101000;
    assign weights1[3][305] = 16'b0000000000010110;
    assign weights1[3][306] = 16'b0000000000100111;
    assign weights1[3][307] = 16'b0000000000100111;
    assign weights1[3][308] = 16'b0000000000000100;
    assign weights1[3][309] = 16'b0000000000000110;
    assign weights1[3][310] = 16'b1111111111101111;
    assign weights1[3][311] = 16'b1111111111111110;
    assign weights1[3][312] = 16'b1111111111111101;
    assign weights1[3][313] = 16'b0000000000000000;
    assign weights1[3][314] = 16'b1111111111111000;
    assign weights1[3][315] = 16'b0000000000000010;
    assign weights1[3][316] = 16'b0000000000001000;
    assign weights1[3][317] = 16'b0000000000100001;
    assign weights1[3][318] = 16'b0000000000100101;
    assign weights1[3][319] = 16'b0000000000011101;
    assign weights1[3][320] = 16'b1111111111010000;
    assign weights1[3][321] = 16'b1111111110101110;
    assign weights1[3][322] = 16'b1111111111011011;
    assign weights1[3][323] = 16'b0000000000001011;
    assign weights1[3][324] = 16'b0000000000011100;
    assign weights1[3][325] = 16'b0000000000011110;
    assign weights1[3][326] = 16'b0000000000100000;
    assign weights1[3][327] = 16'b1111111111101011;
    assign weights1[3][328] = 16'b0000000000000001;
    assign weights1[3][329] = 16'b1111111111000011;
    assign weights1[3][330] = 16'b1111111111000010;
    assign weights1[3][331] = 16'b1111111111001011;
    assign weights1[3][332] = 16'b0000000000000001;
    assign weights1[3][333] = 16'b0000000000110000;
    assign weights1[3][334] = 16'b0000000000101010;
    assign weights1[3][335] = 16'b0000000000011111;
    assign weights1[3][336] = 16'b1111111111111101;
    assign weights1[3][337] = 16'b0000000000001010;
    assign weights1[3][338] = 16'b0000000000001010;
    assign weights1[3][339] = 16'b0000000000010111;
    assign weights1[3][340] = 16'b0000000000000100;
    assign weights1[3][341] = 16'b0000000000000111;
    assign weights1[3][342] = 16'b0000000000000010;
    assign weights1[3][343] = 16'b0000000000101011;
    assign weights1[3][344] = 16'b1111111111110100;
    assign weights1[3][345] = 16'b0000000000001101;
    assign weights1[3][346] = 16'b0000000000100011;
    assign weights1[3][347] = 16'b0000000000011110;
    assign weights1[3][348] = 16'b1111111111011111;
    assign weights1[3][349] = 16'b1111111111001011;
    assign weights1[3][350] = 16'b1111111111011001;
    assign weights1[3][351] = 16'b0000000000000010;
    assign weights1[3][352] = 16'b0000000000001110;
    assign weights1[3][353] = 16'b0000000000100011;
    assign weights1[3][354] = 16'b1111111111111000;
    assign weights1[3][355] = 16'b1111111111111111;
    assign weights1[3][356] = 16'b1111111111111010;
    assign weights1[3][357] = 16'b1111111111000101;
    assign weights1[3][358] = 16'b1111111111100011;
    assign weights1[3][359] = 16'b1111111111111011;
    assign weights1[3][360] = 16'b0000000000110111;
    assign weights1[3][361] = 16'b0000000000011111;
    assign weights1[3][362] = 16'b0000000000011101;
    assign weights1[3][363] = 16'b0000000000001001;
    assign weights1[3][364] = 16'b1111111111111111;
    assign weights1[3][365] = 16'b0000000000001111;
    assign weights1[3][366] = 16'b0000000000001011;
    assign weights1[3][367] = 16'b1111111111111100;
    assign weights1[3][368] = 16'b0000000000001010;
    assign weights1[3][369] = 16'b0000000000001010;
    assign weights1[3][370] = 16'b0000000000010000;
    assign weights1[3][371] = 16'b1111111111100111;
    assign weights1[3][372] = 16'b0000000000001100;
    assign weights1[3][373] = 16'b0000000000000100;
    assign weights1[3][374] = 16'b0000000000010100;
    assign weights1[3][375] = 16'b0000000000100010;
    assign weights1[3][376] = 16'b1111111111111100;
    assign weights1[3][377] = 16'b1111111111101000;
    assign weights1[3][378] = 16'b1111111111111000;
    assign weights1[3][379] = 16'b1111111111111010;
    assign weights1[3][380] = 16'b1111111111111011;
    assign weights1[3][381] = 16'b0000000000000000;
    assign weights1[3][382] = 16'b1111111111111010;
    assign weights1[3][383] = 16'b1111111111111110;
    assign weights1[3][384] = 16'b1111111111011110;
    assign weights1[3][385] = 16'b1111111111011010;
    assign weights1[3][386] = 16'b1111111111011011;
    assign weights1[3][387] = 16'b0000000000001101;
    assign weights1[3][388] = 16'b0000000000011011;
    assign weights1[3][389] = 16'b0000000000001011;
    assign weights1[3][390] = 16'b1111111111111101;
    assign weights1[3][391] = 16'b1111111111111111;
    assign weights1[3][392] = 16'b0000000000000000;
    assign weights1[3][393] = 16'b0000000000001010;
    assign weights1[3][394] = 16'b0000000000001101;
    assign weights1[3][395] = 16'b1111111111110100;
    assign weights1[3][396] = 16'b1111111111110100;
    assign weights1[3][397] = 16'b1111111111111010;
    assign weights1[3][398] = 16'b1111111111101000;
    assign weights1[3][399] = 16'b0000000000000011;
    assign weights1[3][400] = 16'b0000000000010000;
    assign weights1[3][401] = 16'b0000000000000101;
    assign weights1[3][402] = 16'b0000000000001011;
    assign weights1[3][403] = 16'b0000000000011011;
    assign weights1[3][404] = 16'b0000000000001100;
    assign weights1[3][405] = 16'b1111111111101001;
    assign weights1[3][406] = 16'b1111111111101010;
    assign weights1[3][407] = 16'b0000000000000100;
    assign weights1[3][408] = 16'b0000000000001100;
    assign weights1[3][409] = 16'b0000000000001001;
    assign weights1[3][410] = 16'b0000000000000011;
    assign weights1[3][411] = 16'b1111111111111010;
    assign weights1[3][412] = 16'b1111111111100001;
    assign weights1[3][413] = 16'b1111111111110001;
    assign weights1[3][414] = 16'b0000000000000001;
    assign weights1[3][415] = 16'b0000000000010000;
    assign weights1[3][416] = 16'b0000000000010001;
    assign weights1[3][417] = 16'b0000000000010001;
    assign weights1[3][418] = 16'b0000000000000101;
    assign weights1[3][419] = 16'b1111111111110110;
    assign weights1[3][420] = 16'b0000000000001011;
    assign weights1[3][421] = 16'b0000000000001001;
    assign weights1[3][422] = 16'b0000000000001100;
    assign weights1[3][423] = 16'b1111111111111001;
    assign weights1[3][424] = 16'b0000000000001001;
    assign weights1[3][425] = 16'b0000000000000010;
    assign weights1[3][426] = 16'b0000000000010101;
    assign weights1[3][427] = 16'b0000000000000001;
    assign weights1[3][428] = 16'b0000000000001101;
    assign weights1[3][429] = 16'b0000000000001011;
    assign weights1[3][430] = 16'b0000000000000110;
    assign weights1[3][431] = 16'b0000000000001001;
    assign weights1[3][432] = 16'b0000000000000101;
    assign weights1[3][433] = 16'b0000000000001101;
    assign weights1[3][434] = 16'b1111111111110010;
    assign weights1[3][435] = 16'b1111111111111000;
    assign weights1[3][436] = 16'b0000000000000100;
    assign weights1[3][437] = 16'b0000000000000010;
    assign weights1[3][438] = 16'b1111111111110010;
    assign weights1[3][439] = 16'b0000000000000001;
    assign weights1[3][440] = 16'b1111111111101011;
    assign weights1[3][441] = 16'b1111111111110000;
    assign weights1[3][442] = 16'b0000000000010111;
    assign weights1[3][443] = 16'b0000000000011111;
    assign weights1[3][444] = 16'b1111111111111111;
    assign weights1[3][445] = 16'b1111111111110000;
    assign weights1[3][446] = 16'b1111111111111011;
    assign weights1[3][447] = 16'b1111111111111101;
    assign weights1[3][448] = 16'b0000000000000110;
    assign weights1[3][449] = 16'b0000000000000010;
    assign weights1[3][450] = 16'b0000000000000010;
    assign weights1[3][451] = 16'b1111111111111101;
    assign weights1[3][452] = 16'b1111111111111110;
    assign weights1[3][453] = 16'b1111111111111100;
    assign weights1[3][454] = 16'b0000000000000110;
    assign weights1[3][455] = 16'b0000000000000100;
    assign weights1[3][456] = 16'b1111111111110100;
    assign weights1[3][457] = 16'b1111111111111111;
    assign weights1[3][458] = 16'b0000000000001010;
    assign weights1[3][459] = 16'b0000000000000101;
    assign weights1[3][460] = 16'b0000000000000110;
    assign weights1[3][461] = 16'b0000000000000011;
    assign weights1[3][462] = 16'b0000000000001101;
    assign weights1[3][463] = 16'b0000000000000001;
    assign weights1[3][464] = 16'b1111111111101111;
    assign weights1[3][465] = 16'b1111111111111010;
    assign weights1[3][466] = 16'b1111111111110011;
    assign weights1[3][467] = 16'b1111111111111100;
    assign weights1[3][468] = 16'b0000000000000000;
    assign weights1[3][469] = 16'b1111111111111111;
    assign weights1[3][470] = 16'b1111111111111010;
    assign weights1[3][471] = 16'b0000000000000111;
    assign weights1[3][472] = 16'b0000000000000001;
    assign weights1[3][473] = 16'b1111111111101101;
    assign weights1[3][474] = 16'b1111111111111001;
    assign weights1[3][475] = 16'b1111111111111101;
    assign weights1[3][476] = 16'b0000000000000101;
    assign weights1[3][477] = 16'b0000000000000101;
    assign weights1[3][478] = 16'b0000000000001001;
    assign weights1[3][479] = 16'b1111111111110110;
    assign weights1[3][480] = 16'b0000000000000111;
    assign weights1[3][481] = 16'b0000000000100101;
    assign weights1[3][482] = 16'b1111111111101111;
    assign weights1[3][483] = 16'b0000000000010000;
    assign weights1[3][484] = 16'b1111111111101011;
    assign weights1[3][485] = 16'b1111111111111010;
    assign weights1[3][486] = 16'b0000000000000001;
    assign weights1[3][487] = 16'b0000000000000101;
    assign weights1[3][488] = 16'b0000000000000011;
    assign weights1[3][489] = 16'b1111111111110111;
    assign weights1[3][490] = 16'b0000000000000000;
    assign weights1[3][491] = 16'b1111111111110111;
    assign weights1[3][492] = 16'b1111111111111011;
    assign weights1[3][493] = 16'b1111111111110010;
    assign weights1[3][494] = 16'b1111111111111001;
    assign weights1[3][495] = 16'b1111111111111010;
    assign weights1[3][496] = 16'b0000000000001110;
    assign weights1[3][497] = 16'b0000000000001011;
    assign weights1[3][498] = 16'b0000000000000010;
    assign weights1[3][499] = 16'b1111111111110110;
    assign weights1[3][500] = 16'b1111111111110000;
    assign weights1[3][501] = 16'b1111111111110001;
    assign weights1[3][502] = 16'b1111111111101111;
    assign weights1[3][503] = 16'b1111111111111001;
    assign weights1[3][504] = 16'b0000000000000011;
    assign weights1[3][505] = 16'b1111111111111110;
    assign weights1[3][506] = 16'b1111111111111010;
    assign weights1[3][507] = 16'b1111111111110101;
    assign weights1[3][508] = 16'b0000000000011011;
    assign weights1[3][509] = 16'b0000000000000001;
    assign weights1[3][510] = 16'b0000000000000101;
    assign weights1[3][511] = 16'b1111111111111100;
    assign weights1[3][512] = 16'b0000000000001010;
    assign weights1[3][513] = 16'b0000000000000111;
    assign weights1[3][514] = 16'b0000000000010101;
    assign weights1[3][515] = 16'b0000000000010010;
    assign weights1[3][516] = 16'b0000000000000011;
    assign weights1[3][517] = 16'b1111111111111011;
    assign weights1[3][518] = 16'b1111111111110010;
    assign weights1[3][519] = 16'b1111111111101010;
    assign weights1[3][520] = 16'b1111111111110001;
    assign weights1[3][521] = 16'b1111111111111011;
    assign weights1[3][522] = 16'b1111111111111101;
    assign weights1[3][523] = 16'b1111111111111001;
    assign weights1[3][524] = 16'b1111111111110100;
    assign weights1[3][525] = 16'b1111111111101010;
    assign weights1[3][526] = 16'b1111111111110010;
    assign weights1[3][527] = 16'b1111111111100111;
    assign weights1[3][528] = 16'b1111111111110101;
    assign weights1[3][529] = 16'b1111111111111100;
    assign weights1[3][530] = 16'b1111111111111011;
    assign weights1[3][531] = 16'b1111111111111000;
    assign weights1[3][532] = 16'b0000000000000000;
    assign weights1[3][533] = 16'b1111111111111011;
    assign weights1[3][534] = 16'b0000000000000000;
    assign weights1[3][535] = 16'b0000000000000101;
    assign weights1[3][536] = 16'b0000000000000010;
    assign weights1[3][537] = 16'b1111111111111011;
    assign weights1[3][538] = 16'b1111111111110110;
    assign weights1[3][539] = 16'b1111111111111110;
    assign weights1[3][540] = 16'b1111111111111111;
    assign weights1[3][541] = 16'b1111111111110101;
    assign weights1[3][542] = 16'b1111111111110110;
    assign weights1[3][543] = 16'b0000000000001000;
    assign weights1[3][544] = 16'b0000000000000001;
    assign weights1[3][545] = 16'b1111111111111000;
    assign weights1[3][546] = 16'b0000000000000110;
    assign weights1[3][547] = 16'b1111111111101101;
    assign weights1[3][548] = 16'b1111111111111111;
    assign weights1[3][549] = 16'b1111111111111000;
    assign weights1[3][550] = 16'b0000000000000010;
    assign weights1[3][551] = 16'b1111111111111110;
    assign weights1[3][552] = 16'b1111111111101111;
    assign weights1[3][553] = 16'b1111111111111100;
    assign weights1[3][554] = 16'b1111111111110110;
    assign weights1[3][555] = 16'b1111111111101101;
    assign weights1[3][556] = 16'b0000000000000110;
    assign weights1[3][557] = 16'b1111111111111111;
    assign weights1[3][558] = 16'b0000000000001000;
    assign weights1[3][559] = 16'b0000000000000101;
    assign weights1[3][560] = 16'b0000000000000101;
    assign weights1[3][561] = 16'b1111111111110111;
    assign weights1[3][562] = 16'b1111111111111100;
    assign weights1[3][563] = 16'b1111111111111111;
    assign weights1[3][564] = 16'b0000000000000000;
    assign weights1[3][565] = 16'b1111111111110011;
    assign weights1[3][566] = 16'b0000000000001001;
    assign weights1[3][567] = 16'b1111111111101100;
    assign weights1[3][568] = 16'b1111111111110010;
    assign weights1[3][569] = 16'b0000000000000101;
    assign weights1[3][570] = 16'b0000000000000010;
    assign weights1[3][571] = 16'b0000000000000101;
    assign weights1[3][572] = 16'b0000000000000111;
    assign weights1[3][573] = 16'b1111111111111011;
    assign weights1[3][574] = 16'b1111111111100011;
    assign weights1[3][575] = 16'b0000000000000010;
    assign weights1[3][576] = 16'b1111111111110101;
    assign weights1[3][577] = 16'b1111111111110110;
    assign weights1[3][578] = 16'b1111111111101111;
    assign weights1[3][579] = 16'b0000000000000011;
    assign weights1[3][580] = 16'b1111111111111000;
    assign weights1[3][581] = 16'b1111111111110001;
    assign weights1[3][582] = 16'b1111111111110100;
    assign weights1[3][583] = 16'b0000000000000111;
    assign weights1[3][584] = 16'b0000000000010001;
    assign weights1[3][585] = 16'b0000000000001111;
    assign weights1[3][586] = 16'b0000000000001001;
    assign weights1[3][587] = 16'b0000000000001100;
    assign weights1[3][588] = 16'b1111111111111101;
    assign weights1[3][589] = 16'b1111111111111111;
    assign weights1[3][590] = 16'b0000000000000110;
    assign weights1[3][591] = 16'b1111111111111011;
    assign weights1[3][592] = 16'b1111111111110000;
    assign weights1[3][593] = 16'b1111111111110100;
    assign weights1[3][594] = 16'b1111111111111110;
    assign weights1[3][595] = 16'b0000000000000100;
    assign weights1[3][596] = 16'b0000000000101111;
    assign weights1[3][597] = 16'b1111111111110111;
    assign weights1[3][598] = 16'b1111111111111000;
    assign weights1[3][599] = 16'b0000000000000100;
    assign weights1[3][600] = 16'b1111111111110101;
    assign weights1[3][601] = 16'b1111111111111111;
    assign weights1[3][602] = 16'b1111111111111011;
    assign weights1[3][603] = 16'b1111111111110111;
    assign weights1[3][604] = 16'b1111111111111000;
    assign weights1[3][605] = 16'b0000000000000001;
    assign weights1[3][606] = 16'b0000000000001011;
    assign weights1[3][607] = 16'b0000000000000100;
    assign weights1[3][608] = 16'b1111111111111011;
    assign weights1[3][609] = 16'b1111111111011101;
    assign weights1[3][610] = 16'b1111111111111010;
    assign weights1[3][611] = 16'b1111111111111110;
    assign weights1[3][612] = 16'b0000000000001100;
    assign weights1[3][613] = 16'b1111111111111011;
    assign weights1[3][614] = 16'b0000000000001000;
    assign weights1[3][615] = 16'b0000000000001001;
    assign weights1[3][616] = 16'b1111111111111011;
    assign weights1[3][617] = 16'b1111111111111001;
    assign weights1[3][618] = 16'b0000000000000110;
    assign weights1[3][619] = 16'b1111111111110101;
    assign weights1[3][620] = 16'b1111111111111011;
    assign weights1[3][621] = 16'b0000000000001011;
    assign weights1[3][622] = 16'b0000000000001000;
    assign weights1[3][623] = 16'b0000000000000011;
    assign weights1[3][624] = 16'b1111111111111010;
    assign weights1[3][625] = 16'b1111111111110111;
    assign weights1[3][626] = 16'b0000000000000001;
    assign weights1[3][627] = 16'b1111111111101100;
    assign weights1[3][628] = 16'b1111111111111111;
    assign weights1[3][629] = 16'b0000000000000111;
    assign weights1[3][630] = 16'b1111111111111110;
    assign weights1[3][631] = 16'b0000000000000000;
    assign weights1[3][632] = 16'b1111111111110110;
    assign weights1[3][633] = 16'b1111111111110000;
    assign weights1[3][634] = 16'b1111111111011101;
    assign weights1[3][635] = 16'b1111111111111101;
    assign weights1[3][636] = 16'b0000000000010000;
    assign weights1[3][637] = 16'b0000000000000001;
    assign weights1[3][638] = 16'b1111111111101110;
    assign weights1[3][639] = 16'b1111111111111010;
    assign weights1[3][640] = 16'b1111111111111101;
    assign weights1[3][641] = 16'b1111111111110100;
    assign weights1[3][642] = 16'b0000000000000011;
    assign weights1[3][643] = 16'b0000000000000010;
    assign weights1[3][644] = 16'b1111111111111001;
    assign weights1[3][645] = 16'b1111111111111011;
    assign weights1[3][646] = 16'b0000000000000010;
    assign weights1[3][647] = 16'b0000000000001000;
    assign weights1[3][648] = 16'b0000000000000000;
    assign weights1[3][649] = 16'b1111111111111010;
    assign weights1[3][650] = 16'b1111111111011011;
    assign weights1[3][651] = 16'b1111111111111110;
    assign weights1[3][652] = 16'b0000000000001110;
    assign weights1[3][653] = 16'b1111111111111000;
    assign weights1[3][654] = 16'b0000000000001100;
    assign weights1[3][655] = 16'b0000000000000110;
    assign weights1[3][656] = 16'b0000000000000000;
    assign weights1[3][657] = 16'b1111111111111110;
    assign weights1[3][658] = 16'b1111111111110001;
    assign weights1[3][659] = 16'b1111111111110111;
    assign weights1[3][660] = 16'b1111111111110011;
    assign weights1[3][661] = 16'b0000000000000111;
    assign weights1[3][662] = 16'b0000000000011001;
    assign weights1[3][663] = 16'b1111111111110101;
    assign weights1[3][664] = 16'b1111111111111011;
    assign weights1[3][665] = 16'b0000000000000111;
    assign weights1[3][666] = 16'b1111111111110100;
    assign weights1[3][667] = 16'b1111111111110010;
    assign weights1[3][668] = 16'b1111111111111000;
    assign weights1[3][669] = 16'b1111111111110111;
    assign weights1[3][670] = 16'b1111111111111110;
    assign weights1[3][671] = 16'b0000000000000010;
    assign weights1[3][672] = 16'b0000000000000001;
    assign weights1[3][673] = 16'b1111111111111011;
    assign weights1[3][674] = 16'b1111111111111110;
    assign weights1[3][675] = 16'b1111111111111101;
    assign weights1[3][676] = 16'b1111111111110111;
    assign weights1[3][677] = 16'b1111111111101100;
    assign weights1[3][678] = 16'b1111111111110010;
    assign weights1[3][679] = 16'b1111111111111000;
    assign weights1[3][680] = 16'b1111111111100110;
    assign weights1[3][681] = 16'b1111111111111010;
    assign weights1[3][682] = 16'b1111111111100101;
    assign weights1[3][683] = 16'b1111111111110111;
    assign weights1[3][684] = 16'b0000000000010110;
    assign weights1[3][685] = 16'b0000000000000011;
    assign weights1[3][686] = 16'b1111111111111000;
    assign weights1[3][687] = 16'b0000000000000101;
    assign weights1[3][688] = 16'b0000000000000101;
    assign weights1[3][689] = 16'b0000000000010110;
    assign weights1[3][690] = 16'b0000000000001101;
    assign weights1[3][691] = 16'b1111111111110100;
    assign weights1[3][692] = 16'b0000000000000110;
    assign weights1[3][693] = 16'b0000000000001010;
    assign weights1[3][694] = 16'b0000000000000100;
    assign weights1[3][695] = 16'b1111111111111001;
    assign weights1[3][696] = 16'b1111111111111101;
    assign weights1[3][697] = 16'b0000000000000001;
    assign weights1[3][698] = 16'b1111111111111101;
    assign weights1[3][699] = 16'b0000000000000001;
    assign weights1[3][700] = 16'b0000000000000000;
    assign weights1[3][701] = 16'b1111111111111100;
    assign weights1[3][702] = 16'b1111111111110110;
    assign weights1[3][703] = 16'b0000000000000010;
    assign weights1[3][704] = 16'b1111111111111001;
    assign weights1[3][705] = 16'b1111111111111110;
    assign weights1[3][706] = 16'b1111111111111101;
    assign weights1[3][707] = 16'b1111111111110011;
    assign weights1[3][708] = 16'b1111111111110011;
    assign weights1[3][709] = 16'b1111111111100001;
    assign weights1[3][710] = 16'b0000000000010001;
    assign weights1[3][711] = 16'b1111111111110101;
    assign weights1[3][712] = 16'b1111111111101011;
    assign weights1[3][713] = 16'b0000000000011011;
    assign weights1[3][714] = 16'b1111111111100111;
    assign weights1[3][715] = 16'b0000000000001001;
    assign weights1[3][716] = 16'b1111111111110111;
    assign weights1[3][717] = 16'b0000000000000100;
    assign weights1[3][718] = 16'b0000000000001001;
    assign weights1[3][719] = 16'b1111111111111100;
    assign weights1[3][720] = 16'b1111111111110001;
    assign weights1[3][721] = 16'b0000000000000111;
    assign weights1[3][722] = 16'b0000000000000101;
    assign weights1[3][723] = 16'b0000000000000111;
    assign weights1[3][724] = 16'b0000000000000011;
    assign weights1[3][725] = 16'b0000000000000011;
    assign weights1[3][726] = 16'b0000000000000001;
    assign weights1[3][727] = 16'b1111111111111111;
    assign weights1[3][728] = 16'b0000000000000000;
    assign weights1[3][729] = 16'b1111111111111110;
    assign weights1[3][730] = 16'b0000000000000000;
    assign weights1[3][731] = 16'b1111111111111111;
    assign weights1[3][732] = 16'b1111111111111111;
    assign weights1[3][733] = 16'b1111111111111001;
    assign weights1[3][734] = 16'b1111111111110111;
    assign weights1[3][735] = 16'b0000000000010000;
    assign weights1[3][736] = 16'b0000000000000000;
    assign weights1[3][737] = 16'b0000000000000011;
    assign weights1[3][738] = 16'b0000000000000010;
    assign weights1[3][739] = 16'b1111111111111011;
    assign weights1[3][740] = 16'b1111111111111110;
    assign weights1[3][741] = 16'b1111111111111000;
    assign weights1[3][742] = 16'b1111111111110100;
    assign weights1[3][743] = 16'b0000000000000000;
    assign weights1[3][744] = 16'b1111111111110111;
    assign weights1[3][745] = 16'b0000000000000100;
    assign weights1[3][746] = 16'b0000000000000000;
    assign weights1[3][747] = 16'b0000000000000101;
    assign weights1[3][748] = 16'b0000000000010100;
    assign weights1[3][749] = 16'b1111111111111011;
    assign weights1[3][750] = 16'b0000000000010000;
    assign weights1[3][751] = 16'b0000000000001011;
    assign weights1[3][752] = 16'b0000000000000100;
    assign weights1[3][753] = 16'b0000000000001000;
    assign weights1[3][754] = 16'b0000000000000010;
    assign weights1[3][755] = 16'b1111111111111111;
    assign weights1[3][756] = 16'b0000000000000000;
    assign weights1[3][757] = 16'b0000000000000010;
    assign weights1[3][758] = 16'b0000000000000101;
    assign weights1[3][759] = 16'b0000000000001000;
    assign weights1[3][760] = 16'b0000000000001000;
    assign weights1[3][761] = 16'b1111111111110010;
    assign weights1[3][762] = 16'b1111111111110001;
    assign weights1[3][763] = 16'b1111111111110100;
    assign weights1[3][764] = 16'b1111111111111100;
    assign weights1[3][765] = 16'b1111111111111011;
    assign weights1[3][766] = 16'b0000000000001000;
    assign weights1[3][767] = 16'b1111111111111000;
    assign weights1[3][768] = 16'b1111111111111110;
    assign weights1[3][769] = 16'b0000000000001010;
    assign weights1[3][770] = 16'b1111111111111100;
    assign weights1[3][771] = 16'b0000000000000111;
    assign weights1[3][772] = 16'b0000000000010000;
    assign weights1[3][773] = 16'b1111111111111011;
    assign weights1[3][774] = 16'b1111111111111101;
    assign weights1[3][775] = 16'b0000000000000111;
    assign weights1[3][776] = 16'b0000000000000100;
    assign weights1[3][777] = 16'b1111111111110101;
    assign weights1[3][778] = 16'b0000000000000111;
    assign weights1[3][779] = 16'b0000000000001000;
    assign weights1[3][780] = 16'b0000000000000101;
    assign weights1[3][781] = 16'b0000000000000110;
    assign weights1[3][782] = 16'b0000000000000001;
    assign weights1[3][783] = 16'b0000000000000001;
    assign weights1[4][0] = 16'b1111111111111111;
    assign weights1[4][1] = 16'b1111111111111111;
    assign weights1[4][2] = 16'b1111111111111110;
    assign weights1[4][3] = 16'b0000000000000000;
    assign weights1[4][4] = 16'b1111111111111110;
    assign weights1[4][5] = 16'b1111111111111100;
    assign weights1[4][6] = 16'b0000000000000011;
    assign weights1[4][7] = 16'b1111111111111110;
    assign weights1[4][8] = 16'b1111111111111001;
    assign weights1[4][9] = 16'b1111111111110001;
    assign weights1[4][10] = 16'b1111111111110010;
    assign weights1[4][11] = 16'b1111111111110000;
    assign weights1[4][12] = 16'b1111111111101010;
    assign weights1[4][13] = 16'b1111111111110001;
    assign weights1[4][14] = 16'b1111111111101100;
    assign weights1[4][15] = 16'b1111111111101100;
    assign weights1[4][16] = 16'b1111111111101001;
    assign weights1[4][17] = 16'b1111111111101100;
    assign weights1[4][18] = 16'b1111111111110010;
    assign weights1[4][19] = 16'b1111111111110110;
    assign weights1[4][20] = 16'b1111111111110100;
    assign weights1[4][21] = 16'b1111111111110101;
    assign weights1[4][22] = 16'b1111111111110111;
    assign weights1[4][23] = 16'b1111111111111110;
    assign weights1[4][24] = 16'b1111111111111110;
    assign weights1[4][25] = 16'b1111111111111111;
    assign weights1[4][26] = 16'b1111111111111111;
    assign weights1[4][27] = 16'b1111111111111111;
    assign weights1[4][28] = 16'b1111111111111111;
    assign weights1[4][29] = 16'b1111111111111111;
    assign weights1[4][30] = 16'b1111111111111111;
    assign weights1[4][31] = 16'b1111111111111111;
    assign weights1[4][32] = 16'b0000000000000001;
    assign weights1[4][33] = 16'b0000000000000000;
    assign weights1[4][34] = 16'b0000000000001100;
    assign weights1[4][35] = 16'b0000000000000011;
    assign weights1[4][36] = 16'b1111111111110110;
    assign weights1[4][37] = 16'b1111111111110110;
    assign weights1[4][38] = 16'b1111111111110011;
    assign weights1[4][39] = 16'b1111111111110001;
    assign weights1[4][40] = 16'b1111111111110011;
    assign weights1[4][41] = 16'b1111111111100111;
    assign weights1[4][42] = 16'b1111111111110001;
    assign weights1[4][43] = 16'b1111111111101100;
    assign weights1[4][44] = 16'b1111111111110101;
    assign weights1[4][45] = 16'b1111111111100100;
    assign weights1[4][46] = 16'b1111111111111000;
    assign weights1[4][47] = 16'b1111111111101110;
    assign weights1[4][48] = 16'b1111111111101111;
    assign weights1[4][49] = 16'b1111111111101111;
    assign weights1[4][50] = 16'b1111111111110010;
    assign weights1[4][51] = 16'b1111111111110110;
    assign weights1[4][52] = 16'b1111111111111010;
    assign weights1[4][53] = 16'b1111111111111110;
    assign weights1[4][54] = 16'b1111111111111110;
    assign weights1[4][55] = 16'b1111111111111110;
    assign weights1[4][56] = 16'b1111111111111111;
    assign weights1[4][57] = 16'b1111111111111110;
    assign weights1[4][58] = 16'b1111111111111111;
    assign weights1[4][59] = 16'b1111111111111100;
    assign weights1[4][60] = 16'b1111111111111110;
    assign weights1[4][61] = 16'b0000000000000001;
    assign weights1[4][62] = 16'b0000000000000101;
    assign weights1[4][63] = 16'b0000000000001010;
    assign weights1[4][64] = 16'b1111111111111101;
    assign weights1[4][65] = 16'b1111111111110101;
    assign weights1[4][66] = 16'b1111111111111010;
    assign weights1[4][67] = 16'b1111111111111100;
    assign weights1[4][68] = 16'b1111111111111011;
    assign weights1[4][69] = 16'b1111111111111110;
    assign weights1[4][70] = 16'b0000000000000101;
    assign weights1[4][71] = 16'b1111111111110111;
    assign weights1[4][72] = 16'b1111111111110110;
    assign weights1[4][73] = 16'b1111111111101011;
    assign weights1[4][74] = 16'b1111111111110100;
    assign weights1[4][75] = 16'b1111111111110010;
    assign weights1[4][76] = 16'b1111111111101010;
    assign weights1[4][77] = 16'b1111111111100101;
    assign weights1[4][78] = 16'b1111111111101001;
    assign weights1[4][79] = 16'b1111111111101111;
    assign weights1[4][80] = 16'b1111111111110100;
    assign weights1[4][81] = 16'b1111111111111001;
    assign weights1[4][82] = 16'b1111111111111100;
    assign weights1[4][83] = 16'b1111111111111100;
    assign weights1[4][84] = 16'b0000000000000010;
    assign weights1[4][85] = 16'b0000000000000000;
    assign weights1[4][86] = 16'b1111111111111101;
    assign weights1[4][87] = 16'b1111111111111001;
    assign weights1[4][88] = 16'b1111111111111010;
    assign weights1[4][89] = 16'b1111111111111011;
    assign weights1[4][90] = 16'b0000000000000010;
    assign weights1[4][91] = 16'b0000000000000111;
    assign weights1[4][92] = 16'b0000000000000010;
    assign weights1[4][93] = 16'b1111111111111110;
    assign weights1[4][94] = 16'b0000000000001111;
    assign weights1[4][95] = 16'b0000000000000100;
    assign weights1[4][96] = 16'b1111111111100101;
    assign weights1[4][97] = 16'b1111111111110111;
    assign weights1[4][98] = 16'b1111111111011110;
    assign weights1[4][99] = 16'b1111111111110010;
    assign weights1[4][100] = 16'b1111111111011011;
    assign weights1[4][101] = 16'b1111111111010100;
    assign weights1[4][102] = 16'b1111111111011101;
    assign weights1[4][103] = 16'b1111111111100111;
    assign weights1[4][104] = 16'b1111111111001010;
    assign weights1[4][105] = 16'b1111111111011011;
    assign weights1[4][106] = 16'b1111111111011101;
    assign weights1[4][107] = 16'b1111111111100101;
    assign weights1[4][108] = 16'b1111111111110000;
    assign weights1[4][109] = 16'b1111111111110101;
    assign weights1[4][110] = 16'b1111111111110010;
    assign weights1[4][111] = 16'b1111111111110111;
    assign weights1[4][112] = 16'b0000000000000010;
    assign weights1[4][113] = 16'b0000000000000001;
    assign weights1[4][114] = 16'b1111111111111100;
    assign weights1[4][115] = 16'b1111111111111100;
    assign weights1[4][116] = 16'b1111111111110010;
    assign weights1[4][117] = 16'b0000000000000000;
    assign weights1[4][118] = 16'b0000000000000001;
    assign weights1[4][119] = 16'b1111111111111000;
    assign weights1[4][120] = 16'b1111111111111010;
    assign weights1[4][121] = 16'b1111111111110110;
    assign weights1[4][122] = 16'b1111111111011111;
    assign weights1[4][123] = 16'b1111111111010000;
    assign weights1[4][124] = 16'b1111111111110011;
    assign weights1[4][125] = 16'b1111111111010011;
    assign weights1[4][126] = 16'b0000000000000000;
    assign weights1[4][127] = 16'b1111111111100110;
    assign weights1[4][128] = 16'b1111111111100110;
    assign weights1[4][129] = 16'b0000000000001011;
    assign weights1[4][130] = 16'b1111111111101011;
    assign weights1[4][131] = 16'b1111111111100011;
    assign weights1[4][132] = 16'b0000000000000101;
    assign weights1[4][133] = 16'b0000000000001011;
    assign weights1[4][134] = 16'b1111111111100111;
    assign weights1[4][135] = 16'b1111111111011110;
    assign weights1[4][136] = 16'b1111111111100110;
    assign weights1[4][137] = 16'b1111111111111101;
    assign weights1[4][138] = 16'b1111111111111001;
    assign weights1[4][139] = 16'b1111111111111001;
    assign weights1[4][140] = 16'b0000000000000011;
    assign weights1[4][141] = 16'b1111111111111101;
    assign weights1[4][142] = 16'b1111111111111000;
    assign weights1[4][143] = 16'b0000000000000101;
    assign weights1[4][144] = 16'b0000000000001001;
    assign weights1[4][145] = 16'b1111111111011110;
    assign weights1[4][146] = 16'b1111111111100110;
    assign weights1[4][147] = 16'b1111111111110101;
    assign weights1[4][148] = 16'b1111111111111011;
    assign weights1[4][149] = 16'b0000000000001100;
    assign weights1[4][150] = 16'b1111111111111011;
    assign weights1[4][151] = 16'b0000000000010010;
    assign weights1[4][152] = 16'b1111111111101111;
    assign weights1[4][153] = 16'b1111111111111000;
    assign weights1[4][154] = 16'b1111111111111110;
    assign weights1[4][155] = 16'b1111111111101110;
    assign weights1[4][156] = 16'b0000000000000111;
    assign weights1[4][157] = 16'b1111111111111100;
    assign weights1[4][158] = 16'b0000000000000000;
    assign weights1[4][159] = 16'b1111111111011000;
    assign weights1[4][160] = 16'b1111111111110111;
    assign weights1[4][161] = 16'b1111111111100001;
    assign weights1[4][162] = 16'b1111111111110010;
    assign weights1[4][163] = 16'b1111111111010101;
    assign weights1[4][164] = 16'b1111111111111110;
    assign weights1[4][165] = 16'b1111111111111100;
    assign weights1[4][166] = 16'b1111111111111001;
    assign weights1[4][167] = 16'b1111111111111000;
    assign weights1[4][168] = 16'b1111111111111110;
    assign weights1[4][169] = 16'b1111111111111111;
    assign weights1[4][170] = 16'b0000000000000000;
    assign weights1[4][171] = 16'b0000000000000001;
    assign weights1[4][172] = 16'b1111111111110011;
    assign weights1[4][173] = 16'b0000000000000100;
    assign weights1[4][174] = 16'b1111111111101110;
    assign weights1[4][175] = 16'b0000000000000101;
    assign weights1[4][176] = 16'b1111111111110011;
    assign weights1[4][177] = 16'b1111111111111000;
    assign weights1[4][178] = 16'b0000000000000100;
    assign weights1[4][179] = 16'b1111111111011010;
    assign weights1[4][180] = 16'b1111111111111100;
    assign weights1[4][181] = 16'b1111111111110111;
    assign weights1[4][182] = 16'b0000000000001000;
    assign weights1[4][183] = 16'b1111111111100101;
    assign weights1[4][184] = 16'b0000000000000110;
    assign weights1[4][185] = 16'b0000000000000110;
    assign weights1[4][186] = 16'b1111111111101100;
    assign weights1[4][187] = 16'b1111111111111011;
    assign weights1[4][188] = 16'b1111111111100111;
    assign weights1[4][189] = 16'b1111111111110100;
    assign weights1[4][190] = 16'b1111111111101100;
    assign weights1[4][191] = 16'b1111111111011100;
    assign weights1[4][192] = 16'b1111111111101110;
    assign weights1[4][193] = 16'b1111111111011110;
    assign weights1[4][194] = 16'b1111111111100001;
    assign weights1[4][195] = 16'b1111111111101111;
    assign weights1[4][196] = 16'b1111111111111111;
    assign weights1[4][197] = 16'b0000000000000011;
    assign weights1[4][198] = 16'b0000000000001011;
    assign weights1[4][199] = 16'b1111111111101010;
    assign weights1[4][200] = 16'b1111111111101110;
    assign weights1[4][201] = 16'b1111111111101001;
    assign weights1[4][202] = 16'b1111111111111101;
    assign weights1[4][203] = 16'b1111111111110010;
    assign weights1[4][204] = 16'b0000000000011101;
    assign weights1[4][205] = 16'b0000000000000010;
    assign weights1[4][206] = 16'b1111111111011100;
    assign weights1[4][207] = 16'b1111111111110011;
    assign weights1[4][208] = 16'b1111111111110111;
    assign weights1[4][209] = 16'b1111111111111101;
    assign weights1[4][210] = 16'b1111111111101011;
    assign weights1[4][211] = 16'b1111111111101011;
    assign weights1[4][212] = 16'b1111111111111001;
    assign weights1[4][213] = 16'b1111111111011011;
    assign weights1[4][214] = 16'b1111111111101111;
    assign weights1[4][215] = 16'b1111111111101000;
    assign weights1[4][216] = 16'b1111111111101111;
    assign weights1[4][217] = 16'b1111111111111111;
    assign weights1[4][218] = 16'b1111111111101101;
    assign weights1[4][219] = 16'b1111111111011110;
    assign weights1[4][220] = 16'b1111111111101010;
    assign weights1[4][221] = 16'b1111111111010110;
    assign weights1[4][222] = 16'b1111111111110000;
    assign weights1[4][223] = 16'b1111111111011111;
    assign weights1[4][224] = 16'b1111111111111111;
    assign weights1[4][225] = 16'b1111111111111011;
    assign weights1[4][226] = 16'b1111111111111110;
    assign weights1[4][227] = 16'b1111111111111001;
    assign weights1[4][228] = 16'b1111111111110111;
    assign weights1[4][229] = 16'b0000000000010110;
    assign weights1[4][230] = 16'b1111111111110100;
    assign weights1[4][231] = 16'b1111111111101000;
    assign weights1[4][232] = 16'b1111111111100101;
    assign weights1[4][233] = 16'b1111111111100010;
    assign weights1[4][234] = 16'b1111111111111111;
    assign weights1[4][235] = 16'b0000000000001000;
    assign weights1[4][236] = 16'b1111111111101100;
    assign weights1[4][237] = 16'b1111111111101110;
    assign weights1[4][238] = 16'b0000000000000011;
    assign weights1[4][239] = 16'b0000000000011110;
    assign weights1[4][240] = 16'b1111111111101111;
    assign weights1[4][241] = 16'b1111111111111000;
    assign weights1[4][242] = 16'b1111111111100010;
    assign weights1[4][243] = 16'b0000000000001111;
    assign weights1[4][244] = 16'b1111111111100001;
    assign weights1[4][245] = 16'b1111111111111100;
    assign weights1[4][246] = 16'b1111111111101111;
    assign weights1[4][247] = 16'b1111111111101011;
    assign weights1[4][248] = 16'b1111111111100100;
    assign weights1[4][249] = 16'b1111111111100101;
    assign weights1[4][250] = 16'b1111111111101000;
    assign weights1[4][251] = 16'b1111111111100001;
    assign weights1[4][252] = 16'b0000000000000001;
    assign weights1[4][253] = 16'b1111111111111100;
    assign weights1[4][254] = 16'b1111111111110111;
    assign weights1[4][255] = 16'b1111111111110001;
    assign weights1[4][256] = 16'b1111111111010111;
    assign weights1[4][257] = 16'b1111111111101100;
    assign weights1[4][258] = 16'b1111111111010101;
    assign weights1[4][259] = 16'b0000000000000000;
    assign weights1[4][260] = 16'b1111111111010001;
    assign weights1[4][261] = 16'b1111111111110000;
    assign weights1[4][262] = 16'b1111111111010110;
    assign weights1[4][263] = 16'b1111111111101101;
    assign weights1[4][264] = 16'b1111111111001110;
    assign weights1[4][265] = 16'b1111111111010100;
    assign weights1[4][266] = 16'b1111111111100010;
    assign weights1[4][267] = 16'b1111111111100111;
    assign weights1[4][268] = 16'b1111111111101110;
    assign weights1[4][269] = 16'b1111111111111111;
    assign weights1[4][270] = 16'b1111111111110111;
    assign weights1[4][271] = 16'b1111111111110111;
    assign weights1[4][272] = 16'b1111111111100001;
    assign weights1[4][273] = 16'b1111111111111011;
    assign weights1[4][274] = 16'b0000000000000000;
    assign weights1[4][275] = 16'b1111111111101110;
    assign weights1[4][276] = 16'b1111111111100110;
    assign weights1[4][277] = 16'b1111111111101101;
    assign weights1[4][278] = 16'b1111111111100100;
    assign weights1[4][279] = 16'b1111111111011011;
    assign weights1[4][280] = 16'b1111111111111011;
    assign weights1[4][281] = 16'b1111111111110001;
    assign weights1[4][282] = 16'b1111111111101101;
    assign weights1[4][283] = 16'b1111111111001111;
    assign weights1[4][284] = 16'b1111111111011011;
    assign weights1[4][285] = 16'b1111111111001000;
    assign weights1[4][286] = 16'b1111111111011011;
    assign weights1[4][287] = 16'b1111111111100100;
    assign weights1[4][288] = 16'b1111111110111100;
    assign weights1[4][289] = 16'b1111111111010110;
    assign weights1[4][290] = 16'b1111111111000000;
    assign weights1[4][291] = 16'b1111111111001001;
    assign weights1[4][292] = 16'b1111111111011111;
    assign weights1[4][293] = 16'b1111111111011001;
    assign weights1[4][294] = 16'b1111111111011001;
    assign weights1[4][295] = 16'b1111111111011000;
    assign weights1[4][296] = 16'b1111111111001110;
    assign weights1[4][297] = 16'b1111111111110011;
    assign weights1[4][298] = 16'b1111111111101001;
    assign weights1[4][299] = 16'b1111111111010101;
    assign weights1[4][300] = 16'b1111111111011010;
    assign weights1[4][301] = 16'b1111111111110000;
    assign weights1[4][302] = 16'b1111111111100110;
    assign weights1[4][303] = 16'b1111111111010011;
    assign weights1[4][304] = 16'b1111111111100111;
    assign weights1[4][305] = 16'b1111111111011111;
    assign weights1[4][306] = 16'b1111111111100001;
    assign weights1[4][307] = 16'b1111111111011101;
    assign weights1[4][308] = 16'b1111111111111100;
    assign weights1[4][309] = 16'b1111111111101000;
    assign weights1[4][310] = 16'b1111111111011100;
    assign weights1[4][311] = 16'b1111111111010001;
    assign weights1[4][312] = 16'b1111111111100010;
    assign weights1[4][313] = 16'b1111111111001011;
    assign weights1[4][314] = 16'b1111111111010011;
    assign weights1[4][315] = 16'b1111111111001101;
    assign weights1[4][316] = 16'b1111111111000100;
    assign weights1[4][317] = 16'b1111111111010100;
    assign weights1[4][318] = 16'b1111111111000010;
    assign weights1[4][319] = 16'b1111111111001010;
    assign weights1[4][320] = 16'b1111111111010000;
    assign weights1[4][321] = 16'b1111111111010000;
    assign weights1[4][322] = 16'b1111111111011000;
    assign weights1[4][323] = 16'b1111111111000010;
    assign weights1[4][324] = 16'b1111111111011010;
    assign weights1[4][325] = 16'b1111111111001100;
    assign weights1[4][326] = 16'b1111111111010100;
    assign weights1[4][327] = 16'b1111111111100010;
    assign weights1[4][328] = 16'b1111111111101111;
    assign weights1[4][329] = 16'b1111111111001101;
    assign weights1[4][330] = 16'b1111111111010111;
    assign weights1[4][331] = 16'b1111111111011001;
    assign weights1[4][332] = 16'b1111111111100100;
    assign weights1[4][333] = 16'b1111111111011100;
    assign weights1[4][334] = 16'b1111111111100010;
    assign weights1[4][335] = 16'b1111111111011001;
    assign weights1[4][336] = 16'b1111111111111011;
    assign weights1[4][337] = 16'b1111111111100110;
    assign weights1[4][338] = 16'b1111111111011011;
    assign weights1[4][339] = 16'b1111111111100110;
    assign weights1[4][340] = 16'b1111111111011001;
    assign weights1[4][341] = 16'b1111111111010001;
    assign weights1[4][342] = 16'b1111111111100100;
    assign weights1[4][343] = 16'b1111111110111011;
    assign weights1[4][344] = 16'b1111111111001101;
    assign weights1[4][345] = 16'b1111111110110111;
    assign weights1[4][346] = 16'b1111111110101011;
    assign weights1[4][347] = 16'b1111111111010001;
    assign weights1[4][348] = 16'b1111111110101111;
    assign weights1[4][349] = 16'b1111111111001001;
    assign weights1[4][350] = 16'b1111111111000100;
    assign weights1[4][351] = 16'b1111111111000111;
    assign weights1[4][352] = 16'b1111111110110100;
    assign weights1[4][353] = 16'b1111111111010101;
    assign weights1[4][354] = 16'b1111111111010100;
    assign weights1[4][355] = 16'b1111111111011110;
    assign weights1[4][356] = 16'b1111111111101001;
    assign weights1[4][357] = 16'b1111111111011011;
    assign weights1[4][358] = 16'b1111111111001001;
    assign weights1[4][359] = 16'b1111111111010110;
    assign weights1[4][360] = 16'b1111111111011011;
    assign weights1[4][361] = 16'b1111111111011111;
    assign weights1[4][362] = 16'b1111111111100011;
    assign weights1[4][363] = 16'b1111111111100001;
    assign weights1[4][364] = 16'b1111111111111101;
    assign weights1[4][365] = 16'b1111111111101101;
    assign weights1[4][366] = 16'b1111111111011111;
    assign weights1[4][367] = 16'b1111111111101011;
    assign weights1[4][368] = 16'b1111111111001111;
    assign weights1[4][369] = 16'b1111111111010111;
    assign weights1[4][370] = 16'b1111111111010001;
    assign weights1[4][371] = 16'b1111111111000101;
    assign weights1[4][372] = 16'b1111111111100000;
    assign weights1[4][373] = 16'b1111111111000000;
    assign weights1[4][374] = 16'b1111111111010000;
    assign weights1[4][375] = 16'b1111111111010001;
    assign weights1[4][376] = 16'b1111111111001011;
    assign weights1[4][377] = 16'b1111111111001110;
    assign weights1[4][378] = 16'b1111111111000010;
    assign weights1[4][379] = 16'b1111111111001000;
    assign weights1[4][380] = 16'b1111111111000110;
    assign weights1[4][381] = 16'b1111111111010110;
    assign weights1[4][382] = 16'b1111111110111000;
    assign weights1[4][383] = 16'b1111111111001101;
    assign weights1[4][384] = 16'b1111111111011010;
    assign weights1[4][385] = 16'b1111111111010100;
    assign weights1[4][386] = 16'b1111111111011001;
    assign weights1[4][387] = 16'b1111111111100001;
    assign weights1[4][388] = 16'b1111111111100110;
    assign weights1[4][389] = 16'b1111111111100101;
    assign weights1[4][390] = 16'b1111111111100101;
    assign weights1[4][391] = 16'b1111111111010111;
    assign weights1[4][392] = 16'b1111111111111110;
    assign weights1[4][393] = 16'b1111111111111000;
    assign weights1[4][394] = 16'b1111111111110000;
    assign weights1[4][395] = 16'b1111111111101010;
    assign weights1[4][396] = 16'b1111111111100110;
    assign weights1[4][397] = 16'b1111111111011111;
    assign weights1[4][398] = 16'b1111111111101011;
    assign weights1[4][399] = 16'b1111111111100110;
    assign weights1[4][400] = 16'b1111111111111001;
    assign weights1[4][401] = 16'b1111111111011101;
    assign weights1[4][402] = 16'b1111111111101110;
    assign weights1[4][403] = 16'b1111111111100111;
    assign weights1[4][404] = 16'b1111111111010000;
    assign weights1[4][405] = 16'b1111111111100011;
    assign weights1[4][406] = 16'b1111111111000001;
    assign weights1[4][407] = 16'b1111111111001000;
    assign weights1[4][408] = 16'b1111111111001001;
    assign weights1[4][409] = 16'b1111111110111000;
    assign weights1[4][410] = 16'b1111111110111011;
    assign weights1[4][411] = 16'b1111111111001111;
    assign weights1[4][412] = 16'b1111111111001011;
    assign weights1[4][413] = 16'b1111111111011001;
    assign weights1[4][414] = 16'b1111111111010100;
    assign weights1[4][415] = 16'b1111111111010110;
    assign weights1[4][416] = 16'b1111111111001010;
    assign weights1[4][417] = 16'b1111111111010111;
    assign weights1[4][418] = 16'b1111111111010101;
    assign weights1[4][419] = 16'b1111111111010110;
    assign weights1[4][420] = 16'b1111111111111101;
    assign weights1[4][421] = 16'b0000000000000110;
    assign weights1[4][422] = 16'b1111111111110010;
    assign weights1[4][423] = 16'b0000000000000010;
    assign weights1[4][424] = 16'b1111111111110100;
    assign weights1[4][425] = 16'b1111111111010001;
    assign weights1[4][426] = 16'b0000000000001001;
    assign weights1[4][427] = 16'b1111111111011110;
    assign weights1[4][428] = 16'b0000000000000111;
    assign weights1[4][429] = 16'b1111111111111101;
    assign weights1[4][430] = 16'b1111111111110001;
    assign weights1[4][431] = 16'b1111111111110110;
    assign weights1[4][432] = 16'b1111111111110000;
    assign weights1[4][433] = 16'b1111111111010110;
    assign weights1[4][434] = 16'b1111111111101110;
    assign weights1[4][435] = 16'b1111111111100010;
    assign weights1[4][436] = 16'b1111111111010101;
    assign weights1[4][437] = 16'b1111111111011011;
    assign weights1[4][438] = 16'b1111111111000000;
    assign weights1[4][439] = 16'b1111111110111101;
    assign weights1[4][440] = 16'b1111111111001010;
    assign weights1[4][441] = 16'b1111111111001100;
    assign weights1[4][442] = 16'b1111111111001111;
    assign weights1[4][443] = 16'b1111111110110001;
    assign weights1[4][444] = 16'b1111111111001010;
    assign weights1[4][445] = 16'b1111111111001000;
    assign weights1[4][446] = 16'b1111111111010110;
    assign weights1[4][447] = 16'b1111111111011001;
    assign weights1[4][448] = 16'b0000000000011000;
    assign weights1[4][449] = 16'b0000000000001110;
    assign weights1[4][450] = 16'b0000000000010110;
    assign weights1[4][451] = 16'b0000000000011011;
    assign weights1[4][452] = 16'b0000000000001101;
    assign weights1[4][453] = 16'b1111111111111010;
    assign weights1[4][454] = 16'b0000000000000100;
    assign weights1[4][455] = 16'b0000000000010001;
    assign weights1[4][456] = 16'b0000000000001100;
    assign weights1[4][457] = 16'b0000000000001001;
    assign weights1[4][458] = 16'b1111111111110101;
    assign weights1[4][459] = 16'b1111111111001111;
    assign weights1[4][460] = 16'b0000000000000100;
    assign weights1[4][461] = 16'b1111111111110110;
    assign weights1[4][462] = 16'b1111111111101110;
    assign weights1[4][463] = 16'b1111111111110101;
    assign weights1[4][464] = 16'b1111111111110111;
    assign weights1[4][465] = 16'b1111111111100001;
    assign weights1[4][466] = 16'b1111111111100001;
    assign weights1[4][467] = 16'b1111111111101000;
    assign weights1[4][468] = 16'b1111111111011101;
    assign weights1[4][469] = 16'b1111111110110110;
    assign weights1[4][470] = 16'b1111111110110010;
    assign weights1[4][471] = 16'b1111111111000001;
    assign weights1[4][472] = 16'b1111111110110101;
    assign weights1[4][473] = 16'b1111111111010000;
    assign weights1[4][474] = 16'b1111111111011011;
    assign weights1[4][475] = 16'b1111111111011001;
    assign weights1[4][476] = 16'b0000000000011111;
    assign weights1[4][477] = 16'b0000000000010110;
    assign weights1[4][478] = 16'b0000000000101011;
    assign weights1[4][479] = 16'b0000000000101000;
    assign weights1[4][480] = 16'b0000000000010110;
    assign weights1[4][481] = 16'b0000000000111010;
    assign weights1[4][482] = 16'b0000000000110100;
    assign weights1[4][483] = 16'b0000000000110001;
    assign weights1[4][484] = 16'b0000000000101100;
    assign weights1[4][485] = 16'b0000000000001111;
    assign weights1[4][486] = 16'b0000000000011100;
    assign weights1[4][487] = 16'b1111111111111111;
    assign weights1[4][488] = 16'b0000000000000101;
    assign weights1[4][489] = 16'b0000000000001010;
    assign weights1[4][490] = 16'b1111111111111110;
    assign weights1[4][491] = 16'b0000000000001101;
    assign weights1[4][492] = 16'b1111111111111010;
    assign weights1[4][493] = 16'b1111111111110010;
    assign weights1[4][494] = 16'b1111111111100100;
    assign weights1[4][495] = 16'b0000000000000010;
    assign weights1[4][496] = 16'b1111111111111000;
    assign weights1[4][497] = 16'b1111111111101110;
    assign weights1[4][498] = 16'b1111111111110110;
    assign weights1[4][499] = 16'b1111111111101100;
    assign weights1[4][500] = 16'b1111111111110000;
    assign weights1[4][501] = 16'b1111111111110011;
    assign weights1[4][502] = 16'b1111111111100101;
    assign weights1[4][503] = 16'b1111111111110011;
    assign weights1[4][504] = 16'b0000000000011110;
    assign weights1[4][505] = 16'b0000000000101000;
    assign weights1[4][506] = 16'b0000000000101010;
    assign weights1[4][507] = 16'b0000000000100000;
    assign weights1[4][508] = 16'b0000000000111111;
    assign weights1[4][509] = 16'b0000000001000101;
    assign weights1[4][510] = 16'b0000000000101111;
    assign weights1[4][511] = 16'b0000000001001011;
    assign weights1[4][512] = 16'b0000000000110101;
    assign weights1[4][513] = 16'b0000000000110111;
    assign weights1[4][514] = 16'b0000000000011001;
    assign weights1[4][515] = 16'b0000000000110011;
    assign weights1[4][516] = 16'b0000000001001111;
    assign weights1[4][517] = 16'b0000000000011001;
    assign weights1[4][518] = 16'b0000000000100011;
    assign weights1[4][519] = 16'b0000000000010111;
    assign weights1[4][520] = 16'b0000000001000001;
    assign weights1[4][521] = 16'b0000000000010101;
    assign weights1[4][522] = 16'b0000000000011100;
    assign weights1[4][523] = 16'b0000000000101000;
    assign weights1[4][524] = 16'b0000000000011001;
    assign weights1[4][525] = 16'b0000000000001010;
    assign weights1[4][526] = 16'b0000000000100000;
    assign weights1[4][527] = 16'b0000000000101100;
    assign weights1[4][528] = 16'b0000000000100001;
    assign weights1[4][529] = 16'b0000000000000110;
    assign weights1[4][530] = 16'b1111111111110011;
    assign weights1[4][531] = 16'b0000000000001111;
    assign weights1[4][532] = 16'b0000000000101000;
    assign weights1[4][533] = 16'b0000000000101100;
    assign weights1[4][534] = 16'b0000000000011101;
    assign weights1[4][535] = 16'b0000000000100000;
    assign weights1[4][536] = 16'b0000000000100011;
    assign weights1[4][537] = 16'b0000000000110110;
    assign weights1[4][538] = 16'b0000000000111011;
    assign weights1[4][539] = 16'b0000000000111100;
    assign weights1[4][540] = 16'b0000000001001000;
    assign weights1[4][541] = 16'b0000000001000101;
    assign weights1[4][542] = 16'b0000000001000110;
    assign weights1[4][543] = 16'b0000000001011010;
    assign weights1[4][544] = 16'b0000000001001111;
    assign weights1[4][545] = 16'b0000000001001000;
    assign weights1[4][546] = 16'b0000000000111111;
    assign weights1[4][547] = 16'b0000000001001000;
    assign weights1[4][548] = 16'b0000000000101110;
    assign weights1[4][549] = 16'b0000000000100001;
    assign weights1[4][550] = 16'b0000000000110100;
    assign weights1[4][551] = 16'b0000000000101011;
    assign weights1[4][552] = 16'b0000000000011101;
    assign weights1[4][553] = 16'b0000000000011111;
    assign weights1[4][554] = 16'b0000000000100110;
    assign weights1[4][555] = 16'b0000000000110001;
    assign weights1[4][556] = 16'b0000000000110100;
    assign weights1[4][557] = 16'b0000000000011110;
    assign weights1[4][558] = 16'b0000000000011010;
    assign weights1[4][559] = 16'b0000000000100111;
    assign weights1[4][560] = 16'b0000000000010101;
    assign weights1[4][561] = 16'b0000000000011111;
    assign weights1[4][562] = 16'b0000000000011110;
    assign weights1[4][563] = 16'b0000000000111101;
    assign weights1[4][564] = 16'b0000000000111010;
    assign weights1[4][565] = 16'b0000000000101101;
    assign weights1[4][566] = 16'b0000000000110111;
    assign weights1[4][567] = 16'b0000000000111001;
    assign weights1[4][568] = 16'b0000000000101101;
    assign weights1[4][569] = 16'b0000000000101111;
    assign weights1[4][570] = 16'b0000000000110110;
    assign weights1[4][571] = 16'b0000000001001011;
    assign weights1[4][572] = 16'b0000000001001100;
    assign weights1[4][573] = 16'b0000000001001100;
    assign weights1[4][574] = 16'b0000000001011101;
    assign weights1[4][575] = 16'b0000000000110110;
    assign weights1[4][576] = 16'b0000000001000011;
    assign weights1[4][577] = 16'b0000000000110001;
    assign weights1[4][578] = 16'b0000000001001000;
    assign weights1[4][579] = 16'b0000000000111010;
    assign weights1[4][580] = 16'b0000000001000101;
    assign weights1[4][581] = 16'b0000000000100010;
    assign weights1[4][582] = 16'b0000000000100111;
    assign weights1[4][583] = 16'b0000000000110000;
    assign weights1[4][584] = 16'b0000000000111101;
    assign weights1[4][585] = 16'b0000000000101011;
    assign weights1[4][586] = 16'b0000000000110001;
    assign weights1[4][587] = 16'b0000000000100100;
    assign weights1[4][588] = 16'b0000000000000111;
    assign weights1[4][589] = 16'b0000000000010001;
    assign weights1[4][590] = 16'b0000000000101011;
    assign weights1[4][591] = 16'b0000000000110010;
    assign weights1[4][592] = 16'b0000000000100000;
    assign weights1[4][593] = 16'b0000000000100001;
    assign weights1[4][594] = 16'b0000000000100110;
    assign weights1[4][595] = 16'b0000000000100110;
    assign weights1[4][596] = 16'b0000000000100111;
    assign weights1[4][597] = 16'b0000000000100000;
    assign weights1[4][598] = 16'b0000000000101100;
    assign weights1[4][599] = 16'b0000000000011100;
    assign weights1[4][600] = 16'b0000000000010011;
    assign weights1[4][601] = 16'b0000000000100111;
    assign weights1[4][602] = 16'b0000000000101110;
    assign weights1[4][603] = 16'b0000000000101001;
    assign weights1[4][604] = 16'b0000000000111100;
    assign weights1[4][605] = 16'b0000000001010001;
    assign weights1[4][606] = 16'b0000000001000111;
    assign weights1[4][607] = 16'b0000000001001011;
    assign weights1[4][608] = 16'b0000000000101110;
    assign weights1[4][609] = 16'b0000000000111011;
    assign weights1[4][610] = 16'b0000000000110000;
    assign weights1[4][611] = 16'b0000000001100000;
    assign weights1[4][612] = 16'b0000000001001110;
    assign weights1[4][613] = 16'b0000000001000010;
    assign weights1[4][614] = 16'b0000000000101100;
    assign weights1[4][615] = 16'b0000000000100001;
    assign weights1[4][616] = 16'b0000000000001011;
    assign weights1[4][617] = 16'b0000000000001110;
    assign weights1[4][618] = 16'b0000000000001110;
    assign weights1[4][619] = 16'b0000000000010100;
    assign weights1[4][620] = 16'b0000000000010110;
    assign weights1[4][621] = 16'b0000000000100111;
    assign weights1[4][622] = 16'b0000000000010000;
    assign weights1[4][623] = 16'b0000000000100000;
    assign weights1[4][624] = 16'b0000000000110000;
    assign weights1[4][625] = 16'b0000000000010111;
    assign weights1[4][626] = 16'b1111111111111001;
    assign weights1[4][627] = 16'b0000000000010101;
    assign weights1[4][628] = 16'b0000000000010110;
    assign weights1[4][629] = 16'b0000000000001011;
    assign weights1[4][630] = 16'b0000000000011001;
    assign weights1[4][631] = 16'b0000000000100100;
    assign weights1[4][632] = 16'b0000000000011110;
    assign weights1[4][633] = 16'b0000000000101101;
    assign weights1[4][634] = 16'b0000000000111001;
    assign weights1[4][635] = 16'b0000000001000100;
    assign weights1[4][636] = 16'b0000000000110011;
    assign weights1[4][637] = 16'b0000000000111100;
    assign weights1[4][638] = 16'b0000000001000110;
    assign weights1[4][639] = 16'b0000000000111011;
    assign weights1[4][640] = 16'b0000000001000100;
    assign weights1[4][641] = 16'b0000000000110111;
    assign weights1[4][642] = 16'b0000000000100111;
    assign weights1[4][643] = 16'b0000000000011110;
    assign weights1[4][644] = 16'b0000000000000010;
    assign weights1[4][645] = 16'b0000000000000101;
    assign weights1[4][646] = 16'b0000000000001011;
    assign weights1[4][647] = 16'b0000000000001100;
    assign weights1[4][648] = 16'b0000000000001000;
    assign weights1[4][649] = 16'b0000000000011000;
    assign weights1[4][650] = 16'b0000000000011010;
    assign weights1[4][651] = 16'b0000000000001100;
    assign weights1[4][652] = 16'b0000000000100000;
    assign weights1[4][653] = 16'b0000000000100000;
    assign weights1[4][654] = 16'b0000000000011011;
    assign weights1[4][655] = 16'b0000000000100101;
    assign weights1[4][656] = 16'b0000000000100011;
    assign weights1[4][657] = 16'b0000000000000110;
    assign weights1[4][658] = 16'b0000000000001011;
    assign weights1[4][659] = 16'b0000000000010111;
    assign weights1[4][660] = 16'b0000000000010111;
    assign weights1[4][661] = 16'b0000000000000110;
    assign weights1[4][662] = 16'b0000000000100111;
    assign weights1[4][663] = 16'b0000000000111100;
    assign weights1[4][664] = 16'b0000000001000010;
    assign weights1[4][665] = 16'b0000000000111111;
    assign weights1[4][666] = 16'b0000000001000010;
    assign weights1[4][667] = 16'b0000000000100010;
    assign weights1[4][668] = 16'b0000000000111110;
    assign weights1[4][669] = 16'b0000000000110011;
    assign weights1[4][670] = 16'b0000000000011001;
    assign weights1[4][671] = 16'b0000000000010000;
    assign weights1[4][672] = 16'b0000000000000011;
    assign weights1[4][673] = 16'b0000000000000100;
    assign weights1[4][674] = 16'b0000000000001100;
    assign weights1[4][675] = 16'b0000000000000101;
    assign weights1[4][676] = 16'b0000000000000011;
    assign weights1[4][677] = 16'b0000000000000100;
    assign weights1[4][678] = 16'b0000000000000011;
    assign weights1[4][679] = 16'b0000000000000111;
    assign weights1[4][680] = 16'b0000000000000101;
    assign weights1[4][681] = 16'b0000000000000010;
    assign weights1[4][682] = 16'b1111111111110001;
    assign weights1[4][683] = 16'b1111111111111011;
    assign weights1[4][684] = 16'b0000000000010011;
    assign weights1[4][685] = 16'b0000000000100110;
    assign weights1[4][686] = 16'b0000000000010101;
    assign weights1[4][687] = 16'b0000000000000111;
    assign weights1[4][688] = 16'b0000000000011000;
    assign weights1[4][689] = 16'b1111111111111010;
    assign weights1[4][690] = 16'b1111111111111100;
    assign weights1[4][691] = 16'b0000000000000001;
    assign weights1[4][692] = 16'b0000000000010001;
    assign weights1[4][693] = 16'b0000000000001000;
    assign weights1[4][694] = 16'b0000000000100100;
    assign weights1[4][695] = 16'b0000000000010111;
    assign weights1[4][696] = 16'b0000000000110011;
    assign weights1[4][697] = 16'b0000000000110011;
    assign weights1[4][698] = 16'b0000000000010100;
    assign weights1[4][699] = 16'b0000000000001001;
    assign weights1[4][700] = 16'b0000000000000000;
    assign weights1[4][701] = 16'b0000000000000001;
    assign weights1[4][702] = 16'b1111111111110110;
    assign weights1[4][703] = 16'b1111111111101101;
    assign weights1[4][704] = 16'b1111111111101101;
    assign weights1[4][705] = 16'b1111111111111100;
    assign weights1[4][706] = 16'b0000000000000000;
    assign weights1[4][707] = 16'b1111111111101011;
    assign weights1[4][708] = 16'b0000000000001000;
    assign weights1[4][709] = 16'b0000000000000001;
    assign weights1[4][710] = 16'b0000000000000101;
    assign weights1[4][711] = 16'b1111111111111111;
    assign weights1[4][712] = 16'b1111111111101111;
    assign weights1[4][713] = 16'b1111111111111111;
    assign weights1[4][714] = 16'b1111111111111101;
    assign weights1[4][715] = 16'b0000000000000110;
    assign weights1[4][716] = 16'b0000000000000110;
    assign weights1[4][717] = 16'b1111111111110110;
    assign weights1[4][718] = 16'b0000000000000000;
    assign weights1[4][719] = 16'b1111111111101000;
    assign weights1[4][720] = 16'b0000000000000100;
    assign weights1[4][721] = 16'b1111111111110001;
    assign weights1[4][722] = 16'b0000000000000000;
    assign weights1[4][723] = 16'b0000000000001111;
    assign weights1[4][724] = 16'b0000000000100101;
    assign weights1[4][725] = 16'b0000000000100011;
    assign weights1[4][726] = 16'b0000000000001001;
    assign weights1[4][727] = 16'b0000000000000100;
    assign weights1[4][728] = 16'b1111111111111110;
    assign weights1[4][729] = 16'b1111111111111111;
    assign weights1[4][730] = 16'b1111111111110111;
    assign weights1[4][731] = 16'b1111111111110000;
    assign weights1[4][732] = 16'b1111111111110011;
    assign weights1[4][733] = 16'b1111111111110001;
    assign weights1[4][734] = 16'b1111111111110010;
    assign weights1[4][735] = 16'b1111111111110011;
    assign weights1[4][736] = 16'b1111111111110011;
    assign weights1[4][737] = 16'b1111111111101111;
    assign weights1[4][738] = 16'b1111111111101011;
    assign weights1[4][739] = 16'b1111111111101001;
    assign weights1[4][740] = 16'b0000000000000110;
    assign weights1[4][741] = 16'b1111111111111011;
    assign weights1[4][742] = 16'b0000000000010111;
    assign weights1[4][743] = 16'b0000000000000011;
    assign weights1[4][744] = 16'b1111111111111010;
    assign weights1[4][745] = 16'b1111111111111010;
    assign weights1[4][746] = 16'b1111111111111001;
    assign weights1[4][747] = 16'b1111111111111001;
    assign weights1[4][748] = 16'b0000000000001110;
    assign weights1[4][749] = 16'b1111111111101110;
    assign weights1[4][750] = 16'b0000000000001001;
    assign weights1[4][751] = 16'b0000000000000110;
    assign weights1[4][752] = 16'b0000000000001001;
    assign weights1[4][753] = 16'b0000000000010000;
    assign weights1[4][754] = 16'b0000000000000001;
    assign weights1[4][755] = 16'b0000000000000000;
    assign weights1[4][756] = 16'b0000000000000001;
    assign weights1[4][757] = 16'b1111111111111100;
    assign weights1[4][758] = 16'b1111111111111100;
    assign weights1[4][759] = 16'b1111111111110011;
    assign weights1[4][760] = 16'b1111111111111010;
    assign weights1[4][761] = 16'b1111111111101111;
    assign weights1[4][762] = 16'b1111111111101001;
    assign weights1[4][763] = 16'b1111111111101001;
    assign weights1[4][764] = 16'b1111111111100110;
    assign weights1[4][765] = 16'b1111111111100011;
    assign weights1[4][766] = 16'b1111111111101111;
    assign weights1[4][767] = 16'b1111111111101101;
    assign weights1[4][768] = 16'b1111111111110001;
    assign weights1[4][769] = 16'b1111111111111000;
    assign weights1[4][770] = 16'b1111111111110001;
    assign weights1[4][771] = 16'b1111111111100101;
    assign weights1[4][772] = 16'b1111111111101001;
    assign weights1[4][773] = 16'b1111111111111111;
    assign weights1[4][774] = 16'b0000000000000101;
    assign weights1[4][775] = 16'b0000000000001101;
    assign weights1[4][776] = 16'b1111111111110101;
    assign weights1[4][777] = 16'b0000000000000110;
    assign weights1[4][778] = 16'b0000000000000011;
    assign weights1[4][779] = 16'b0000000000000100;
    assign weights1[4][780] = 16'b1111111111111101;
    assign weights1[4][781] = 16'b1111111111111111;
    assign weights1[4][782] = 16'b1111111111111011;
    assign weights1[4][783] = 16'b0000000000000001;
    assign weights1[5][0] = 16'b0000000000000001;
    assign weights1[5][1] = 16'b0000000000000001;
    assign weights1[5][2] = 16'b0000000000000000;
    assign weights1[5][3] = 16'b0000000000000101;
    assign weights1[5][4] = 16'b0000000000001001;
    assign weights1[5][5] = 16'b0000000000001101;
    assign weights1[5][6] = 16'b0000000000000110;
    assign weights1[5][7] = 16'b0000000000010110;
    assign weights1[5][8] = 16'b0000000000100101;
    assign weights1[5][9] = 16'b0000000000001100;
    assign weights1[5][10] = 16'b0000000000000011;
    assign weights1[5][11] = 16'b1111111111110111;
    assign weights1[5][12] = 16'b1111111111101110;
    assign weights1[5][13] = 16'b1111111111010011;
    assign weights1[5][14] = 16'b1111111111011110;
    assign weights1[5][15] = 16'b1111111111011011;
    assign weights1[5][16] = 16'b1111111111011000;
    assign weights1[5][17] = 16'b1111111111100011;
    assign weights1[5][18] = 16'b1111111111101010;
    assign weights1[5][19] = 16'b1111111111110010;
    assign weights1[5][20] = 16'b1111111111111001;
    assign weights1[5][21] = 16'b1111111111111010;
    assign weights1[5][22] = 16'b1111111111111011;
    assign weights1[5][23] = 16'b0000000000000000;
    assign weights1[5][24] = 16'b0000000000000000;
    assign weights1[5][25] = 16'b0000000000000000;
    assign weights1[5][26] = 16'b0000000000000000;
    assign weights1[5][27] = 16'b0000000000000000;
    assign weights1[5][28] = 16'b0000000000000010;
    assign weights1[5][29] = 16'b0000000000000100;
    assign weights1[5][30] = 16'b0000000000001010;
    assign weights1[5][31] = 16'b0000000000000101;
    assign weights1[5][32] = 16'b0000000000010010;
    assign weights1[5][33] = 16'b0000000000011111;
    assign weights1[5][34] = 16'b0000000000100100;
    assign weights1[5][35] = 16'b0000000000100001;
    assign weights1[5][36] = 16'b0000000000100001;
    assign weights1[5][37] = 16'b0000000000000111;
    assign weights1[5][38] = 16'b0000000000000101;
    assign weights1[5][39] = 16'b1111111111111101;
    assign weights1[5][40] = 16'b1111111111110001;
    assign weights1[5][41] = 16'b1111111111101000;
    assign weights1[5][42] = 16'b1111111111100111;
    assign weights1[5][43] = 16'b1111111111100010;
    assign weights1[5][44] = 16'b1111111111011100;
    assign weights1[5][45] = 16'b1111111111011001;
    assign weights1[5][46] = 16'b1111111111011011;
    assign weights1[5][47] = 16'b1111111111100001;
    assign weights1[5][48] = 16'b1111111111110011;
    assign weights1[5][49] = 16'b1111111111110101;
    assign weights1[5][50] = 16'b1111111111111011;
    assign weights1[5][51] = 16'b1111111111111100;
    assign weights1[5][52] = 16'b1111111111111111;
    assign weights1[5][53] = 16'b0000000000000000;
    assign weights1[5][54] = 16'b0000000000000000;
    assign weights1[5][55] = 16'b0000000000000000;
    assign weights1[5][56] = 16'b0000000000000110;
    assign weights1[5][57] = 16'b0000000000001001;
    assign weights1[5][58] = 16'b0000000000001011;
    assign weights1[5][59] = 16'b0000000000010100;
    assign weights1[5][60] = 16'b0000000000010100;
    assign weights1[5][61] = 16'b0000000000100100;
    assign weights1[5][62] = 16'b0000000000100000;
    assign weights1[5][63] = 16'b0000000000010110;
    assign weights1[5][64] = 16'b0000000000010011;
    assign weights1[5][65] = 16'b0000000000001000;
    assign weights1[5][66] = 16'b0000000000001100;
    assign weights1[5][67] = 16'b0000000000001010;
    assign weights1[5][68] = 16'b0000000000000110;
    assign weights1[5][69] = 16'b1111111111101001;
    assign weights1[5][70] = 16'b1111111111100010;
    assign weights1[5][71] = 16'b1111111111100000;
    assign weights1[5][72] = 16'b1111111111101000;
    assign weights1[5][73] = 16'b1111111111001111;
    assign weights1[5][74] = 16'b1111111111000100;
    assign weights1[5][75] = 16'b1111111111010000;
    assign weights1[5][76] = 16'b1111111111011111;
    assign weights1[5][77] = 16'b1111111111110100;
    assign weights1[5][78] = 16'b1111111111111011;
    assign weights1[5][79] = 16'b1111111111111101;
    assign weights1[5][80] = 16'b0000000000000000;
    assign weights1[5][81] = 16'b0000000000000001;
    assign weights1[5][82] = 16'b0000000000000000;
    assign weights1[5][83] = 16'b0000000000000000;
    assign weights1[5][84] = 16'b0000000000001100;
    assign weights1[5][85] = 16'b0000000000011000;
    assign weights1[5][86] = 16'b0000000000011000;
    assign weights1[5][87] = 16'b0000000000001111;
    assign weights1[5][88] = 16'b0000000000100010;
    assign weights1[5][89] = 16'b0000000000011010;
    assign weights1[5][90] = 16'b0000000000100111;
    assign weights1[5][91] = 16'b0000000000100001;
    assign weights1[5][92] = 16'b0000000000010101;
    assign weights1[5][93] = 16'b0000000000000011;
    assign weights1[5][94] = 16'b0000000000010110;
    assign weights1[5][95] = 16'b1111111111111100;
    assign weights1[5][96] = 16'b1111111111100110;
    assign weights1[5][97] = 16'b1111111111100101;
    assign weights1[5][98] = 16'b1111111111100110;
    assign weights1[5][99] = 16'b1111111110111110;
    assign weights1[5][100] = 16'b1111111111100100;
    assign weights1[5][101] = 16'b1111111111010010;
    assign weights1[5][102] = 16'b1111111110110010;
    assign weights1[5][103] = 16'b1111111111001000;
    assign weights1[5][104] = 16'b1111111111100001;
    assign weights1[5][105] = 16'b1111111111110000;
    assign weights1[5][106] = 16'b1111111111110111;
    assign weights1[5][107] = 16'b1111111111111001;
    assign weights1[5][108] = 16'b0000000000000000;
    assign weights1[5][109] = 16'b0000000000000000;
    assign weights1[5][110] = 16'b0000000000000000;
    assign weights1[5][111] = 16'b0000000000000000;
    assign weights1[5][112] = 16'b0000000000001100;
    assign weights1[5][113] = 16'b0000000000011100;
    assign weights1[5][114] = 16'b0000000000010011;
    assign weights1[5][115] = 16'b0000000000010011;
    assign weights1[5][116] = 16'b0000000000010001;
    assign weights1[5][117] = 16'b0000000000010100;
    assign weights1[5][118] = 16'b0000000000010101;
    assign weights1[5][119] = 16'b0000000000011000;
    assign weights1[5][120] = 16'b0000000000011100;
    assign weights1[5][121] = 16'b0000000000001100;
    assign weights1[5][122] = 16'b0000000000010111;
    assign weights1[5][123] = 16'b0000000000011010;
    assign weights1[5][124] = 16'b0000000000010110;
    assign weights1[5][125] = 16'b0000000000011010;
    assign weights1[5][126] = 16'b0000000000000001;
    assign weights1[5][127] = 16'b1111111111100100;
    assign weights1[5][128] = 16'b1111111111000000;
    assign weights1[5][129] = 16'b1111111110101000;
    assign weights1[5][130] = 16'b1111111110100111;
    assign weights1[5][131] = 16'b1111111111000010;
    assign weights1[5][132] = 16'b1111111111011010;
    assign weights1[5][133] = 16'b1111111111101101;
    assign weights1[5][134] = 16'b1111111111110011;
    assign weights1[5][135] = 16'b1111111111110110;
    assign weights1[5][136] = 16'b1111111111111110;
    assign weights1[5][137] = 16'b0000000000000000;
    assign weights1[5][138] = 16'b0000000000000000;
    assign weights1[5][139] = 16'b0000000000000000;
    assign weights1[5][140] = 16'b0000000000001100;
    assign weights1[5][141] = 16'b0000000000011101;
    assign weights1[5][142] = 16'b0000000000010110;
    assign weights1[5][143] = 16'b0000000000011000;
    assign weights1[5][144] = 16'b0000000000001010;
    assign weights1[5][145] = 16'b0000000000011110;
    assign weights1[5][146] = 16'b0000000000001110;
    assign weights1[5][147] = 16'b0000000000010111;
    assign weights1[5][148] = 16'b0000000000010111;
    assign weights1[5][149] = 16'b0000000000000001;
    assign weights1[5][150] = 16'b0000000000011011;
    assign weights1[5][151] = 16'b0000000000010011;
    assign weights1[5][152] = 16'b0000000000001111;
    assign weights1[5][153] = 16'b0000000000010010;
    assign weights1[5][154] = 16'b1111111111111001;
    assign weights1[5][155] = 16'b0000000000000110;
    assign weights1[5][156] = 16'b1111111111111001;
    assign weights1[5][157] = 16'b1111111110110101;
    assign weights1[5][158] = 16'b1111111110101001;
    assign weights1[5][159] = 16'b1111111110101111;
    assign weights1[5][160] = 16'b1111111111011000;
    assign weights1[5][161] = 16'b1111111111110001;
    assign weights1[5][162] = 16'b1111111111110010;
    assign weights1[5][163] = 16'b1111111111110100;
    assign weights1[5][164] = 16'b1111111111111011;
    assign weights1[5][165] = 16'b1111111111111011;
    assign weights1[5][166] = 16'b1111111111111100;
    assign weights1[5][167] = 16'b0000000000000000;
    assign weights1[5][168] = 16'b0000000000001101;
    assign weights1[5][169] = 16'b0000000000010101;
    assign weights1[5][170] = 16'b0000000000011110;
    assign weights1[5][171] = 16'b0000000000011111;
    assign weights1[5][172] = 16'b0000000000010100;
    assign weights1[5][173] = 16'b0000000000011001;
    assign weights1[5][174] = 16'b0000000000011011;
    assign weights1[5][175] = 16'b0000000000101110;
    assign weights1[5][176] = 16'b0000000000010001;
    assign weights1[5][177] = 16'b0000000000001101;
    assign weights1[5][178] = 16'b0000000000100010;
    assign weights1[5][179] = 16'b0000000000100000;
    assign weights1[5][180] = 16'b0000000000001100;
    assign weights1[5][181] = 16'b0000000000010010;
    assign weights1[5][182] = 16'b1111111111110101;
    assign weights1[5][183] = 16'b0000000000000011;
    assign weights1[5][184] = 16'b1111111111110000;
    assign weights1[5][185] = 16'b1111111111000100;
    assign weights1[5][186] = 16'b1111111101111010;
    assign weights1[5][187] = 16'b1111111110010100;
    assign weights1[5][188] = 16'b1111111111011010;
    assign weights1[5][189] = 16'b1111111111101001;
    assign weights1[5][190] = 16'b1111111111101100;
    assign weights1[5][191] = 16'b1111111111110010;
    assign weights1[5][192] = 16'b1111111111110010;
    assign weights1[5][193] = 16'b1111111111110111;
    assign weights1[5][194] = 16'b1111111111111011;
    assign weights1[5][195] = 16'b0000000000000000;
    assign weights1[5][196] = 16'b0000000000010101;
    assign weights1[5][197] = 16'b0000000000100010;
    assign weights1[5][198] = 16'b0000000000101000;
    assign weights1[5][199] = 16'b0000000000010000;
    assign weights1[5][200] = 16'b0000000000001111;
    assign weights1[5][201] = 16'b1111111111110111;
    assign weights1[5][202] = 16'b0000000000000101;
    assign weights1[5][203] = 16'b1111111111101010;
    assign weights1[5][204] = 16'b1111111111111101;
    assign weights1[5][205] = 16'b0000000000010000;
    assign weights1[5][206] = 16'b0000000000010001;
    assign weights1[5][207] = 16'b0000000000110101;
    assign weights1[5][208] = 16'b0000000000011101;
    assign weights1[5][209] = 16'b0000000000000010;
    assign weights1[5][210] = 16'b0000000000010011;
    assign weights1[5][211] = 16'b0000000000001011;
    assign weights1[5][212] = 16'b0000000000001101;
    assign weights1[5][213] = 16'b1111111110111001;
    assign weights1[5][214] = 16'b1111111101100010;
    assign weights1[5][215] = 16'b1111111110010111;
    assign weights1[5][216] = 16'b1111111111010010;
    assign weights1[5][217] = 16'b1111111111101011;
    assign weights1[5][218] = 16'b1111111111101111;
    assign weights1[5][219] = 16'b1111111111101111;
    assign weights1[5][220] = 16'b1111111111110100;
    assign weights1[5][221] = 16'b1111111111110011;
    assign weights1[5][222] = 16'b1111111111111011;
    assign weights1[5][223] = 16'b0000000000000000;
    assign weights1[5][224] = 16'b0000000000011110;
    assign weights1[5][225] = 16'b0000000000100000;
    assign weights1[5][226] = 16'b0000000000000010;
    assign weights1[5][227] = 16'b0000000000001000;
    assign weights1[5][228] = 16'b0000000000000100;
    assign weights1[5][229] = 16'b1111111111111000;
    assign weights1[5][230] = 16'b1111111111111100;
    assign weights1[5][231] = 16'b0000000000001100;
    assign weights1[5][232] = 16'b1111111111110100;
    assign weights1[5][233] = 16'b0000000000000111;
    assign weights1[5][234] = 16'b0000000000111111;
    assign weights1[5][235] = 16'b0000000000100100;
    assign weights1[5][236] = 16'b0000000000101000;
    assign weights1[5][237] = 16'b0000000000110011;
    assign weights1[5][238] = 16'b0000000000101110;
    assign weights1[5][239] = 16'b0000000000001101;
    assign weights1[5][240] = 16'b1111111111101001;
    assign weights1[5][241] = 16'b1111111111010011;
    assign weights1[5][242] = 16'b1111111101110111;
    assign weights1[5][243] = 16'b1111111110101111;
    assign weights1[5][244] = 16'b1111111111001010;
    assign weights1[5][245] = 16'b1111111111011100;
    assign weights1[5][246] = 16'b1111111111100101;
    assign weights1[5][247] = 16'b1111111111101000;
    assign weights1[5][248] = 16'b1111111111101111;
    assign weights1[5][249] = 16'b1111111111110010;
    assign weights1[5][250] = 16'b1111111111110110;
    assign weights1[5][251] = 16'b1111111111111001;
    assign weights1[5][252] = 16'b0000000000010011;
    assign weights1[5][253] = 16'b0000000000010000;
    assign weights1[5][254] = 16'b0000000000010000;
    assign weights1[5][255] = 16'b0000000000000011;
    assign weights1[5][256] = 16'b0000000000000110;
    assign weights1[5][257] = 16'b0000000000001110;
    assign weights1[5][258] = 16'b1111111111110101;
    assign weights1[5][259] = 16'b1111111111101010;
    assign weights1[5][260] = 16'b1111111111101111;
    assign weights1[5][261] = 16'b0000000000011000;
    assign weights1[5][262] = 16'b0000000000101100;
    assign weights1[5][263] = 16'b0000000000011100;
    assign weights1[5][264] = 16'b0000000000101000;
    assign weights1[5][265] = 16'b0000000000111111;
    assign weights1[5][266] = 16'b0000000000101010;
    assign weights1[5][267] = 16'b0000000000011111;
    assign weights1[5][268] = 16'b1111111111010101;
    assign weights1[5][269] = 16'b1111111110110110;
    assign weights1[5][270] = 16'b1111111101111010;
    assign weights1[5][271] = 16'b1111111110111011;
    assign weights1[5][272] = 16'b1111111111000110;
    assign weights1[5][273] = 16'b1111111111011010;
    assign weights1[5][274] = 16'b1111111111100001;
    assign weights1[5][275] = 16'b1111111111011100;
    assign weights1[5][276] = 16'b1111111111011111;
    assign weights1[5][277] = 16'b1111111111110001;
    assign weights1[5][278] = 16'b1111111111110110;
    assign weights1[5][279] = 16'b1111111111111111;
    assign weights1[5][280] = 16'b0000000000011010;
    assign weights1[5][281] = 16'b0000000000100100;
    assign weights1[5][282] = 16'b0000000000011111;
    assign weights1[5][283] = 16'b0000000000000010;
    assign weights1[5][284] = 16'b1111111111111001;
    assign weights1[5][285] = 16'b1111111111110010;
    assign weights1[5][286] = 16'b1111111111110110;
    assign weights1[5][287] = 16'b1111111111110111;
    assign weights1[5][288] = 16'b1111111111111001;
    assign weights1[5][289] = 16'b1111111111111001;
    assign weights1[5][290] = 16'b0000000000101001;
    assign weights1[5][291] = 16'b0000000000101111;
    assign weights1[5][292] = 16'b0000000000101111;
    assign weights1[5][293] = 16'b0000000000110110;
    assign weights1[5][294] = 16'b0000000000100011;
    assign weights1[5][295] = 16'b0000000000000001;
    assign weights1[5][296] = 16'b1111111111101000;
    assign weights1[5][297] = 16'b1111111110111011;
    assign weights1[5][298] = 16'b1111111110010101;
    assign weights1[5][299] = 16'b1111111111000101;
    assign weights1[5][300] = 16'b1111111111000100;
    assign weights1[5][301] = 16'b1111111111011101;
    assign weights1[5][302] = 16'b1111111111100111;
    assign weights1[5][303] = 16'b1111111111011100;
    assign weights1[5][304] = 16'b1111111111100001;
    assign weights1[5][305] = 16'b1111111111110100;
    assign weights1[5][306] = 16'b1111111111111001;
    assign weights1[5][307] = 16'b1111111111110111;
    assign weights1[5][308] = 16'b0000000000011011;
    assign weights1[5][309] = 16'b0000000000010100;
    assign weights1[5][310] = 16'b0000000000001000;
    assign weights1[5][311] = 16'b0000000000001000;
    assign weights1[5][312] = 16'b1111111111111101;
    assign weights1[5][313] = 16'b0000000000000001;
    assign weights1[5][314] = 16'b1111111111100101;
    assign weights1[5][315] = 16'b1111111111110010;
    assign weights1[5][316] = 16'b1111111111100110;
    assign weights1[5][317] = 16'b1111111111101010;
    assign weights1[5][318] = 16'b0000000000000010;
    assign weights1[5][319] = 16'b0000000000100100;
    assign weights1[5][320] = 16'b0000000000011101;
    assign weights1[5][321] = 16'b0000000000111101;
    assign weights1[5][322] = 16'b0000000000110100;
    assign weights1[5][323] = 16'b1111111111111100;
    assign weights1[5][324] = 16'b1111111111011100;
    assign weights1[5][325] = 16'b1111111111001110;
    assign weights1[5][326] = 16'b1111111110101101;
    assign weights1[5][327] = 16'b1111111111000111;
    assign weights1[5][328] = 16'b1111111111010010;
    assign weights1[5][329] = 16'b1111111111001100;
    assign weights1[5][330] = 16'b1111111111100011;
    assign weights1[5][331] = 16'b1111111111101011;
    assign weights1[5][332] = 16'b1111111111101001;
    assign weights1[5][333] = 16'b1111111111111100;
    assign weights1[5][334] = 16'b1111111111101110;
    assign weights1[5][335] = 16'b1111111111110110;
    assign weights1[5][336] = 16'b0000000000011100;
    assign weights1[5][337] = 16'b0000000000010001;
    assign weights1[5][338] = 16'b1111111111111110;
    assign weights1[5][339] = 16'b1111111111111010;
    assign weights1[5][340] = 16'b1111111111110110;
    assign weights1[5][341] = 16'b1111111111110000;
    assign weights1[5][342] = 16'b1111111111101101;
    assign weights1[5][343] = 16'b1111111111011011;
    assign weights1[5][344] = 16'b1111111111100000;
    assign weights1[5][345] = 16'b1111111111110100;
    assign weights1[5][346] = 16'b1111111111111011;
    assign weights1[5][347] = 16'b0000000000010100;
    assign weights1[5][348] = 16'b0000000000100010;
    assign weights1[5][349] = 16'b0000000000101001;
    assign weights1[5][350] = 16'b0000000000010110;
    assign weights1[5][351] = 16'b0000000000000000;
    assign weights1[5][352] = 16'b1111111111001001;
    assign weights1[5][353] = 16'b1111111111011110;
    assign weights1[5][354] = 16'b1111111111100001;
    assign weights1[5][355] = 16'b1111111111110001;
    assign weights1[5][356] = 16'b1111111111110101;
    assign weights1[5][357] = 16'b1111111111100001;
    assign weights1[5][358] = 16'b1111111111100001;
    assign weights1[5][359] = 16'b1111111111100001;
    assign weights1[5][360] = 16'b1111111111101101;
    assign weights1[5][361] = 16'b1111111111110101;
    assign weights1[5][362] = 16'b1111111111101110;
    assign weights1[5][363] = 16'b1111111111110101;
    assign weights1[5][364] = 16'b0000000000001110;
    assign weights1[5][365] = 16'b0000000000000000;
    assign weights1[5][366] = 16'b0000000000000111;
    assign weights1[5][367] = 16'b1111111111111001;
    assign weights1[5][368] = 16'b1111111111110101;
    assign weights1[5][369] = 16'b1111111111101110;
    assign weights1[5][370] = 16'b1111111111111001;
    assign weights1[5][371] = 16'b1111111111011011;
    assign weights1[5][372] = 16'b1111111111101111;
    assign weights1[5][373] = 16'b1111111111110111;
    assign weights1[5][374] = 16'b0000000000000011;
    assign weights1[5][375] = 16'b0000000000101101;
    assign weights1[5][376] = 16'b0000000000100111;
    assign weights1[5][377] = 16'b0000000000010000;
    assign weights1[5][378] = 16'b0000000000010000;
    assign weights1[5][379] = 16'b1111111111110011;
    assign weights1[5][380] = 16'b1111111111011010;
    assign weights1[5][381] = 16'b1111111111111010;
    assign weights1[5][382] = 16'b1111111111010001;
    assign weights1[5][383] = 16'b1111111111101110;
    assign weights1[5][384] = 16'b1111111111010001;
    assign weights1[5][385] = 16'b1111111111101110;
    assign weights1[5][386] = 16'b1111111111100100;
    assign weights1[5][387] = 16'b1111111111111011;
    assign weights1[5][388] = 16'b1111111111101010;
    assign weights1[5][389] = 16'b1111111111101001;
    assign weights1[5][390] = 16'b1111111111101101;
    assign weights1[5][391] = 16'b1111111111111100;
    assign weights1[5][392] = 16'b0000000000001010;
    assign weights1[5][393] = 16'b1111111111111000;
    assign weights1[5][394] = 16'b1111111111110101;
    assign weights1[5][395] = 16'b1111111111110000;
    assign weights1[5][396] = 16'b1111111111101000;
    assign weights1[5][397] = 16'b1111111111101011;
    assign weights1[5][398] = 16'b1111111111100100;
    assign weights1[5][399] = 16'b1111111111011101;
    assign weights1[5][400] = 16'b1111111111101101;
    assign weights1[5][401] = 16'b0000000000000011;
    assign weights1[5][402] = 16'b1111111111111100;
    assign weights1[5][403] = 16'b0000000000001001;
    assign weights1[5][404] = 16'b0000000000011111;
    assign weights1[5][405] = 16'b0000000000001011;
    assign weights1[5][406] = 16'b0000000000000110;
    assign weights1[5][407] = 16'b1111111111110100;
    assign weights1[5][408] = 16'b1111111111101000;
    assign weights1[5][409] = 16'b1111111111100101;
    assign weights1[5][410] = 16'b1111111111011010;
    assign weights1[5][411] = 16'b1111111111111101;
    assign weights1[5][412] = 16'b1111111111100011;
    assign weights1[5][413] = 16'b1111111111110010;
    assign weights1[5][414] = 16'b1111111111100101;
    assign weights1[5][415] = 16'b1111111111111010;
    assign weights1[5][416] = 16'b1111111111111100;
    assign weights1[5][417] = 16'b1111111111110010;
    assign weights1[5][418] = 16'b1111111111101101;
    assign weights1[5][419] = 16'b1111111111110110;
    assign weights1[5][420] = 16'b0000000000001001;
    assign weights1[5][421] = 16'b1111111111110001;
    assign weights1[5][422] = 16'b0000000000000101;
    assign weights1[5][423] = 16'b1111111111110110;
    assign weights1[5][424] = 16'b1111111111110111;
    assign weights1[5][425] = 16'b1111111111100111;
    assign weights1[5][426] = 16'b1111111111110110;
    assign weights1[5][427] = 16'b1111111111111000;
    assign weights1[5][428] = 16'b1111111111111010;
    assign weights1[5][429] = 16'b1111111111111111;
    assign weights1[5][430] = 16'b1111111111111010;
    assign weights1[5][431] = 16'b0000000000001101;
    assign weights1[5][432] = 16'b1111111111111101;
    assign weights1[5][433] = 16'b0000000000011001;
    assign weights1[5][434] = 16'b1111111111110110;
    assign weights1[5][435] = 16'b1111111111100100;
    assign weights1[5][436] = 16'b1111111111011011;
    assign weights1[5][437] = 16'b1111111111101010;
    assign weights1[5][438] = 16'b1111111111011100;
    assign weights1[5][439] = 16'b1111111111110111;
    assign weights1[5][440] = 16'b1111111111110000;
    assign weights1[5][441] = 16'b1111111111111010;
    assign weights1[5][442] = 16'b1111111111110111;
    assign weights1[5][443] = 16'b1111111111100010;
    assign weights1[5][444] = 16'b0000000000010111;
    assign weights1[5][445] = 16'b0000000000001011;
    assign weights1[5][446] = 16'b0000000000000100;
    assign weights1[5][447] = 16'b1111111111101011;
    assign weights1[5][448] = 16'b0000000000001100;
    assign weights1[5][449] = 16'b1111111111111000;
    assign weights1[5][450] = 16'b1111111111111100;
    assign weights1[5][451] = 16'b1111111111101100;
    assign weights1[5][452] = 16'b1111111111101101;
    assign weights1[5][453] = 16'b1111111111111000;
    assign weights1[5][454] = 16'b1111111111110010;
    assign weights1[5][455] = 16'b1111111111111011;
    assign weights1[5][456] = 16'b0000000000010001;
    assign weights1[5][457] = 16'b1111111111111000;
    assign weights1[5][458] = 16'b1111111111111110;
    assign weights1[5][459] = 16'b0000000000000011;
    assign weights1[5][460] = 16'b0000000000000110;
    assign weights1[5][461] = 16'b0000000000000000;
    assign weights1[5][462] = 16'b0000000000001010;
    assign weights1[5][463] = 16'b1111111111100010;
    assign weights1[5][464] = 16'b1111111111110111;
    assign weights1[5][465] = 16'b1111111111011010;
    assign weights1[5][466] = 16'b1111111111100011;
    assign weights1[5][467] = 16'b0000000000001100;
    assign weights1[5][468] = 16'b1111111111111110;
    assign weights1[5][469] = 16'b0000000000010010;
    assign weights1[5][470] = 16'b0000000000010000;
    assign weights1[5][471] = 16'b1111111111111100;
    assign weights1[5][472] = 16'b0000000000001000;
    assign weights1[5][473] = 16'b0000000000001010;
    assign weights1[5][474] = 16'b1111111111111111;
    assign weights1[5][475] = 16'b1111111111111101;
    assign weights1[5][476] = 16'b0000000000001100;
    assign weights1[5][477] = 16'b0000000000000001;
    assign weights1[5][478] = 16'b0000000000000110;
    assign weights1[5][479] = 16'b0000000000001010;
    assign weights1[5][480] = 16'b0000000000001010;
    assign weights1[5][481] = 16'b1111111111110011;
    assign weights1[5][482] = 16'b1111111111101111;
    assign weights1[5][483] = 16'b0000000000001010;
    assign weights1[5][484] = 16'b1111111111110100;
    assign weights1[5][485] = 16'b0000000000000010;
    assign weights1[5][486] = 16'b1111111111110001;
    assign weights1[5][487] = 16'b1111111111101010;
    assign weights1[5][488] = 16'b1111111111110001;
    assign weights1[5][489] = 16'b1111111111110101;
    assign weights1[5][490] = 16'b0000000000000001;
    assign weights1[5][491] = 16'b1111111111101101;
    assign weights1[5][492] = 16'b1111111111111010;
    assign weights1[5][493] = 16'b0000000000000110;
    assign weights1[5][494] = 16'b1111111111111001;
    assign weights1[5][495] = 16'b0000000000001101;
    assign weights1[5][496] = 16'b1111111111101000;
    assign weights1[5][497] = 16'b0000000000010110;
    assign weights1[5][498] = 16'b0000000000011110;
    assign weights1[5][499] = 16'b0000000000010100;
    assign weights1[5][500] = 16'b1111111111101110;
    assign weights1[5][501] = 16'b0000000000000010;
    assign weights1[5][502] = 16'b1111111111110010;
    assign weights1[5][503] = 16'b1111111111110011;
    assign weights1[5][504] = 16'b0000000000001011;
    assign weights1[5][505] = 16'b0000000000001001;
    assign weights1[5][506] = 16'b0000000000001111;
    assign weights1[5][507] = 16'b0000000000000010;
    assign weights1[5][508] = 16'b1111111111111100;
    assign weights1[5][509] = 16'b0000000000010001;
    assign weights1[5][510] = 16'b0000000000001100;
    assign weights1[5][511] = 16'b1111111111110010;
    assign weights1[5][512] = 16'b1111111111111110;
    assign weights1[5][513] = 16'b0000000000000110;
    assign weights1[5][514] = 16'b1111111111111011;
    assign weights1[5][515] = 16'b1111111111110110;
    assign weights1[5][516] = 16'b1111111111110000;
    assign weights1[5][517] = 16'b0000000000000101;
    assign weights1[5][518] = 16'b0000000000010101;
    assign weights1[5][519] = 16'b0000000000001011;
    assign weights1[5][520] = 16'b1111111111110000;
    assign weights1[5][521] = 16'b1111111111110100;
    assign weights1[5][522] = 16'b1111111111111010;
    assign weights1[5][523] = 16'b1111111111110101;
    assign weights1[5][524] = 16'b0000000000000001;
    assign weights1[5][525] = 16'b0000000000001111;
    assign weights1[5][526] = 16'b0000000000100111;
    assign weights1[5][527] = 16'b0000000000100011;
    assign weights1[5][528] = 16'b0000000000000011;
    assign weights1[5][529] = 16'b1111111111101101;
    assign weights1[5][530] = 16'b1111111111110100;
    assign weights1[5][531] = 16'b1111111111111010;
    assign weights1[5][532] = 16'b0000000000001011;
    assign weights1[5][533] = 16'b0000000000010001;
    assign weights1[5][534] = 16'b0000000000100010;
    assign weights1[5][535] = 16'b0000000000001000;
    assign weights1[5][536] = 16'b0000000000001101;
    assign weights1[5][537] = 16'b0000000000000100;
    assign weights1[5][538] = 16'b1111111111111000;
    assign weights1[5][539] = 16'b1111111111101010;
    assign weights1[5][540] = 16'b1111111111111000;
    assign weights1[5][541] = 16'b1111111111100101;
    assign weights1[5][542] = 16'b0000000000000100;
    assign weights1[5][543] = 16'b1111111111101000;
    assign weights1[5][544] = 16'b1111111111101010;
    assign weights1[5][545] = 16'b1111111111111110;
    assign weights1[5][546] = 16'b1111111111101101;
    assign weights1[5][547] = 16'b0000000000001101;
    assign weights1[5][548] = 16'b1111111111110011;
    assign weights1[5][549] = 16'b1111111111101110;
    assign weights1[5][550] = 16'b0000000000000011;
    assign weights1[5][551] = 16'b0000000000000001;
    assign weights1[5][552] = 16'b1111111111101110;
    assign weights1[5][553] = 16'b1111111111110101;
    assign weights1[5][554] = 16'b0000000000000010;
    assign weights1[5][555] = 16'b0000000000000011;
    assign weights1[5][556] = 16'b1111111111111001;
    assign weights1[5][557] = 16'b1111111111111000;
    assign weights1[5][558] = 16'b1111111111110100;
    assign weights1[5][559] = 16'b1111111111110101;
    assign weights1[5][560] = 16'b0000000000010010;
    assign weights1[5][561] = 16'b0000000000010110;
    assign weights1[5][562] = 16'b0000000000010011;
    assign weights1[5][563] = 16'b0000000000001011;
    assign weights1[5][564] = 16'b0000000000000110;
    assign weights1[5][565] = 16'b0000000000000110;
    assign weights1[5][566] = 16'b1111111111110010;
    assign weights1[5][567] = 16'b0000000000000101;
    assign weights1[5][568] = 16'b0000000000000001;
    assign weights1[5][569] = 16'b0000000000000001;
    assign weights1[5][570] = 16'b0000000000000001;
    assign weights1[5][571] = 16'b1111111111110100;
    assign weights1[5][572] = 16'b1111111111110100;
    assign weights1[5][573] = 16'b1111111111111010;
    assign weights1[5][574] = 16'b0000000000001001;
    assign weights1[5][575] = 16'b0000000000000100;
    assign weights1[5][576] = 16'b1111111111111010;
    assign weights1[5][577] = 16'b0000000000001011;
    assign weights1[5][578] = 16'b1111111111100011;
    assign weights1[5][579] = 16'b1111111111101011;
    assign weights1[5][580] = 16'b1111111111111100;
    assign weights1[5][581] = 16'b1111111111111001;
    assign weights1[5][582] = 16'b0000000000001101;
    assign weights1[5][583] = 16'b1111111111111110;
    assign weights1[5][584] = 16'b1111111111110101;
    assign weights1[5][585] = 16'b0000000000000110;
    assign weights1[5][586] = 16'b1111111111110100;
    assign weights1[5][587] = 16'b1111111111111000;
    assign weights1[5][588] = 16'b0000000000010100;
    assign weights1[5][589] = 16'b0000000000010000;
    assign weights1[5][590] = 16'b0000000000001001;
    assign weights1[5][591] = 16'b1111111111111111;
    assign weights1[5][592] = 16'b1111111111101010;
    assign weights1[5][593] = 16'b1111111111101001;
    assign weights1[5][594] = 16'b1111111111110110;
    assign weights1[5][595] = 16'b0000000000000100;
    assign weights1[5][596] = 16'b1111111111110101;
    assign weights1[5][597] = 16'b0000000000000000;
    assign weights1[5][598] = 16'b0000000000000100;
    assign weights1[5][599] = 16'b1111111111110100;
    assign weights1[5][600] = 16'b1111111111101111;
    assign weights1[5][601] = 16'b1111111111100000;
    assign weights1[5][602] = 16'b0000000000000010;
    assign weights1[5][603] = 16'b0000000000010000;
    assign weights1[5][604] = 16'b1111111111110010;
    assign weights1[5][605] = 16'b1111111111111110;
    assign weights1[5][606] = 16'b0000000000000100;
    assign weights1[5][607] = 16'b1111111111110011;
    assign weights1[5][608] = 16'b1111111111101010;
    assign weights1[5][609] = 16'b1111111111011110;
    assign weights1[5][610] = 16'b1111111111101111;
    assign weights1[5][611] = 16'b1111111111100110;
    assign weights1[5][612] = 16'b1111111111110110;
    assign weights1[5][613] = 16'b1111111111111001;
    assign weights1[5][614] = 16'b1111111111111000;
    assign weights1[5][615] = 16'b1111111111111000;
    assign weights1[5][616] = 16'b0000000000001100;
    assign weights1[5][617] = 16'b0000000000011001;
    assign weights1[5][618] = 16'b0000000000000101;
    assign weights1[5][619] = 16'b0000000000001011;
    assign weights1[5][620] = 16'b1111111111111111;
    assign weights1[5][621] = 16'b1111111111110011;
    assign weights1[5][622] = 16'b1111111111110100;
    assign weights1[5][623] = 16'b1111111111110110;
    assign weights1[5][624] = 16'b1111111111111000;
    assign weights1[5][625] = 16'b0000000000000101;
    assign weights1[5][626] = 16'b1111111111110100;
    assign weights1[5][627] = 16'b0000000000001010;
    assign weights1[5][628] = 16'b0000000000000110;
    assign weights1[5][629] = 16'b1111111111110111;
    assign weights1[5][630] = 16'b1111111111101101;
    assign weights1[5][631] = 16'b1111111111110010;
    assign weights1[5][632] = 16'b1111111111101010;
    assign weights1[5][633] = 16'b1111111111110010;
    assign weights1[5][634] = 16'b0000000000001011;
    assign weights1[5][635] = 16'b1111111111111000;
    assign weights1[5][636] = 16'b0000000000011110;
    assign weights1[5][637] = 16'b1111111111111010;
    assign weights1[5][638] = 16'b1111111111011100;
    assign weights1[5][639] = 16'b1111111111111010;
    assign weights1[5][640] = 16'b0000000000000000;
    assign weights1[5][641] = 16'b1111111111111001;
    assign weights1[5][642] = 16'b1111111111110111;
    assign weights1[5][643] = 16'b1111111111111010;
    assign weights1[5][644] = 16'b0000000000000101;
    assign weights1[5][645] = 16'b0000000000001011;
    assign weights1[5][646] = 16'b0000000000001111;
    assign weights1[5][647] = 16'b0000000000001001;
    assign weights1[5][648] = 16'b0000000000001000;
    assign weights1[5][649] = 16'b0000000000000110;
    assign weights1[5][650] = 16'b0000000000001010;
    assign weights1[5][651] = 16'b1111111111110001;
    assign weights1[5][652] = 16'b1111111111111011;
    assign weights1[5][653] = 16'b0000000000000110;
    assign weights1[5][654] = 16'b0000000000010000;
    assign weights1[5][655] = 16'b0000000000000100;
    assign weights1[5][656] = 16'b1111111111111001;
    assign weights1[5][657] = 16'b1111111111111010;
    assign weights1[5][658] = 16'b1111111111111100;
    assign weights1[5][659] = 16'b0000000000011100;
    assign weights1[5][660] = 16'b1111111111110100;
    assign weights1[5][661] = 16'b0000000000001001;
    assign weights1[5][662] = 16'b1111111111101000;
    assign weights1[5][663] = 16'b1111111111111011;
    assign weights1[5][664] = 16'b1111111111110111;
    assign weights1[5][665] = 16'b1111111111110011;
    assign weights1[5][666] = 16'b1111111111111001;
    assign weights1[5][667] = 16'b1111111111101100;
    assign weights1[5][668] = 16'b1111111111111111;
    assign weights1[5][669] = 16'b1111111111111011;
    assign weights1[5][670] = 16'b0000000000000010;
    assign weights1[5][671] = 16'b0000000000000000;
    assign weights1[5][672] = 16'b0000000000000100;
    assign weights1[5][673] = 16'b0000000000001011;
    assign weights1[5][674] = 16'b0000000000000100;
    assign weights1[5][675] = 16'b0000000000000100;
    assign weights1[5][676] = 16'b1111111111111110;
    assign weights1[5][677] = 16'b0000000000000010;
    assign weights1[5][678] = 16'b1111111111111011;
    assign weights1[5][679] = 16'b0000000000000110;
    assign weights1[5][680] = 16'b0000000000011001;
    assign weights1[5][681] = 16'b0000000000000010;
    assign weights1[5][682] = 16'b1111111111111110;
    assign weights1[5][683] = 16'b1111111111110101;
    assign weights1[5][684] = 16'b1111111111100011;
    assign weights1[5][685] = 16'b0000000000000010;
    assign weights1[5][686] = 16'b1111111111101011;
    assign weights1[5][687] = 16'b1111111111110010;
    assign weights1[5][688] = 16'b1111111111101000;
    assign weights1[5][689] = 16'b1111111111111101;
    assign weights1[5][690] = 16'b1111111111100010;
    assign weights1[5][691] = 16'b1111111111111001;
    assign weights1[5][692] = 16'b1111111111101111;
    assign weights1[5][693] = 16'b1111111111111101;
    assign weights1[5][694] = 16'b1111111111110001;
    assign weights1[5][695] = 16'b1111111111111110;
    assign weights1[5][696] = 16'b1111111111111101;
    assign weights1[5][697] = 16'b1111111111111100;
    assign weights1[5][698] = 16'b0000000000000100;
    assign weights1[5][699] = 16'b0000000000000100;
    assign weights1[5][700] = 16'b1111111111111101;
    assign weights1[5][701] = 16'b0000000000001110;
    assign weights1[5][702] = 16'b0000000000010000;
    assign weights1[5][703] = 16'b0000000000001010;
    assign weights1[5][704] = 16'b0000000000001000;
    assign weights1[5][705] = 16'b0000000000001100;
    assign weights1[5][706] = 16'b0000000000000010;
    assign weights1[5][707] = 16'b0000000000000110;
    assign weights1[5][708] = 16'b1111111111111111;
    assign weights1[5][709] = 16'b1111111111100101;
    assign weights1[5][710] = 16'b1111111111111111;
    assign weights1[5][711] = 16'b1111111111101000;
    assign weights1[5][712] = 16'b1111111111110111;
    assign weights1[5][713] = 16'b1111111111110101;
    assign weights1[5][714] = 16'b1111111111111110;
    assign weights1[5][715] = 16'b1111111111110101;
    assign weights1[5][716] = 16'b0000000000001111;
    assign weights1[5][717] = 16'b0000000000010101;
    assign weights1[5][718] = 16'b0000000000001010;
    assign weights1[5][719] = 16'b1111111111111110;
    assign weights1[5][720] = 16'b1111111111101111;
    assign weights1[5][721] = 16'b1111111111111111;
    assign weights1[5][722] = 16'b1111111111111000;
    assign weights1[5][723] = 16'b1111111111111010;
    assign weights1[5][724] = 16'b1111111111111111;
    assign weights1[5][725] = 16'b0000000000000001;
    assign weights1[5][726] = 16'b1111111111111101;
    assign weights1[5][727] = 16'b0000000000000001;
    assign weights1[5][728] = 16'b0000000000000001;
    assign weights1[5][729] = 16'b0000000000000110;
    assign weights1[5][730] = 16'b0000000000010010;
    assign weights1[5][731] = 16'b0000000000010001;
    assign weights1[5][732] = 16'b0000000000000100;
    assign weights1[5][733] = 16'b0000000000000011;
    assign weights1[5][734] = 16'b0000000000010110;
    assign weights1[5][735] = 16'b0000000000001001;
    assign weights1[5][736] = 16'b0000000000000011;
    assign weights1[5][737] = 16'b1111111111111101;
    assign weights1[5][738] = 16'b0000000000011100;
    assign weights1[5][739] = 16'b1111111111110100;
    assign weights1[5][740] = 16'b0000000000001100;
    assign weights1[5][741] = 16'b0000000000001101;
    assign weights1[5][742] = 16'b1111111111110001;
    assign weights1[5][743] = 16'b1111111111110001;
    assign weights1[5][744] = 16'b0000000000000111;
    assign weights1[5][745] = 16'b0000000000011000;
    assign weights1[5][746] = 16'b0000000000010011;
    assign weights1[5][747] = 16'b0000000000010011;
    assign weights1[5][748] = 16'b0000000000000110;
    assign weights1[5][749] = 16'b0000000000010011;
    assign weights1[5][750] = 16'b1111111111111011;
    assign weights1[5][751] = 16'b1111111111111010;
    assign weights1[5][752] = 16'b0000000000000000;
    assign weights1[5][753] = 16'b0000000000000000;
    assign weights1[5][754] = 16'b1111111111111110;
    assign weights1[5][755] = 16'b1111111111111111;
    assign weights1[5][756] = 16'b0000000000000101;
    assign weights1[5][757] = 16'b0000000000000110;
    assign weights1[5][758] = 16'b0000000000001100;
    assign weights1[5][759] = 16'b0000000000010001;
    assign weights1[5][760] = 16'b0000000000010001;
    assign weights1[5][761] = 16'b0000000000010011;
    assign weights1[5][762] = 16'b0000000000001111;
    assign weights1[5][763] = 16'b0000000000000110;
    assign weights1[5][764] = 16'b0000000000001011;
    assign weights1[5][765] = 16'b0000000000000100;
    assign weights1[5][766] = 16'b0000000000001101;
    assign weights1[5][767] = 16'b1111111111111111;
    assign weights1[5][768] = 16'b0000000000001001;
    assign weights1[5][769] = 16'b0000000000001111;
    assign weights1[5][770] = 16'b1111111111111100;
    assign weights1[5][771] = 16'b0000000000010000;
    assign weights1[5][772] = 16'b0000000000001111;
    assign weights1[5][773] = 16'b0000000000010011;
    assign weights1[5][774] = 16'b0000000000010010;
    assign weights1[5][775] = 16'b0000000000000010;
    assign weights1[5][776] = 16'b0000000000000110;
    assign weights1[5][777] = 16'b0000000000000011;
    assign weights1[5][778] = 16'b1111111111111101;
    assign weights1[5][779] = 16'b1111111111111011;
    assign weights1[5][780] = 16'b0000000000000000;
    assign weights1[5][781] = 16'b0000000000000001;
    assign weights1[5][782] = 16'b1111111111111111;
    assign weights1[5][783] = 16'b1111111111111111;
    assign weights1[6][0] = 16'b0000000000000000;
    assign weights1[6][1] = 16'b0000000000000000;
    assign weights1[6][2] = 16'b0000000000000000;
    assign weights1[6][3] = 16'b0000000000000000;
    assign weights1[6][4] = 16'b0000000000000000;
    assign weights1[6][5] = 16'b0000000000000000;
    assign weights1[6][6] = 16'b0000000000000000;
    assign weights1[6][7] = 16'b0000000000000000;
    assign weights1[6][8] = 16'b0000000000000000;
    assign weights1[6][9] = 16'b0000000000000000;
    assign weights1[6][10] = 16'b0000000000000000;
    assign weights1[6][11] = 16'b0000000000000000;
    assign weights1[6][12] = 16'b0000000000000000;
    assign weights1[6][13] = 16'b0000000000000000;
    assign weights1[6][14] = 16'b0000000000000000;
    assign weights1[6][15] = 16'b0000000000000000;
    assign weights1[6][16] = 16'b0000000000000000;
    assign weights1[6][17] = 16'b0000000000000000;
    assign weights1[6][18] = 16'b0000000000000000;
    assign weights1[6][19] = 16'b0000000000000000;
    assign weights1[6][20] = 16'b0000000000000000;
    assign weights1[6][21] = 16'b0000000000000000;
    assign weights1[6][22] = 16'b0000000000000000;
    assign weights1[6][23] = 16'b0000000000000000;
    assign weights1[6][24] = 16'b0000000000000000;
    assign weights1[6][25] = 16'b0000000000000000;
    assign weights1[6][26] = 16'b0000000000000000;
    assign weights1[6][27] = 16'b0000000000000000;
    assign weights1[6][28] = 16'b0000000000000000;
    assign weights1[6][29] = 16'b0000000000000000;
    assign weights1[6][30] = 16'b0000000000000000;
    assign weights1[6][31] = 16'b0000000000000000;
    assign weights1[6][32] = 16'b0000000000000000;
    assign weights1[6][33] = 16'b0000000000000000;
    assign weights1[6][34] = 16'b0000000000000000;
    assign weights1[6][35] = 16'b0000000000000000;
    assign weights1[6][36] = 16'b0000000000000000;
    assign weights1[6][37] = 16'b0000000000000000;
    assign weights1[6][38] = 16'b0000000000000000;
    assign weights1[6][39] = 16'b0000000000000000;
    assign weights1[6][40] = 16'b0000000000000000;
    assign weights1[6][41] = 16'b0000000000000000;
    assign weights1[6][42] = 16'b0000000000000000;
    assign weights1[6][43] = 16'b0000000000000000;
    assign weights1[6][44] = 16'b0000000000000000;
    assign weights1[6][45] = 16'b0000000000000000;
    assign weights1[6][46] = 16'b0000000000000000;
    assign weights1[6][47] = 16'b0000000000000000;
    assign weights1[6][48] = 16'b0000000000000000;
    assign weights1[6][49] = 16'b0000000000000000;
    assign weights1[6][50] = 16'b0000000000000000;
    assign weights1[6][51] = 16'b0000000000000000;
    assign weights1[6][52] = 16'b0000000000000000;
    assign weights1[6][53] = 16'b0000000000000000;
    assign weights1[6][54] = 16'b0000000000000000;
    assign weights1[6][55] = 16'b0000000000000000;
    assign weights1[6][56] = 16'b0000000000000000;
    assign weights1[6][57] = 16'b0000000000000000;
    assign weights1[6][58] = 16'b0000000000000000;
    assign weights1[6][59] = 16'b0000000000000000;
    assign weights1[6][60] = 16'b0000000000000000;
    assign weights1[6][61] = 16'b0000000000000000;
    assign weights1[6][62] = 16'b0000000000000000;
    assign weights1[6][63] = 16'b0000000000000000;
    assign weights1[6][64] = 16'b0000000000000000;
    assign weights1[6][65] = 16'b0000000000000000;
    assign weights1[6][66] = 16'b0000000000000000;
    assign weights1[6][67] = 16'b0000000000000000;
    assign weights1[6][68] = 16'b0000000000000000;
    assign weights1[6][69] = 16'b0000000000000000;
    assign weights1[6][70] = 16'b0000000000000000;
    assign weights1[6][71] = 16'b0000000000000000;
    assign weights1[6][72] = 16'b0000000000000000;
    assign weights1[6][73] = 16'b0000000000000000;
    assign weights1[6][74] = 16'b0000000000000000;
    assign weights1[6][75] = 16'b0000000000000000;
    assign weights1[6][76] = 16'b0000000000000000;
    assign weights1[6][77] = 16'b0000000000000000;
    assign weights1[6][78] = 16'b0000000000000000;
    assign weights1[6][79] = 16'b0000000000000000;
    assign weights1[6][80] = 16'b0000000000000000;
    assign weights1[6][81] = 16'b0000000000000000;
    assign weights1[6][82] = 16'b0000000000000000;
    assign weights1[6][83] = 16'b0000000000000000;
    assign weights1[6][84] = 16'b0000000000000000;
    assign weights1[6][85] = 16'b0000000000000000;
    assign weights1[6][86] = 16'b0000000000000000;
    assign weights1[6][87] = 16'b0000000000000000;
    assign weights1[6][88] = 16'b0000000000000000;
    assign weights1[6][89] = 16'b0000000000000000;
    assign weights1[6][90] = 16'b0000000000000000;
    assign weights1[6][91] = 16'b0000000000000000;
    assign weights1[6][92] = 16'b0000000000000000;
    assign weights1[6][93] = 16'b0000000000000000;
    assign weights1[6][94] = 16'b0000000000000000;
    assign weights1[6][95] = 16'b0000000000000000;
    assign weights1[6][96] = 16'b0000000000000000;
    assign weights1[6][97] = 16'b0000000000000000;
    assign weights1[6][98] = 16'b0000000000000000;
    assign weights1[6][99] = 16'b0000000000000000;
    assign weights1[6][100] = 16'b0000000000000000;
    assign weights1[6][101] = 16'b0000000000000000;
    assign weights1[6][102] = 16'b0000000000000000;
    assign weights1[6][103] = 16'b0000000000000000;
    assign weights1[6][104] = 16'b0000000000000000;
    assign weights1[6][105] = 16'b0000000000000000;
    assign weights1[6][106] = 16'b0000000000000000;
    assign weights1[6][107] = 16'b0000000000000000;
    assign weights1[6][108] = 16'b0000000000000000;
    assign weights1[6][109] = 16'b0000000000000000;
    assign weights1[6][110] = 16'b0000000000000000;
    assign weights1[6][111] = 16'b0000000000000000;
    assign weights1[6][112] = 16'b0000000000000000;
    assign weights1[6][113] = 16'b0000000000000000;
    assign weights1[6][114] = 16'b0000000000000000;
    assign weights1[6][115] = 16'b0000000000000000;
    assign weights1[6][116] = 16'b0000000000000000;
    assign weights1[6][117] = 16'b0000000000000000;
    assign weights1[6][118] = 16'b0000000000000000;
    assign weights1[6][119] = 16'b0000000000000000;
    assign weights1[6][120] = 16'b0000000000000000;
    assign weights1[6][121] = 16'b0000000000000000;
    assign weights1[6][122] = 16'b0000000000000000;
    assign weights1[6][123] = 16'b0000000000000000;
    assign weights1[6][124] = 16'b0000000000000000;
    assign weights1[6][125] = 16'b0000000000000000;
    assign weights1[6][126] = 16'b0000000000000000;
    assign weights1[6][127] = 16'b0000000000000000;
    assign weights1[6][128] = 16'b0000000000000000;
    assign weights1[6][129] = 16'b0000000000000000;
    assign weights1[6][130] = 16'b0000000000000000;
    assign weights1[6][131] = 16'b0000000000000000;
    assign weights1[6][132] = 16'b0000000000000000;
    assign weights1[6][133] = 16'b0000000000000000;
    assign weights1[6][134] = 16'b0000000000000000;
    assign weights1[6][135] = 16'b0000000000000000;
    assign weights1[6][136] = 16'b0000000000000000;
    assign weights1[6][137] = 16'b0000000000000000;
    assign weights1[6][138] = 16'b0000000000000000;
    assign weights1[6][139] = 16'b0000000000000000;
    assign weights1[6][140] = 16'b0000000000000000;
    assign weights1[6][141] = 16'b0000000000000000;
    assign weights1[6][142] = 16'b0000000000000000;
    assign weights1[6][143] = 16'b0000000000000000;
    assign weights1[6][144] = 16'b0000000000000000;
    assign weights1[6][145] = 16'b0000000000000000;
    assign weights1[6][146] = 16'b0000000000000000;
    assign weights1[6][147] = 16'b0000000000000000;
    assign weights1[6][148] = 16'b0000000000000000;
    assign weights1[6][149] = 16'b0000000000000000;
    assign weights1[6][150] = 16'b0000000000000000;
    assign weights1[6][151] = 16'b0000000000000000;
    assign weights1[6][152] = 16'b0000000000000000;
    assign weights1[6][153] = 16'b0000000000000000;
    assign weights1[6][154] = 16'b0000000000000000;
    assign weights1[6][155] = 16'b0000000000000000;
    assign weights1[6][156] = 16'b0000000000000000;
    assign weights1[6][157] = 16'b0000000000000000;
    assign weights1[6][158] = 16'b0000000000000000;
    assign weights1[6][159] = 16'b0000000000000000;
    assign weights1[6][160] = 16'b0000000000000000;
    assign weights1[6][161] = 16'b0000000000000000;
    assign weights1[6][162] = 16'b0000000000000000;
    assign weights1[6][163] = 16'b0000000000000000;
    assign weights1[6][164] = 16'b0000000000000000;
    assign weights1[6][165] = 16'b0000000000000000;
    assign weights1[6][166] = 16'b0000000000000000;
    assign weights1[6][167] = 16'b0000000000000000;
    assign weights1[6][168] = 16'b0000000000000000;
    assign weights1[6][169] = 16'b0000000000000000;
    assign weights1[6][170] = 16'b0000000000000000;
    assign weights1[6][171] = 16'b0000000000000000;
    assign weights1[6][172] = 16'b0000000000000000;
    assign weights1[6][173] = 16'b0000000000000000;
    assign weights1[6][174] = 16'b0000000000000000;
    assign weights1[6][175] = 16'b0000000000000000;
    assign weights1[6][176] = 16'b0000000000000000;
    assign weights1[6][177] = 16'b0000000000000000;
    assign weights1[6][178] = 16'b0000000000000000;
    assign weights1[6][179] = 16'b0000000000000000;
    assign weights1[6][180] = 16'b0000000000000000;
    assign weights1[6][181] = 16'b0000000000000000;
    assign weights1[6][182] = 16'b0000000000000000;
    assign weights1[6][183] = 16'b0000000000000000;
    assign weights1[6][184] = 16'b0000000000000000;
    assign weights1[6][185] = 16'b0000000000000000;
    assign weights1[6][186] = 16'b0000000000000000;
    assign weights1[6][187] = 16'b0000000000000000;
    assign weights1[6][188] = 16'b0000000000000000;
    assign weights1[6][189] = 16'b0000000000000000;
    assign weights1[6][190] = 16'b0000000000000000;
    assign weights1[6][191] = 16'b0000000000000000;
    assign weights1[6][192] = 16'b0000000000000000;
    assign weights1[6][193] = 16'b0000000000000000;
    assign weights1[6][194] = 16'b0000000000000000;
    assign weights1[6][195] = 16'b0000000000000000;
    assign weights1[6][196] = 16'b0000000000000000;
    assign weights1[6][197] = 16'b0000000000000000;
    assign weights1[6][198] = 16'b0000000000000000;
    assign weights1[6][199] = 16'b0000000000000000;
    assign weights1[6][200] = 16'b0000000000000000;
    assign weights1[6][201] = 16'b0000000000000000;
    assign weights1[6][202] = 16'b0000000000000000;
    assign weights1[6][203] = 16'b0000000000000000;
    assign weights1[6][204] = 16'b0000000000000000;
    assign weights1[6][205] = 16'b0000000000000000;
    assign weights1[6][206] = 16'b0000000000000000;
    assign weights1[6][207] = 16'b0000000000000000;
    assign weights1[6][208] = 16'b0000000000000000;
    assign weights1[6][209] = 16'b0000000000000000;
    assign weights1[6][210] = 16'b0000000000000000;
    assign weights1[6][211] = 16'b0000000000000000;
    assign weights1[6][212] = 16'b0000000000000000;
    assign weights1[6][213] = 16'b0000000000000000;
    assign weights1[6][214] = 16'b0000000000000000;
    assign weights1[6][215] = 16'b0000000000000000;
    assign weights1[6][216] = 16'b0000000000000000;
    assign weights1[6][217] = 16'b0000000000000000;
    assign weights1[6][218] = 16'b0000000000000000;
    assign weights1[6][219] = 16'b0000000000000000;
    assign weights1[6][220] = 16'b0000000000000000;
    assign weights1[6][221] = 16'b0000000000000000;
    assign weights1[6][222] = 16'b0000000000000000;
    assign weights1[6][223] = 16'b0000000000000000;
    assign weights1[6][224] = 16'b0000000000000000;
    assign weights1[6][225] = 16'b0000000000000000;
    assign weights1[6][226] = 16'b0000000000000000;
    assign weights1[6][227] = 16'b0000000000000000;
    assign weights1[6][228] = 16'b0000000000000000;
    assign weights1[6][229] = 16'b0000000000000000;
    assign weights1[6][230] = 16'b0000000000000000;
    assign weights1[6][231] = 16'b0000000000000000;
    assign weights1[6][232] = 16'b0000000000000000;
    assign weights1[6][233] = 16'b0000000000000000;
    assign weights1[6][234] = 16'b0000000000000000;
    assign weights1[6][235] = 16'b0000000000000000;
    assign weights1[6][236] = 16'b0000000000000000;
    assign weights1[6][237] = 16'b0000000000000000;
    assign weights1[6][238] = 16'b0000000000000000;
    assign weights1[6][239] = 16'b0000000000000000;
    assign weights1[6][240] = 16'b0000000000000000;
    assign weights1[6][241] = 16'b0000000000000000;
    assign weights1[6][242] = 16'b0000000000000000;
    assign weights1[6][243] = 16'b0000000000000000;
    assign weights1[6][244] = 16'b0000000000000000;
    assign weights1[6][245] = 16'b0000000000000000;
    assign weights1[6][246] = 16'b0000000000000000;
    assign weights1[6][247] = 16'b0000000000000000;
    assign weights1[6][248] = 16'b0000000000000000;
    assign weights1[6][249] = 16'b0000000000000000;
    assign weights1[6][250] = 16'b0000000000000000;
    assign weights1[6][251] = 16'b0000000000000000;
    assign weights1[6][252] = 16'b0000000000000000;
    assign weights1[6][253] = 16'b0000000000000000;
    assign weights1[6][254] = 16'b0000000000000000;
    assign weights1[6][255] = 16'b0000000000000000;
    assign weights1[6][256] = 16'b0000000000000000;
    assign weights1[6][257] = 16'b0000000000000000;
    assign weights1[6][258] = 16'b0000000000000000;
    assign weights1[6][259] = 16'b0000000000000000;
    assign weights1[6][260] = 16'b0000000000000000;
    assign weights1[6][261] = 16'b0000000000000000;
    assign weights1[6][262] = 16'b0000000000000000;
    assign weights1[6][263] = 16'b0000000000000000;
    assign weights1[6][264] = 16'b0000000000000000;
    assign weights1[6][265] = 16'b0000000000000000;
    assign weights1[6][266] = 16'b0000000000000000;
    assign weights1[6][267] = 16'b0000000000000000;
    assign weights1[6][268] = 16'b0000000000000000;
    assign weights1[6][269] = 16'b0000000000000000;
    assign weights1[6][270] = 16'b0000000000000000;
    assign weights1[6][271] = 16'b0000000000000000;
    assign weights1[6][272] = 16'b0000000000000000;
    assign weights1[6][273] = 16'b0000000000000000;
    assign weights1[6][274] = 16'b0000000000000000;
    assign weights1[6][275] = 16'b0000000000000000;
    assign weights1[6][276] = 16'b0000000000000000;
    assign weights1[6][277] = 16'b0000000000000000;
    assign weights1[6][278] = 16'b0000000000000000;
    assign weights1[6][279] = 16'b0000000000000000;
    assign weights1[6][280] = 16'b0000000000000000;
    assign weights1[6][281] = 16'b0000000000000000;
    assign weights1[6][282] = 16'b0000000000000000;
    assign weights1[6][283] = 16'b0000000000000000;
    assign weights1[6][284] = 16'b0000000000000000;
    assign weights1[6][285] = 16'b0000000000000000;
    assign weights1[6][286] = 16'b0000000000000000;
    assign weights1[6][287] = 16'b0000000000000000;
    assign weights1[6][288] = 16'b0000000000000000;
    assign weights1[6][289] = 16'b0000000000000000;
    assign weights1[6][290] = 16'b0000000000000000;
    assign weights1[6][291] = 16'b0000000000000000;
    assign weights1[6][292] = 16'b0000000000000000;
    assign weights1[6][293] = 16'b0000000000000000;
    assign weights1[6][294] = 16'b0000000000000000;
    assign weights1[6][295] = 16'b0000000000000000;
    assign weights1[6][296] = 16'b0000000000000000;
    assign weights1[6][297] = 16'b0000000000000000;
    assign weights1[6][298] = 16'b0000000000000000;
    assign weights1[6][299] = 16'b0000000000000000;
    assign weights1[6][300] = 16'b0000000000000000;
    assign weights1[6][301] = 16'b0000000000000000;
    assign weights1[6][302] = 16'b0000000000000000;
    assign weights1[6][303] = 16'b0000000000000000;
    assign weights1[6][304] = 16'b0000000000000000;
    assign weights1[6][305] = 16'b0000000000000000;
    assign weights1[6][306] = 16'b0000000000000000;
    assign weights1[6][307] = 16'b0000000000000000;
    assign weights1[6][308] = 16'b0000000000000000;
    assign weights1[6][309] = 16'b0000000000000000;
    assign weights1[6][310] = 16'b0000000000000000;
    assign weights1[6][311] = 16'b0000000000000000;
    assign weights1[6][312] = 16'b0000000000000000;
    assign weights1[6][313] = 16'b0000000000000000;
    assign weights1[6][314] = 16'b0000000000000000;
    assign weights1[6][315] = 16'b0000000000000000;
    assign weights1[6][316] = 16'b0000000000000000;
    assign weights1[6][317] = 16'b0000000000000000;
    assign weights1[6][318] = 16'b0000000000000000;
    assign weights1[6][319] = 16'b0000000000000000;
    assign weights1[6][320] = 16'b0000000000000000;
    assign weights1[6][321] = 16'b0000000000000000;
    assign weights1[6][322] = 16'b0000000000000000;
    assign weights1[6][323] = 16'b0000000000000000;
    assign weights1[6][324] = 16'b0000000000000000;
    assign weights1[6][325] = 16'b0000000000000000;
    assign weights1[6][326] = 16'b0000000000000000;
    assign weights1[6][327] = 16'b0000000000000000;
    assign weights1[6][328] = 16'b0000000000000000;
    assign weights1[6][329] = 16'b0000000000000000;
    assign weights1[6][330] = 16'b0000000000000000;
    assign weights1[6][331] = 16'b0000000000000000;
    assign weights1[6][332] = 16'b0000000000000000;
    assign weights1[6][333] = 16'b0000000000000000;
    assign weights1[6][334] = 16'b0000000000000000;
    assign weights1[6][335] = 16'b0000000000000000;
    assign weights1[6][336] = 16'b0000000000000000;
    assign weights1[6][337] = 16'b0000000000000000;
    assign weights1[6][338] = 16'b0000000000000000;
    assign weights1[6][339] = 16'b0000000000000000;
    assign weights1[6][340] = 16'b0000000000000000;
    assign weights1[6][341] = 16'b0000000000000000;
    assign weights1[6][342] = 16'b0000000000000000;
    assign weights1[6][343] = 16'b0000000000000000;
    assign weights1[6][344] = 16'b0000000000000000;
    assign weights1[6][345] = 16'b0000000000000000;
    assign weights1[6][346] = 16'b0000000000000000;
    assign weights1[6][347] = 16'b0000000000000000;
    assign weights1[6][348] = 16'b0000000000000000;
    assign weights1[6][349] = 16'b0000000000000000;
    assign weights1[6][350] = 16'b0000000000000000;
    assign weights1[6][351] = 16'b0000000000000000;
    assign weights1[6][352] = 16'b0000000000000000;
    assign weights1[6][353] = 16'b0000000000000000;
    assign weights1[6][354] = 16'b0000000000000000;
    assign weights1[6][355] = 16'b0000000000000000;
    assign weights1[6][356] = 16'b0000000000000000;
    assign weights1[6][357] = 16'b0000000000000000;
    assign weights1[6][358] = 16'b0000000000000000;
    assign weights1[6][359] = 16'b0000000000000000;
    assign weights1[6][360] = 16'b0000000000000000;
    assign weights1[6][361] = 16'b0000000000000000;
    assign weights1[6][362] = 16'b0000000000000000;
    assign weights1[6][363] = 16'b0000000000000000;
    assign weights1[6][364] = 16'b0000000000000000;
    assign weights1[6][365] = 16'b0000000000000000;
    assign weights1[6][366] = 16'b0000000000000000;
    assign weights1[6][367] = 16'b0000000000000000;
    assign weights1[6][368] = 16'b0000000000000000;
    assign weights1[6][369] = 16'b0000000000000000;
    assign weights1[6][370] = 16'b0000000000000000;
    assign weights1[6][371] = 16'b0000000000000000;
    assign weights1[6][372] = 16'b0000000000000000;
    assign weights1[6][373] = 16'b0000000000000000;
    assign weights1[6][374] = 16'b0000000000000000;
    assign weights1[6][375] = 16'b0000000000000000;
    assign weights1[6][376] = 16'b0000000000000000;
    assign weights1[6][377] = 16'b0000000000000000;
    assign weights1[6][378] = 16'b0000000000000000;
    assign weights1[6][379] = 16'b0000000000000000;
    assign weights1[6][380] = 16'b0000000000000000;
    assign weights1[6][381] = 16'b0000000000000000;
    assign weights1[6][382] = 16'b0000000000000000;
    assign weights1[6][383] = 16'b0000000000000000;
    assign weights1[6][384] = 16'b0000000000000000;
    assign weights1[6][385] = 16'b0000000000000000;
    assign weights1[6][386] = 16'b0000000000000000;
    assign weights1[6][387] = 16'b0000000000000000;
    assign weights1[6][388] = 16'b0000000000000000;
    assign weights1[6][389] = 16'b0000000000000000;
    assign weights1[6][390] = 16'b0000000000000000;
    assign weights1[6][391] = 16'b0000000000000000;
    assign weights1[6][392] = 16'b0000000000000000;
    assign weights1[6][393] = 16'b0000000000000000;
    assign weights1[6][394] = 16'b0000000000000000;
    assign weights1[6][395] = 16'b0000000000000000;
    assign weights1[6][396] = 16'b0000000000000000;
    assign weights1[6][397] = 16'b0000000000000000;
    assign weights1[6][398] = 16'b0000000000000000;
    assign weights1[6][399] = 16'b0000000000000000;
    assign weights1[6][400] = 16'b0000000000000000;
    assign weights1[6][401] = 16'b0000000000000000;
    assign weights1[6][402] = 16'b0000000000000000;
    assign weights1[6][403] = 16'b0000000000000000;
    assign weights1[6][404] = 16'b0000000000000000;
    assign weights1[6][405] = 16'b0000000000000000;
    assign weights1[6][406] = 16'b0000000000000000;
    assign weights1[6][407] = 16'b0000000000000000;
    assign weights1[6][408] = 16'b0000000000000000;
    assign weights1[6][409] = 16'b0000000000000000;
    assign weights1[6][410] = 16'b0000000000000000;
    assign weights1[6][411] = 16'b0000000000000000;
    assign weights1[6][412] = 16'b0000000000000000;
    assign weights1[6][413] = 16'b0000000000000000;
    assign weights1[6][414] = 16'b0000000000000000;
    assign weights1[6][415] = 16'b0000000000000000;
    assign weights1[6][416] = 16'b0000000000000000;
    assign weights1[6][417] = 16'b0000000000000000;
    assign weights1[6][418] = 16'b0000000000000000;
    assign weights1[6][419] = 16'b0000000000000000;
    assign weights1[6][420] = 16'b0000000000000000;
    assign weights1[6][421] = 16'b0000000000000000;
    assign weights1[6][422] = 16'b0000000000000000;
    assign weights1[6][423] = 16'b0000000000000000;
    assign weights1[6][424] = 16'b0000000000000000;
    assign weights1[6][425] = 16'b0000000000000000;
    assign weights1[6][426] = 16'b0000000000000000;
    assign weights1[6][427] = 16'b0000000000000000;
    assign weights1[6][428] = 16'b0000000000000000;
    assign weights1[6][429] = 16'b0000000000000000;
    assign weights1[6][430] = 16'b0000000000000000;
    assign weights1[6][431] = 16'b0000000000000000;
    assign weights1[6][432] = 16'b0000000000000000;
    assign weights1[6][433] = 16'b0000000000000000;
    assign weights1[6][434] = 16'b0000000000000000;
    assign weights1[6][435] = 16'b0000000000000000;
    assign weights1[6][436] = 16'b0000000000000000;
    assign weights1[6][437] = 16'b0000000000000000;
    assign weights1[6][438] = 16'b0000000000000000;
    assign weights1[6][439] = 16'b0000000000000000;
    assign weights1[6][440] = 16'b0000000000000000;
    assign weights1[6][441] = 16'b0000000000000000;
    assign weights1[6][442] = 16'b0000000000000000;
    assign weights1[6][443] = 16'b0000000000000000;
    assign weights1[6][444] = 16'b0000000000000000;
    assign weights1[6][445] = 16'b0000000000000000;
    assign weights1[6][446] = 16'b0000000000000000;
    assign weights1[6][447] = 16'b0000000000000000;
    assign weights1[6][448] = 16'b0000000000000000;
    assign weights1[6][449] = 16'b0000000000000000;
    assign weights1[6][450] = 16'b0000000000000000;
    assign weights1[6][451] = 16'b0000000000000000;
    assign weights1[6][452] = 16'b0000000000000000;
    assign weights1[6][453] = 16'b0000000000000000;
    assign weights1[6][454] = 16'b0000000000000000;
    assign weights1[6][455] = 16'b0000000000000000;
    assign weights1[6][456] = 16'b0000000000000000;
    assign weights1[6][457] = 16'b0000000000000000;
    assign weights1[6][458] = 16'b0000000000000000;
    assign weights1[6][459] = 16'b0000000000000000;
    assign weights1[6][460] = 16'b0000000000000000;
    assign weights1[6][461] = 16'b0000000000000000;
    assign weights1[6][462] = 16'b0000000000000000;
    assign weights1[6][463] = 16'b0000000000000000;
    assign weights1[6][464] = 16'b0000000000000000;
    assign weights1[6][465] = 16'b0000000000000000;
    assign weights1[6][466] = 16'b0000000000000000;
    assign weights1[6][467] = 16'b0000000000000000;
    assign weights1[6][468] = 16'b0000000000000000;
    assign weights1[6][469] = 16'b0000000000000000;
    assign weights1[6][470] = 16'b0000000000000000;
    assign weights1[6][471] = 16'b0000000000000000;
    assign weights1[6][472] = 16'b0000000000000000;
    assign weights1[6][473] = 16'b0000000000000000;
    assign weights1[6][474] = 16'b0000000000000000;
    assign weights1[6][475] = 16'b0000000000000000;
    assign weights1[6][476] = 16'b0000000000000000;
    assign weights1[6][477] = 16'b0000000000000000;
    assign weights1[6][478] = 16'b0000000000000000;
    assign weights1[6][479] = 16'b0000000000000000;
    assign weights1[6][480] = 16'b0000000000000000;
    assign weights1[6][481] = 16'b0000000000000000;
    assign weights1[6][482] = 16'b0000000000000000;
    assign weights1[6][483] = 16'b0000000000000000;
    assign weights1[6][484] = 16'b0000000000000000;
    assign weights1[6][485] = 16'b0000000000000000;
    assign weights1[6][486] = 16'b0000000000000000;
    assign weights1[6][487] = 16'b0000000000000000;
    assign weights1[6][488] = 16'b0000000000000000;
    assign weights1[6][489] = 16'b0000000000000000;
    assign weights1[6][490] = 16'b0000000000000000;
    assign weights1[6][491] = 16'b0000000000000000;
    assign weights1[6][492] = 16'b0000000000000000;
    assign weights1[6][493] = 16'b0000000000000000;
    assign weights1[6][494] = 16'b0000000000000000;
    assign weights1[6][495] = 16'b0000000000000000;
    assign weights1[6][496] = 16'b0000000000000000;
    assign weights1[6][497] = 16'b0000000000000000;
    assign weights1[6][498] = 16'b0000000000000000;
    assign weights1[6][499] = 16'b0000000000000000;
    assign weights1[6][500] = 16'b0000000000000000;
    assign weights1[6][501] = 16'b0000000000000000;
    assign weights1[6][502] = 16'b0000000000000000;
    assign weights1[6][503] = 16'b0000000000000000;
    assign weights1[6][504] = 16'b0000000000000000;
    assign weights1[6][505] = 16'b0000000000000000;
    assign weights1[6][506] = 16'b0000000000000000;
    assign weights1[6][507] = 16'b0000000000000000;
    assign weights1[6][508] = 16'b0000000000000000;
    assign weights1[6][509] = 16'b0000000000000000;
    assign weights1[6][510] = 16'b0000000000000000;
    assign weights1[6][511] = 16'b0000000000000000;
    assign weights1[6][512] = 16'b0000000000000000;
    assign weights1[6][513] = 16'b0000000000000000;
    assign weights1[6][514] = 16'b0000000000000000;
    assign weights1[6][515] = 16'b0000000000000000;
    assign weights1[6][516] = 16'b0000000000000000;
    assign weights1[6][517] = 16'b0000000000000000;
    assign weights1[6][518] = 16'b0000000000000000;
    assign weights1[6][519] = 16'b0000000000000000;
    assign weights1[6][520] = 16'b0000000000000000;
    assign weights1[6][521] = 16'b0000000000000000;
    assign weights1[6][522] = 16'b0000000000000000;
    assign weights1[6][523] = 16'b0000000000000000;
    assign weights1[6][524] = 16'b0000000000000000;
    assign weights1[6][525] = 16'b0000000000000000;
    assign weights1[6][526] = 16'b0000000000000000;
    assign weights1[6][527] = 16'b0000000000000000;
    assign weights1[6][528] = 16'b0000000000000000;
    assign weights1[6][529] = 16'b0000000000000000;
    assign weights1[6][530] = 16'b0000000000000000;
    assign weights1[6][531] = 16'b0000000000000000;
    assign weights1[6][532] = 16'b0000000000000000;
    assign weights1[6][533] = 16'b0000000000000000;
    assign weights1[6][534] = 16'b0000000000000000;
    assign weights1[6][535] = 16'b0000000000000000;
    assign weights1[6][536] = 16'b0000000000000000;
    assign weights1[6][537] = 16'b0000000000000000;
    assign weights1[6][538] = 16'b0000000000000000;
    assign weights1[6][539] = 16'b0000000000000000;
    assign weights1[6][540] = 16'b0000000000000000;
    assign weights1[6][541] = 16'b0000000000000000;
    assign weights1[6][542] = 16'b0000000000000000;
    assign weights1[6][543] = 16'b0000000000000000;
    assign weights1[6][544] = 16'b0000000000000000;
    assign weights1[6][545] = 16'b0000000000000000;
    assign weights1[6][546] = 16'b0000000000000000;
    assign weights1[6][547] = 16'b0000000000000000;
    assign weights1[6][548] = 16'b0000000000000000;
    assign weights1[6][549] = 16'b0000000000000000;
    assign weights1[6][550] = 16'b0000000000000000;
    assign weights1[6][551] = 16'b0000000000000000;
    assign weights1[6][552] = 16'b0000000000000000;
    assign weights1[6][553] = 16'b0000000000000000;
    assign weights1[6][554] = 16'b0000000000000000;
    assign weights1[6][555] = 16'b0000000000000000;
    assign weights1[6][556] = 16'b0000000000000000;
    assign weights1[6][557] = 16'b0000000000000000;
    assign weights1[6][558] = 16'b0000000000000000;
    assign weights1[6][559] = 16'b0000000000000000;
    assign weights1[6][560] = 16'b0000000000000000;
    assign weights1[6][561] = 16'b0000000000000000;
    assign weights1[6][562] = 16'b0000000000000000;
    assign weights1[6][563] = 16'b0000000000000000;
    assign weights1[6][564] = 16'b0000000000000000;
    assign weights1[6][565] = 16'b0000000000000000;
    assign weights1[6][566] = 16'b0000000000000000;
    assign weights1[6][567] = 16'b0000000000000000;
    assign weights1[6][568] = 16'b0000000000000000;
    assign weights1[6][569] = 16'b0000000000000000;
    assign weights1[6][570] = 16'b0000000000000000;
    assign weights1[6][571] = 16'b0000000000000000;
    assign weights1[6][572] = 16'b0000000000000000;
    assign weights1[6][573] = 16'b0000000000000000;
    assign weights1[6][574] = 16'b0000000000000000;
    assign weights1[6][575] = 16'b0000000000000000;
    assign weights1[6][576] = 16'b0000000000000000;
    assign weights1[6][577] = 16'b0000000000000000;
    assign weights1[6][578] = 16'b0000000000000000;
    assign weights1[6][579] = 16'b0000000000000000;
    assign weights1[6][580] = 16'b0000000000000000;
    assign weights1[6][581] = 16'b0000000000000000;
    assign weights1[6][582] = 16'b0000000000000000;
    assign weights1[6][583] = 16'b0000000000000000;
    assign weights1[6][584] = 16'b0000000000000000;
    assign weights1[6][585] = 16'b0000000000000000;
    assign weights1[6][586] = 16'b0000000000000000;
    assign weights1[6][587] = 16'b0000000000000000;
    assign weights1[6][588] = 16'b0000000000000000;
    assign weights1[6][589] = 16'b0000000000000000;
    assign weights1[6][590] = 16'b0000000000000000;
    assign weights1[6][591] = 16'b0000000000000000;
    assign weights1[6][592] = 16'b0000000000000000;
    assign weights1[6][593] = 16'b0000000000000000;
    assign weights1[6][594] = 16'b0000000000000000;
    assign weights1[6][595] = 16'b0000000000000000;
    assign weights1[6][596] = 16'b0000000000000000;
    assign weights1[6][597] = 16'b0000000000000000;
    assign weights1[6][598] = 16'b0000000000000000;
    assign weights1[6][599] = 16'b0000000000000000;
    assign weights1[6][600] = 16'b0000000000000000;
    assign weights1[6][601] = 16'b0000000000000000;
    assign weights1[6][602] = 16'b0000000000000000;
    assign weights1[6][603] = 16'b0000000000000000;
    assign weights1[6][604] = 16'b0000000000000000;
    assign weights1[6][605] = 16'b0000000000000000;
    assign weights1[6][606] = 16'b0000000000000000;
    assign weights1[6][607] = 16'b0000000000000000;
    assign weights1[6][608] = 16'b0000000000000000;
    assign weights1[6][609] = 16'b0000000000000000;
    assign weights1[6][610] = 16'b0000000000000000;
    assign weights1[6][611] = 16'b0000000000000000;
    assign weights1[6][612] = 16'b0000000000000000;
    assign weights1[6][613] = 16'b0000000000000000;
    assign weights1[6][614] = 16'b0000000000000000;
    assign weights1[6][615] = 16'b0000000000000000;
    assign weights1[6][616] = 16'b0000000000000000;
    assign weights1[6][617] = 16'b0000000000000000;
    assign weights1[6][618] = 16'b0000000000000000;
    assign weights1[6][619] = 16'b0000000000000000;
    assign weights1[6][620] = 16'b0000000000000000;
    assign weights1[6][621] = 16'b0000000000000000;
    assign weights1[6][622] = 16'b0000000000000000;
    assign weights1[6][623] = 16'b0000000000000000;
    assign weights1[6][624] = 16'b0000000000000000;
    assign weights1[6][625] = 16'b0000000000000000;
    assign weights1[6][626] = 16'b0000000000000000;
    assign weights1[6][627] = 16'b0000000000000000;
    assign weights1[6][628] = 16'b0000000000000000;
    assign weights1[6][629] = 16'b0000000000000000;
    assign weights1[6][630] = 16'b0000000000000000;
    assign weights1[6][631] = 16'b0000000000000000;
    assign weights1[6][632] = 16'b0000000000000000;
    assign weights1[6][633] = 16'b0000000000000000;
    assign weights1[6][634] = 16'b0000000000000000;
    assign weights1[6][635] = 16'b0000000000000000;
    assign weights1[6][636] = 16'b0000000000000000;
    assign weights1[6][637] = 16'b0000000000000000;
    assign weights1[6][638] = 16'b0000000000000000;
    assign weights1[6][639] = 16'b0000000000000000;
    assign weights1[6][640] = 16'b0000000000000000;
    assign weights1[6][641] = 16'b0000000000000000;
    assign weights1[6][642] = 16'b0000000000000000;
    assign weights1[6][643] = 16'b0000000000000000;
    assign weights1[6][644] = 16'b0000000000000000;
    assign weights1[6][645] = 16'b0000000000000000;
    assign weights1[6][646] = 16'b0000000000000000;
    assign weights1[6][647] = 16'b0000000000000000;
    assign weights1[6][648] = 16'b0000000000000000;
    assign weights1[6][649] = 16'b0000000000000000;
    assign weights1[6][650] = 16'b0000000000000000;
    assign weights1[6][651] = 16'b0000000000000000;
    assign weights1[6][652] = 16'b0000000000000000;
    assign weights1[6][653] = 16'b0000000000000000;
    assign weights1[6][654] = 16'b0000000000000000;
    assign weights1[6][655] = 16'b0000000000000000;
    assign weights1[6][656] = 16'b0000000000000000;
    assign weights1[6][657] = 16'b0000000000000000;
    assign weights1[6][658] = 16'b0000000000000000;
    assign weights1[6][659] = 16'b0000000000000000;
    assign weights1[6][660] = 16'b0000000000000000;
    assign weights1[6][661] = 16'b0000000000000000;
    assign weights1[6][662] = 16'b0000000000000000;
    assign weights1[6][663] = 16'b0000000000000000;
    assign weights1[6][664] = 16'b0000000000000000;
    assign weights1[6][665] = 16'b0000000000000000;
    assign weights1[6][666] = 16'b0000000000000000;
    assign weights1[6][667] = 16'b0000000000000000;
    assign weights1[6][668] = 16'b0000000000000000;
    assign weights1[6][669] = 16'b0000000000000000;
    assign weights1[6][670] = 16'b0000000000000000;
    assign weights1[6][671] = 16'b0000000000000000;
    assign weights1[6][672] = 16'b0000000000000000;
    assign weights1[6][673] = 16'b0000000000000000;
    assign weights1[6][674] = 16'b0000000000000000;
    assign weights1[6][675] = 16'b0000000000000000;
    assign weights1[6][676] = 16'b0000000000000000;
    assign weights1[6][677] = 16'b0000000000000000;
    assign weights1[6][678] = 16'b0000000000000000;
    assign weights1[6][679] = 16'b0000000000000000;
    assign weights1[6][680] = 16'b0000000000000000;
    assign weights1[6][681] = 16'b0000000000000000;
    assign weights1[6][682] = 16'b0000000000000000;
    assign weights1[6][683] = 16'b0000000000000000;
    assign weights1[6][684] = 16'b0000000000000000;
    assign weights1[6][685] = 16'b0000000000000000;
    assign weights1[6][686] = 16'b0000000000000000;
    assign weights1[6][687] = 16'b0000000000000000;
    assign weights1[6][688] = 16'b0000000000000000;
    assign weights1[6][689] = 16'b0000000000000000;
    assign weights1[6][690] = 16'b0000000000000000;
    assign weights1[6][691] = 16'b0000000000000000;
    assign weights1[6][692] = 16'b0000000000000000;
    assign weights1[6][693] = 16'b0000000000000000;
    assign weights1[6][694] = 16'b0000000000000000;
    assign weights1[6][695] = 16'b0000000000000000;
    assign weights1[6][696] = 16'b0000000000000000;
    assign weights1[6][697] = 16'b0000000000000000;
    assign weights1[6][698] = 16'b0000000000000000;
    assign weights1[6][699] = 16'b0000000000000000;
    assign weights1[6][700] = 16'b0000000000000000;
    assign weights1[6][701] = 16'b0000000000000000;
    assign weights1[6][702] = 16'b0000000000000000;
    assign weights1[6][703] = 16'b0000000000000000;
    assign weights1[6][704] = 16'b0000000000000000;
    assign weights1[6][705] = 16'b0000000000000000;
    assign weights1[6][706] = 16'b0000000000000000;
    assign weights1[6][707] = 16'b0000000000000000;
    assign weights1[6][708] = 16'b0000000000000000;
    assign weights1[6][709] = 16'b0000000000000000;
    assign weights1[6][710] = 16'b0000000000000000;
    assign weights1[6][711] = 16'b0000000000000000;
    assign weights1[6][712] = 16'b0000000000000000;
    assign weights1[6][713] = 16'b0000000000000000;
    assign weights1[6][714] = 16'b0000000000000000;
    assign weights1[6][715] = 16'b0000000000000000;
    assign weights1[6][716] = 16'b0000000000000000;
    assign weights1[6][717] = 16'b0000000000000000;
    assign weights1[6][718] = 16'b0000000000000000;
    assign weights1[6][719] = 16'b0000000000000000;
    assign weights1[6][720] = 16'b0000000000000000;
    assign weights1[6][721] = 16'b0000000000000000;
    assign weights1[6][722] = 16'b0000000000000000;
    assign weights1[6][723] = 16'b0000000000000000;
    assign weights1[6][724] = 16'b0000000000000000;
    assign weights1[6][725] = 16'b0000000000000000;
    assign weights1[6][726] = 16'b0000000000000000;
    assign weights1[6][727] = 16'b0000000000000000;
    assign weights1[6][728] = 16'b0000000000000000;
    assign weights1[6][729] = 16'b0000000000000000;
    assign weights1[6][730] = 16'b0000000000000000;
    assign weights1[6][731] = 16'b0000000000000000;
    assign weights1[6][732] = 16'b0000000000000000;
    assign weights1[6][733] = 16'b0000000000000000;
    assign weights1[6][734] = 16'b0000000000000000;
    assign weights1[6][735] = 16'b0000000000000000;
    assign weights1[6][736] = 16'b0000000000000000;
    assign weights1[6][737] = 16'b0000000000000000;
    assign weights1[6][738] = 16'b0000000000000000;
    assign weights1[6][739] = 16'b0000000000000000;
    assign weights1[6][740] = 16'b0000000000000000;
    assign weights1[6][741] = 16'b0000000000000000;
    assign weights1[6][742] = 16'b0000000000000000;
    assign weights1[6][743] = 16'b0000000000000000;
    assign weights1[6][744] = 16'b0000000000000000;
    assign weights1[6][745] = 16'b0000000000000000;
    assign weights1[6][746] = 16'b0000000000000000;
    assign weights1[6][747] = 16'b0000000000000000;
    assign weights1[6][748] = 16'b0000000000000000;
    assign weights1[6][749] = 16'b0000000000000000;
    assign weights1[6][750] = 16'b0000000000000000;
    assign weights1[6][751] = 16'b0000000000000000;
    assign weights1[6][752] = 16'b0000000000000000;
    assign weights1[6][753] = 16'b0000000000000000;
    assign weights1[6][754] = 16'b0000000000000000;
    assign weights1[6][755] = 16'b0000000000000000;
    assign weights1[6][756] = 16'b0000000000000000;
    assign weights1[6][757] = 16'b0000000000000000;
    assign weights1[6][758] = 16'b0000000000000000;
    assign weights1[6][759] = 16'b0000000000000000;
    assign weights1[6][760] = 16'b0000000000000000;
    assign weights1[6][761] = 16'b0000000000000000;
    assign weights1[6][762] = 16'b0000000000000000;
    assign weights1[6][763] = 16'b0000000000000000;
    assign weights1[6][764] = 16'b0000000000000000;
    assign weights1[6][765] = 16'b0000000000000000;
    assign weights1[6][766] = 16'b0000000000000000;
    assign weights1[6][767] = 16'b0000000000000000;
    assign weights1[6][768] = 16'b0000000000000000;
    assign weights1[6][769] = 16'b0000000000000000;
    assign weights1[6][770] = 16'b0000000000000000;
    assign weights1[6][771] = 16'b0000000000000000;
    assign weights1[6][772] = 16'b0000000000000000;
    assign weights1[6][773] = 16'b0000000000000000;
    assign weights1[6][774] = 16'b0000000000000000;
    assign weights1[6][775] = 16'b0000000000000000;
    assign weights1[6][776] = 16'b0000000000000000;
    assign weights1[6][777] = 16'b0000000000000000;
    assign weights1[6][778] = 16'b0000000000000000;
    assign weights1[6][779] = 16'b0000000000000000;
    assign weights1[6][780] = 16'b0000000000000000;
    assign weights1[6][781] = 16'b0000000000000000;
    assign weights1[6][782] = 16'b0000000000000000;
    assign weights1[6][783] = 16'b0000000000000000;
    assign weights1[7][0] = 16'b0000000000000000;
    assign weights1[7][1] = 16'b0000000000000000;
    assign weights1[7][2] = 16'b0000000000000000;
    assign weights1[7][3] = 16'b0000000000000010;
    assign weights1[7][4] = 16'b1111111111111111;
    assign weights1[7][5] = 16'b1111111111111101;
    assign weights1[7][6] = 16'b1111111111111000;
    assign weights1[7][7] = 16'b1111111111110011;
    assign weights1[7][8] = 16'b1111111111111010;
    assign weights1[7][9] = 16'b1111111111110010;
    assign weights1[7][10] = 16'b1111111111011110;
    assign weights1[7][11] = 16'b1111111111101111;
    assign weights1[7][12] = 16'b1111111111111110;
    assign weights1[7][13] = 16'b1111111111111111;
    assign weights1[7][14] = 16'b0000000000001001;
    assign weights1[7][15] = 16'b0000000000000101;
    assign weights1[7][16] = 16'b1111111111110111;
    assign weights1[7][17] = 16'b1111111111111101;
    assign weights1[7][18] = 16'b1111111111110100;
    assign weights1[7][19] = 16'b1111111111101100;
    assign weights1[7][20] = 16'b1111111111110111;
    assign weights1[7][21] = 16'b0000000000000000;
    assign weights1[7][22] = 16'b0000000000000100;
    assign weights1[7][23] = 16'b0000000000000011;
    assign weights1[7][24] = 16'b0000000000000000;
    assign weights1[7][25] = 16'b0000000000000010;
    assign weights1[7][26] = 16'b0000000000000011;
    assign weights1[7][27] = 16'b0000000000000000;
    assign weights1[7][28] = 16'b0000000000000001;
    assign weights1[7][29] = 16'b0000000000000001;
    assign weights1[7][30] = 16'b0000000000000001;
    assign weights1[7][31] = 16'b1111111111111101;
    assign weights1[7][32] = 16'b1111111111111000;
    assign weights1[7][33] = 16'b1111111111111011;
    assign weights1[7][34] = 16'b1111111111111000;
    assign weights1[7][35] = 16'b1111111111110011;
    assign weights1[7][36] = 16'b1111111111111100;
    assign weights1[7][37] = 16'b1111111111111011;
    assign weights1[7][38] = 16'b1111111111101110;
    assign weights1[7][39] = 16'b1111111111111111;
    assign weights1[7][40] = 16'b1111111111111111;
    assign weights1[7][41] = 16'b1111111111110101;
    assign weights1[7][42] = 16'b0000000000000011;
    assign weights1[7][43] = 16'b1111111111110001;
    assign weights1[7][44] = 16'b1111111111110110;
    assign weights1[7][45] = 16'b1111111111111010;
    assign weights1[7][46] = 16'b0000000000000101;
    assign weights1[7][47] = 16'b1111111111110101;
    assign weights1[7][48] = 16'b1111111111110110;
    assign weights1[7][49] = 16'b1111111111111101;
    assign weights1[7][50] = 16'b1111111111111100;
    assign weights1[7][51] = 16'b0000000000000000;
    assign weights1[7][52] = 16'b1111111111111110;
    assign weights1[7][53] = 16'b0000000000000101;
    assign weights1[7][54] = 16'b0000000000000010;
    assign weights1[7][55] = 16'b0000000000000011;
    assign weights1[7][56] = 16'b0000000000000001;
    assign weights1[7][57] = 16'b0000000000000001;
    assign weights1[7][58] = 16'b1111111111111100;
    assign weights1[7][59] = 16'b1111111111111100;
    assign weights1[7][60] = 16'b1111111111110011;
    assign weights1[7][61] = 16'b1111111111110000;
    assign weights1[7][62] = 16'b1111111111110000;
    assign weights1[7][63] = 16'b1111111111110011;
    assign weights1[7][64] = 16'b1111111111110011;
    assign weights1[7][65] = 16'b1111111111110101;
    assign weights1[7][66] = 16'b1111111111111101;
    assign weights1[7][67] = 16'b1111111111111010;
    assign weights1[7][68] = 16'b1111111111111000;
    assign weights1[7][69] = 16'b0000000000000001;
    assign weights1[7][70] = 16'b1111111111110110;
    assign weights1[7][71] = 16'b0000000000000010;
    assign weights1[7][72] = 16'b1111111111110010;
    assign weights1[7][73] = 16'b1111111111110101;
    assign weights1[7][74] = 16'b1111111111111111;
    assign weights1[7][75] = 16'b0000000000000010;
    assign weights1[7][76] = 16'b0000000000000011;
    assign weights1[7][77] = 16'b1111111111111110;
    assign weights1[7][78] = 16'b1111111111111010;
    assign weights1[7][79] = 16'b1111111111111110;
    assign weights1[7][80] = 16'b1111111111111110;
    assign weights1[7][81] = 16'b0000000000000001;
    assign weights1[7][82] = 16'b0000000000000010;
    assign weights1[7][83] = 16'b0000000000000010;
    assign weights1[7][84] = 16'b0000000000000001;
    assign weights1[7][85] = 16'b0000000000000001;
    assign weights1[7][86] = 16'b0000000000000010;
    assign weights1[7][87] = 16'b1111111111111001;
    assign weights1[7][88] = 16'b1111111111111000;
    assign weights1[7][89] = 16'b1111111111110000;
    assign weights1[7][90] = 16'b1111111111101001;
    assign weights1[7][91] = 16'b1111111111111101;
    assign weights1[7][92] = 16'b1111111111101011;
    assign weights1[7][93] = 16'b0000000000000101;
    assign weights1[7][94] = 16'b1111111111111100;
    assign weights1[7][95] = 16'b0000000000001011;
    assign weights1[7][96] = 16'b1111111111111011;
    assign weights1[7][97] = 16'b0000000000011110;
    assign weights1[7][98] = 16'b0000000000000110;
    assign weights1[7][99] = 16'b0000000000000000;
    assign weights1[7][100] = 16'b1111111111111011;
    assign weights1[7][101] = 16'b1111111111110101;
    assign weights1[7][102] = 16'b0000000000000000;
    assign weights1[7][103] = 16'b1111111111110111;
    assign weights1[7][104] = 16'b0000000000001010;
    assign weights1[7][105] = 16'b1111111111111100;
    assign weights1[7][106] = 16'b0000000000000001;
    assign weights1[7][107] = 16'b1111111111101000;
    assign weights1[7][108] = 16'b1111111111101001;
    assign weights1[7][109] = 16'b1111111111110011;
    assign weights1[7][110] = 16'b1111111111110010;
    assign weights1[7][111] = 16'b0000000000000001;
    assign weights1[7][112] = 16'b0000000000000000;
    assign weights1[7][113] = 16'b0000000000000000;
    assign weights1[7][114] = 16'b1111111111111101;
    assign weights1[7][115] = 16'b1111111111101111;
    assign weights1[7][116] = 16'b0000000000000011;
    assign weights1[7][117] = 16'b1111111111110100;
    assign weights1[7][118] = 16'b1111111111110100;
    assign weights1[7][119] = 16'b1111111111110011;
    assign weights1[7][120] = 16'b0000000000000011;
    assign weights1[7][121] = 16'b1111111111110010;
    assign weights1[7][122] = 16'b1111111111100111;
    assign weights1[7][123] = 16'b1111111111100110;
    assign weights1[7][124] = 16'b0000000000000100;
    assign weights1[7][125] = 16'b1111111111111110;
    assign weights1[7][126] = 16'b1111111111101011;
    assign weights1[7][127] = 16'b1111111111111111;
    assign weights1[7][128] = 16'b1111111111110101;
    assign weights1[7][129] = 16'b0000000000001101;
    assign weights1[7][130] = 16'b0000000000000110;
    assign weights1[7][131] = 16'b1111111111111111;
    assign weights1[7][132] = 16'b1111111111101100;
    assign weights1[7][133] = 16'b1111111111101110;
    assign weights1[7][134] = 16'b1111111111111000;
    assign weights1[7][135] = 16'b0000000000010111;
    assign weights1[7][136] = 16'b1111111111111100;
    assign weights1[7][137] = 16'b1111111111101110;
    assign weights1[7][138] = 16'b1111111111110111;
    assign weights1[7][139] = 16'b1111111111111000;
    assign weights1[7][140] = 16'b1111111111111110;
    assign weights1[7][141] = 16'b1111111111111001;
    assign weights1[7][142] = 16'b1111111111111101;
    assign weights1[7][143] = 16'b1111111111110010;
    assign weights1[7][144] = 16'b1111111111110010;
    assign weights1[7][145] = 16'b1111111111100110;
    assign weights1[7][146] = 16'b1111111111110111;
    assign weights1[7][147] = 16'b1111111111101111;
    assign weights1[7][148] = 16'b1111111111110011;
    assign weights1[7][149] = 16'b0000000000000101;
    assign weights1[7][150] = 16'b1111111111111001;
    assign weights1[7][151] = 16'b0000000000000111;
    assign weights1[7][152] = 16'b1111111111111111;
    assign weights1[7][153] = 16'b0000000000010001;
    assign weights1[7][154] = 16'b1111111111111010;
    assign weights1[7][155] = 16'b1111111111110101;
    assign weights1[7][156] = 16'b1111111111111101;
    assign weights1[7][157] = 16'b1111111111110001;
    assign weights1[7][158] = 16'b1111111111101011;
    assign weights1[7][159] = 16'b1111111111111101;
    assign weights1[7][160] = 16'b1111111111011010;
    assign weights1[7][161] = 16'b1111111111110101;
    assign weights1[7][162] = 16'b1111111111111000;
    assign weights1[7][163] = 16'b1111111111110100;
    assign weights1[7][164] = 16'b1111111111111011;
    assign weights1[7][165] = 16'b1111111111111110;
    assign weights1[7][166] = 16'b1111111111110000;
    assign weights1[7][167] = 16'b1111111111110101;
    assign weights1[7][168] = 16'b1111111111111001;
    assign weights1[7][169] = 16'b1111111111111010;
    assign weights1[7][170] = 16'b0000000000001011;
    assign weights1[7][171] = 16'b1111111111110001;
    assign weights1[7][172] = 16'b0000000000000010;
    assign weights1[7][173] = 16'b0000000000000110;
    assign weights1[7][174] = 16'b0000000000010011;
    assign weights1[7][175] = 16'b1111111111110100;
    assign weights1[7][176] = 16'b1111111111111101;
    assign weights1[7][177] = 16'b0000000000001010;
    assign weights1[7][178] = 16'b0000000000000000;
    assign weights1[7][179] = 16'b0000000000000011;
    assign weights1[7][180] = 16'b1111111111111101;
    assign weights1[7][181] = 16'b1111111111111010;
    assign weights1[7][182] = 16'b0000000000010101;
    assign weights1[7][183] = 16'b0000000000001001;
    assign weights1[7][184] = 16'b0000000000001011;
    assign weights1[7][185] = 16'b0000000000001001;
    assign weights1[7][186] = 16'b0000000000000001;
    assign weights1[7][187] = 16'b1111111111101110;
    assign weights1[7][188] = 16'b1111111111110111;
    assign weights1[7][189] = 16'b1111111111111100;
    assign weights1[7][190] = 16'b1111111111110101;
    assign weights1[7][191] = 16'b0000000000000111;
    assign weights1[7][192] = 16'b1111111111111110;
    assign weights1[7][193] = 16'b1111111111111111;
    assign weights1[7][194] = 16'b1111111111110111;
    assign weights1[7][195] = 16'b1111111111110010;
    assign weights1[7][196] = 16'b1111111111111101;
    assign weights1[7][197] = 16'b1111111111110100;
    assign weights1[7][198] = 16'b1111111111111000;
    assign weights1[7][199] = 16'b1111111111111101;
    assign weights1[7][200] = 16'b1111111111111110;
    assign weights1[7][201] = 16'b1111111111111110;
    assign weights1[7][202] = 16'b0000000000000101;
    assign weights1[7][203] = 16'b0000000000000001;
    assign weights1[7][204] = 16'b1111111111111111;
    assign weights1[7][205] = 16'b1111111111101111;
    assign weights1[7][206] = 16'b1111111111111010;
    assign weights1[7][207] = 16'b0000000000001101;
    assign weights1[7][208] = 16'b1111111111111111;
    assign weights1[7][209] = 16'b1111111111111100;
    assign weights1[7][210] = 16'b1111111111110110;
    assign weights1[7][211] = 16'b1111111111111001;
    assign weights1[7][212] = 16'b1111111111111000;
    assign weights1[7][213] = 16'b0000000000000000;
    assign weights1[7][214] = 16'b0000000000000110;
    assign weights1[7][215] = 16'b1111111111111110;
    assign weights1[7][216] = 16'b0000000000010010;
    assign weights1[7][217] = 16'b0000000000001101;
    assign weights1[7][218] = 16'b0000000000001100;
    assign weights1[7][219] = 16'b1111111111110110;
    assign weights1[7][220] = 16'b1111111111111101;
    assign weights1[7][221] = 16'b0000000000001111;
    assign weights1[7][222] = 16'b1111111111101101;
    assign weights1[7][223] = 16'b1111111111111100;
    assign weights1[7][224] = 16'b1111111111111000;
    assign weights1[7][225] = 16'b1111111111110100;
    assign weights1[7][226] = 16'b1111111111111100;
    assign weights1[7][227] = 16'b1111111111111101;
    assign weights1[7][228] = 16'b1111111111110111;
    assign weights1[7][229] = 16'b1111111111111011;
    assign weights1[7][230] = 16'b0000000000000100;
    assign weights1[7][231] = 16'b0000000000000110;
    assign weights1[7][232] = 16'b1111111111110000;
    assign weights1[7][233] = 16'b1111111111111010;
    assign weights1[7][234] = 16'b1111111111111000;
    assign weights1[7][235] = 16'b1111111111110001;
    assign weights1[7][236] = 16'b0000000000000101;
    assign weights1[7][237] = 16'b1111111111111100;
    assign weights1[7][238] = 16'b0000000000010100;
    assign weights1[7][239] = 16'b0000000000001111;
    assign weights1[7][240] = 16'b0000000000010110;
    assign weights1[7][241] = 16'b0000000000100111;
    assign weights1[7][242] = 16'b0000000000001101;
    assign weights1[7][243] = 16'b0000000000001010;
    assign weights1[7][244] = 16'b0000000000000110;
    assign weights1[7][245] = 16'b0000000000100111;
    assign weights1[7][246] = 16'b0000000000010110;
    assign weights1[7][247] = 16'b0000000000010010;
    assign weights1[7][248] = 16'b0000000000011001;
    assign weights1[7][249] = 16'b0000000000001101;
    assign weights1[7][250] = 16'b0000000000000110;
    assign weights1[7][251] = 16'b0000000000110000;
    assign weights1[7][252] = 16'b1111111111110110;
    assign weights1[7][253] = 16'b0000000000000000;
    assign weights1[7][254] = 16'b1111111111111111;
    assign weights1[7][255] = 16'b1111111111110101;
    assign weights1[7][256] = 16'b1111111111111101;
    assign weights1[7][257] = 16'b0000000000000010;
    assign weights1[7][258] = 16'b1111111111110001;
    assign weights1[7][259] = 16'b1111111111111011;
    assign weights1[7][260] = 16'b1111111111111110;
    assign weights1[7][261] = 16'b0000000000000000;
    assign weights1[7][262] = 16'b1111111111111011;
    assign weights1[7][263] = 16'b1111111111110010;
    assign weights1[7][264] = 16'b1111111111111000;
    assign weights1[7][265] = 16'b1111111111111011;
    assign weights1[7][266] = 16'b0000000000000000;
    assign weights1[7][267] = 16'b0000000000011001;
    assign weights1[7][268] = 16'b0000000000000011;
    assign weights1[7][269] = 16'b0000000000001110;
    assign weights1[7][270] = 16'b0000000000000110;
    assign weights1[7][271] = 16'b0000000000011100;
    assign weights1[7][272] = 16'b0000000000000111;
    assign weights1[7][273] = 16'b0000000000100001;
    assign weights1[7][274] = 16'b1111111111111101;
    assign weights1[7][275] = 16'b0000000000100010;
    assign weights1[7][276] = 16'b0000000000111000;
    assign weights1[7][277] = 16'b0000000000101101;
    assign weights1[7][278] = 16'b0000000000011111;
    assign weights1[7][279] = 16'b0000000001000000;
    assign weights1[7][280] = 16'b1111111111101110;
    assign weights1[7][281] = 16'b0000000000000011;
    assign weights1[7][282] = 16'b1111111111110110;
    assign weights1[7][283] = 16'b1111111111110010;
    assign weights1[7][284] = 16'b1111111111110101;
    assign weights1[7][285] = 16'b0000000000010110;
    assign weights1[7][286] = 16'b1111111111111001;
    assign weights1[7][287] = 16'b0000000000001010;
    assign weights1[7][288] = 16'b1111111111110011;
    assign weights1[7][289] = 16'b0000000000000011;
    assign weights1[7][290] = 16'b1111111111110000;
    assign weights1[7][291] = 16'b0000000000001000;
    assign weights1[7][292] = 16'b1111111111101111;
    assign weights1[7][293] = 16'b1111111111111100;
    assign weights1[7][294] = 16'b0000000000000000;
    assign weights1[7][295] = 16'b0000000000010010;
    assign weights1[7][296] = 16'b0000000000001011;
    assign weights1[7][297] = 16'b0000000000001101;
    assign weights1[7][298] = 16'b0000000000100001;
    assign weights1[7][299] = 16'b0000000000100000;
    assign weights1[7][300] = 16'b0000000000001000;
    assign weights1[7][301] = 16'b1111111111111111;
    assign weights1[7][302] = 16'b1111111111101010;
    assign weights1[7][303] = 16'b0000000000100001;
    assign weights1[7][304] = 16'b0000000001011000;
    assign weights1[7][305] = 16'b0000000000111110;
    assign weights1[7][306] = 16'b0000000000110101;
    assign weights1[7][307] = 16'b0000000000110011;
    assign weights1[7][308] = 16'b1111111111110011;
    assign weights1[7][309] = 16'b1111111111110111;
    assign weights1[7][310] = 16'b0000000000000111;
    assign weights1[7][311] = 16'b1111111111111101;
    assign weights1[7][312] = 16'b1111111111110011;
    assign weights1[7][313] = 16'b0000000000000001;
    assign weights1[7][314] = 16'b0000000000001101;
    assign weights1[7][315] = 16'b1111111111110001;
    assign weights1[7][316] = 16'b0000000000001010;
    assign weights1[7][317] = 16'b0000000000000010;
    assign weights1[7][318] = 16'b1111111111111111;
    assign weights1[7][319] = 16'b1111111111100100;
    assign weights1[7][320] = 16'b1111111111100001;
    assign weights1[7][321] = 16'b1111111111111000;
    assign weights1[7][322] = 16'b1111111111110011;
    assign weights1[7][323] = 16'b0000000000001001;
    assign weights1[7][324] = 16'b0000000000011101;
    assign weights1[7][325] = 16'b0000000000100101;
    assign weights1[7][326] = 16'b0000000000110110;
    assign weights1[7][327] = 16'b0000000000110110;
    assign weights1[7][328] = 16'b0000000000111110;
    assign weights1[7][329] = 16'b0000000001010000;
    assign weights1[7][330] = 16'b0000000000110011;
    assign weights1[7][331] = 16'b0000000001010101;
    assign weights1[7][332] = 16'b0000000000111001;
    assign weights1[7][333] = 16'b0000000000111100;
    assign weights1[7][334] = 16'b0000000000101001;
    assign weights1[7][335] = 16'b0000000000010110;
    assign weights1[7][336] = 16'b1111111111111010;
    assign weights1[7][337] = 16'b1111111111110111;
    assign weights1[7][338] = 16'b0000000000001100;
    assign weights1[7][339] = 16'b1111111111111001;
    assign weights1[7][340] = 16'b1111111111110111;
    assign weights1[7][341] = 16'b0000000000001010;
    assign weights1[7][342] = 16'b0000000000000111;
    assign weights1[7][343] = 16'b0000000000001001;
    assign weights1[7][344] = 16'b0000000000010110;
    assign weights1[7][345] = 16'b0000000000010001;
    assign weights1[7][346] = 16'b0000000000001100;
    assign weights1[7][347] = 16'b1111111111111000;
    assign weights1[7][348] = 16'b1111111111101000;
    assign weights1[7][349] = 16'b1111111110110010;
    assign weights1[7][350] = 16'b1111111111001000;
    assign weights1[7][351] = 16'b1111111111110110;
    assign weights1[7][352] = 16'b0000000000000010;
    assign weights1[7][353] = 16'b0000000000011100;
    assign weights1[7][354] = 16'b0000000000101000;
    assign weights1[7][355] = 16'b0000000000101000;
    assign weights1[7][356] = 16'b0000000001001111;
    assign weights1[7][357] = 16'b0000000001001101;
    assign weights1[7][358] = 16'b0000000001011100;
    assign weights1[7][359] = 16'b0000000000100101;
    assign weights1[7][360] = 16'b0000000000111100;
    assign weights1[7][361] = 16'b0000000000110010;
    assign weights1[7][362] = 16'b0000000000010010;
    assign weights1[7][363] = 16'b0000000000010010;
    assign weights1[7][364] = 16'b0000000000000001;
    assign weights1[7][365] = 16'b1111111111111000;
    assign weights1[7][366] = 16'b0000000000000100;
    assign weights1[7][367] = 16'b0000000000001001;
    assign weights1[7][368] = 16'b1111111111111001;
    assign weights1[7][369] = 16'b1111111111111000;
    assign weights1[7][370] = 16'b0000000000000100;
    assign weights1[7][371] = 16'b0000000000000000;
    assign weights1[7][372] = 16'b0000000000010010;
    assign weights1[7][373] = 16'b0000000000000110;
    assign weights1[7][374] = 16'b0000000000010111;
    assign weights1[7][375] = 16'b0000000000100100;
    assign weights1[7][376] = 16'b1111111111101000;
    assign weights1[7][377] = 16'b1111111111000101;
    assign weights1[7][378] = 16'b1111111101111110;
    assign weights1[7][379] = 16'b1111111110001011;
    assign weights1[7][380] = 16'b1111111110011100;
    assign weights1[7][381] = 16'b1111111110101000;
    assign weights1[7][382] = 16'b1111111111011110;
    assign weights1[7][383] = 16'b1111111111101100;
    assign weights1[7][384] = 16'b1111111111111101;
    assign weights1[7][385] = 16'b0000000000001100;
    assign weights1[7][386] = 16'b1111111111111010;
    assign weights1[7][387] = 16'b0000000000001101;
    assign weights1[7][388] = 16'b1111111111110110;
    assign weights1[7][389] = 16'b0000000000000110;
    assign weights1[7][390] = 16'b1111111111101000;
    assign weights1[7][391] = 16'b1111111111101101;
    assign weights1[7][392] = 16'b0000000000001100;
    assign weights1[7][393] = 16'b0000000000000010;
    assign weights1[7][394] = 16'b0000000000000010;
    assign weights1[7][395] = 16'b0000000000001001;
    assign weights1[7][396] = 16'b1111111111110111;
    assign weights1[7][397] = 16'b1111111111110101;
    assign weights1[7][398] = 16'b1111111111110101;
    assign weights1[7][399] = 16'b0000000000000000;
    assign weights1[7][400] = 16'b0000000000001001;
    assign weights1[7][401] = 16'b0000000000000111;
    assign weights1[7][402] = 16'b0000000000000110;
    assign weights1[7][403] = 16'b0000000000010110;
    assign weights1[7][404] = 16'b0000000000011111;
    assign weights1[7][405] = 16'b0000000000000010;
    assign weights1[7][406] = 16'b1111111111010111;
    assign weights1[7][407] = 16'b1111111110001100;
    assign weights1[7][408] = 16'b1111111101001010;
    assign weights1[7][409] = 16'b1111111101001111;
    assign weights1[7][410] = 16'b1111111101000000;
    assign weights1[7][411] = 16'b1111111101110101;
    assign weights1[7][412] = 16'b1111111101101100;
    assign weights1[7][413] = 16'b1111111110011100;
    assign weights1[7][414] = 16'b1111111110100100;
    assign weights1[7][415] = 16'b1111111110101011;
    assign weights1[7][416] = 16'b1111111110110000;
    assign weights1[7][417] = 16'b1111111111001100;
    assign weights1[7][418] = 16'b1111111110111110;
    assign weights1[7][419] = 16'b1111111110111010;
    assign weights1[7][420] = 16'b0000000000001001;
    assign weights1[7][421] = 16'b0000000000010111;
    assign weights1[7][422] = 16'b0000000000010001;
    assign weights1[7][423] = 16'b1111111111111100;
    assign weights1[7][424] = 16'b1111111111111110;
    assign weights1[7][425] = 16'b1111111111111000;
    assign weights1[7][426] = 16'b0000000000001010;
    assign weights1[7][427] = 16'b0000000000001000;
    assign weights1[7][428] = 16'b0000000000000111;
    assign weights1[7][429] = 16'b0000000000000011;
    assign weights1[7][430] = 16'b0000000000001111;
    assign weights1[7][431] = 16'b0000000000011000;
    assign weights1[7][432] = 16'b0000000000000110;
    assign weights1[7][433] = 16'b0000000000010100;
    assign weights1[7][434] = 16'b0000000000101011;
    assign weights1[7][435] = 16'b1111111111100100;
    assign weights1[7][436] = 16'b1111111110011011;
    assign weights1[7][437] = 16'b1111111101101000;
    assign weights1[7][438] = 16'b1111111100101110;
    assign weights1[7][439] = 16'b1111111100010010;
    assign weights1[7][440] = 16'b1111111100111001;
    assign weights1[7][441] = 16'b1111111101110100;
    assign weights1[7][442] = 16'b1111111101100110;
    assign weights1[7][443] = 16'b1111111110100000;
    assign weights1[7][444] = 16'b1111111110100111;
    assign weights1[7][445] = 16'b1111111110110001;
    assign weights1[7][446] = 16'b1111111111000001;
    assign weights1[7][447] = 16'b1111111110101011;
    assign weights1[7][448] = 16'b0000000000001001;
    assign weights1[7][449] = 16'b0000000000001001;
    assign weights1[7][450] = 16'b0000000000001100;
    assign weights1[7][451] = 16'b1111111111111101;
    assign weights1[7][452] = 16'b0000000000000111;
    assign weights1[7][453] = 16'b1111111111101110;
    assign weights1[7][454] = 16'b1111111111111111;
    assign weights1[7][455] = 16'b0000000000001101;
    assign weights1[7][456] = 16'b0000000000001111;
    assign weights1[7][457] = 16'b0000000000000110;
    assign weights1[7][458] = 16'b1111111111110101;
    assign weights1[7][459] = 16'b1111111111111000;
    assign weights1[7][460] = 16'b0000000000010001;
    assign weights1[7][461] = 16'b0000000000001011;
    assign weights1[7][462] = 16'b0000000000001011;
    assign weights1[7][463] = 16'b0000000000001110;
    assign weights1[7][464] = 16'b1111111111111111;
    assign weights1[7][465] = 16'b1111111111011011;
    assign weights1[7][466] = 16'b1111111110011100;
    assign weights1[7][467] = 16'b1111111101001011;
    assign weights1[7][468] = 16'b1111111100110101;
    assign weights1[7][469] = 16'b1111111101100000;
    assign weights1[7][470] = 16'b1111111101111101;
    assign weights1[7][471] = 16'b1111111110010101;
    assign weights1[7][472] = 16'b1111111110110001;
    assign weights1[7][473] = 16'b1111111110110000;
    assign weights1[7][474] = 16'b1111111110111011;
    assign weights1[7][475] = 16'b1111111110110111;
    assign weights1[7][476] = 16'b0000000000000011;
    assign weights1[7][477] = 16'b1111111111111100;
    assign weights1[7][478] = 16'b0000000000000111;
    assign weights1[7][479] = 16'b0000000000001100;
    assign weights1[7][480] = 16'b0000000000001001;
    assign weights1[7][481] = 16'b0000000000001110;
    assign weights1[7][482] = 16'b1111111111110101;
    assign weights1[7][483] = 16'b0000000000000010;
    assign weights1[7][484] = 16'b1111111111111001;
    assign weights1[7][485] = 16'b0000000000000001;
    assign weights1[7][486] = 16'b1111111111111110;
    assign weights1[7][487] = 16'b0000000000001000;
    assign weights1[7][488] = 16'b1111111111110111;
    assign weights1[7][489] = 16'b1111111111111010;
    assign weights1[7][490] = 16'b0000000000010000;
    assign weights1[7][491] = 16'b0000000000011010;
    assign weights1[7][492] = 16'b0000000000001010;
    assign weights1[7][493] = 16'b0000000000010101;
    assign weights1[7][494] = 16'b0000000000100001;
    assign weights1[7][495] = 16'b1111111111000010;
    assign weights1[7][496] = 16'b1111111101101000;
    assign weights1[7][497] = 16'b1111111101110001;
    assign weights1[7][498] = 16'b1111111110000110;
    assign weights1[7][499] = 16'b1111111110010001;
    assign weights1[7][500] = 16'b1111111110011110;
    assign weights1[7][501] = 16'b1111111110111001;
    assign weights1[7][502] = 16'b1111111111000110;
    assign weights1[7][503] = 16'b1111111111001000;
    assign weights1[7][504] = 16'b1111111111111111;
    assign weights1[7][505] = 16'b0000000000000100;
    assign weights1[7][506] = 16'b0000000000001000;
    assign weights1[7][507] = 16'b0000000000010011;
    assign weights1[7][508] = 16'b0000000000001100;
    assign weights1[7][509] = 16'b1111111111111111;
    assign weights1[7][510] = 16'b0000000000000001;
    assign weights1[7][511] = 16'b1111111111100110;
    assign weights1[7][512] = 16'b0000000000000000;
    assign weights1[7][513] = 16'b1111111111110010;
    assign weights1[7][514] = 16'b0000000000000000;
    assign weights1[7][515] = 16'b1111111111111011;
    assign weights1[7][516] = 16'b0000000000010010;
    assign weights1[7][517] = 16'b1111111111111010;
    assign weights1[7][518] = 16'b0000000000010001;
    assign weights1[7][519] = 16'b0000000000010101;
    assign weights1[7][520] = 16'b0000000000011011;
    assign weights1[7][521] = 16'b0000000000001101;
    assign weights1[7][522] = 16'b0000000000100011;
    assign weights1[7][523] = 16'b0000000000010011;
    assign weights1[7][524] = 16'b1111111111001100;
    assign weights1[7][525] = 16'b1111111110001010;
    assign weights1[7][526] = 16'b1111111110000100;
    assign weights1[7][527] = 16'b1111111110011000;
    assign weights1[7][528] = 16'b1111111110101110;
    assign weights1[7][529] = 16'b1111111110111100;
    assign weights1[7][530] = 16'b1111111111001000;
    assign weights1[7][531] = 16'b1111111111000111;
    assign weights1[7][532] = 16'b1111111111110010;
    assign weights1[7][533] = 16'b0000000000010000;
    assign weights1[7][534] = 16'b1111111111111111;
    assign weights1[7][535] = 16'b0000000000000100;
    assign weights1[7][536] = 16'b1111111111111000;
    assign weights1[7][537] = 16'b0000000000010010;
    assign weights1[7][538] = 16'b0000000000000010;
    assign weights1[7][539] = 16'b0000000000010100;
    assign weights1[7][540] = 16'b1111111111111110;
    assign weights1[7][541] = 16'b0000000000000011;
    assign weights1[7][542] = 16'b1111111111111110;
    assign weights1[7][543] = 16'b1111111111101111;
    assign weights1[7][544] = 16'b0000000000000000;
    assign weights1[7][545] = 16'b0000000000001001;
    assign weights1[7][546] = 16'b0000000000000111;
    assign weights1[7][547] = 16'b0000000000001110;
    assign weights1[7][548] = 16'b0000000000011001;
    assign weights1[7][549] = 16'b0000000000001111;
    assign weights1[7][550] = 16'b0000000000100101;
    assign weights1[7][551] = 16'b0000000000101110;
    assign weights1[7][552] = 16'b1111111111111001;
    assign weights1[7][553] = 16'b1111111111000110;
    assign weights1[7][554] = 16'b1111111110100101;
    assign weights1[7][555] = 16'b1111111110100010;
    assign weights1[7][556] = 16'b1111111110110011;
    assign weights1[7][557] = 16'b1111111110111101;
    assign weights1[7][558] = 16'b1111111111001011;
    assign weights1[7][559] = 16'b1111111111010001;
    assign weights1[7][560] = 16'b1111111111111110;
    assign weights1[7][561] = 16'b0000000000001001;
    assign weights1[7][562] = 16'b0000000000000110;
    assign weights1[7][563] = 16'b1111111111111110;
    assign weights1[7][564] = 16'b1111111111110001;
    assign weights1[7][565] = 16'b1111111111111001;
    assign weights1[7][566] = 16'b0000000000001000;
    assign weights1[7][567] = 16'b1111111111111100;
    assign weights1[7][568] = 16'b0000000000000001;
    assign weights1[7][569] = 16'b1111111111110101;
    assign weights1[7][570] = 16'b1111111111111110;
    assign weights1[7][571] = 16'b0000000000000101;
    assign weights1[7][572] = 16'b0000000000000110;
    assign weights1[7][573] = 16'b0000000000010000;
    assign weights1[7][574] = 16'b0000000000001011;
    assign weights1[7][575] = 16'b0000000000001000;
    assign weights1[7][576] = 16'b0000000000101000;
    assign weights1[7][577] = 16'b0000000000000101;
    assign weights1[7][578] = 16'b0000000000010011;
    assign weights1[7][579] = 16'b0000000000101000;
    assign weights1[7][580] = 16'b0000000000001110;
    assign weights1[7][581] = 16'b1111111111100110;
    assign weights1[7][582] = 16'b1111111110111110;
    assign weights1[7][583] = 16'b1111111110111010;
    assign weights1[7][584] = 16'b1111111110111110;
    assign weights1[7][585] = 16'b1111111111001111;
    assign weights1[7][586] = 16'b1111111111001111;
    assign weights1[7][587] = 16'b1111111111010010;
    assign weights1[7][588] = 16'b1111111111111111;
    assign weights1[7][589] = 16'b1111111111111110;
    assign weights1[7][590] = 16'b0000000000001001;
    assign weights1[7][591] = 16'b0000000000000110;
    assign weights1[7][592] = 16'b1111111111111100;
    assign weights1[7][593] = 16'b1111111111110111;
    assign weights1[7][594] = 16'b0000000000001010;
    assign weights1[7][595] = 16'b0000000000001010;
    assign weights1[7][596] = 16'b0000000000000100;
    assign weights1[7][597] = 16'b1111111111111101;
    assign weights1[7][598] = 16'b1111111111111111;
    assign weights1[7][599] = 16'b0000000000000000;
    assign weights1[7][600] = 16'b1111111111101100;
    assign weights1[7][601] = 16'b1111111111111110;
    assign weights1[7][602] = 16'b1111111111111101;
    assign weights1[7][603] = 16'b0000000000001010;
    assign weights1[7][604] = 16'b0000000000011001;
    assign weights1[7][605] = 16'b0000000000011100;
    assign weights1[7][606] = 16'b0000000000000100;
    assign weights1[7][607] = 16'b0000000000010110;
    assign weights1[7][608] = 16'b0000000000000100;
    assign weights1[7][609] = 16'b1111111111110110;
    assign weights1[7][610] = 16'b1111111111100011;
    assign weights1[7][611] = 16'b1111111111001010;
    assign weights1[7][612] = 16'b1111111111001111;
    assign weights1[7][613] = 16'b1111111111010101;
    assign weights1[7][614] = 16'b1111111111010110;
    assign weights1[7][615] = 16'b1111111111011100;
    assign weights1[7][616] = 16'b1111111111111111;
    assign weights1[7][617] = 16'b0000000000000010;
    assign weights1[7][618] = 16'b0000000000000101;
    assign weights1[7][619] = 16'b0000000000000100;
    assign weights1[7][620] = 16'b0000000000001000;
    assign weights1[7][621] = 16'b0000000000001011;
    assign weights1[7][622] = 16'b1111111111111111;
    assign weights1[7][623] = 16'b0000000000001111;
    assign weights1[7][624] = 16'b0000000000000011;
    assign weights1[7][625] = 16'b0000000000001000;
    assign weights1[7][626] = 16'b0000000000001000;
    assign weights1[7][627] = 16'b0000000000000101;
    assign weights1[7][628] = 16'b0000000000000111;
    assign weights1[7][629] = 16'b0000000000000011;
    assign weights1[7][630] = 16'b0000000000000111;
    assign weights1[7][631] = 16'b1111111111110011;
    assign weights1[7][632] = 16'b1111111111111111;
    assign weights1[7][633] = 16'b0000000000011110;
    assign weights1[7][634] = 16'b0000000000100000;
    assign weights1[7][635] = 16'b0000000000100011;
    assign weights1[7][636] = 16'b0000000000010001;
    assign weights1[7][637] = 16'b0000000000011000;
    assign weights1[7][638] = 16'b1111111111100111;
    assign weights1[7][639] = 16'b1111111111001100;
    assign weights1[7][640] = 16'b1111111111011010;
    assign weights1[7][641] = 16'b1111111111010011;
    assign weights1[7][642] = 16'b1111111111100001;
    assign weights1[7][643] = 16'b1111111111100011;
    assign weights1[7][644] = 16'b0000000000000101;
    assign weights1[7][645] = 16'b0000000000001011;
    assign weights1[7][646] = 16'b0000000000001100;
    assign weights1[7][647] = 16'b0000000000011000;
    assign weights1[7][648] = 16'b0000000000000100;
    assign weights1[7][649] = 16'b0000000000000110;
    assign weights1[7][650] = 16'b0000000000001110;
    assign weights1[7][651] = 16'b0000000000011000;
    assign weights1[7][652] = 16'b0000000000001010;
    assign weights1[7][653] = 16'b0000000000001000;
    assign weights1[7][654] = 16'b0000000000001001;
    assign weights1[7][655] = 16'b0000000000010100;
    assign weights1[7][656] = 16'b0000000000010110;
    assign weights1[7][657] = 16'b0000000000000000;
    assign weights1[7][658] = 16'b1111111111111111;
    assign weights1[7][659] = 16'b0000000000010001;
    assign weights1[7][660] = 16'b0000000000001111;
    assign weights1[7][661] = 16'b0000000000000011;
    assign weights1[7][662] = 16'b0000000000010111;
    assign weights1[7][663] = 16'b0000000000100111;
    assign weights1[7][664] = 16'b0000000000100101;
    assign weights1[7][665] = 16'b1111111111111100;
    assign weights1[7][666] = 16'b1111111111100101;
    assign weights1[7][667] = 16'b1111111111011000;
    assign weights1[7][668] = 16'b1111111111001111;
    assign weights1[7][669] = 16'b1111111111011011;
    assign weights1[7][670] = 16'b1111111111100100;
    assign weights1[7][671] = 16'b1111111111101110;
    assign weights1[7][672] = 16'b1111111111111011;
    assign weights1[7][673] = 16'b1111111111111111;
    assign weights1[7][674] = 16'b1111111111111110;
    assign weights1[7][675] = 16'b0000000000010000;
    assign weights1[7][676] = 16'b0000000000011000;
    assign weights1[7][677] = 16'b1111111111111110;
    assign weights1[7][678] = 16'b1111111111111001;
    assign weights1[7][679] = 16'b1111111111111110;
    assign weights1[7][680] = 16'b1111111111111110;
    assign weights1[7][681] = 16'b0000000000001111;
    assign weights1[7][682] = 16'b0000000000001011;
    assign weights1[7][683] = 16'b0000000000001000;
    assign weights1[7][684] = 16'b0000000000010000;
    assign weights1[7][685] = 16'b0000000000011011;
    assign weights1[7][686] = 16'b0000000000011111;
    assign weights1[7][687] = 16'b0000000000000111;
    assign weights1[7][688] = 16'b0000000000011001;
    assign weights1[7][689] = 16'b0000000000010010;
    assign weights1[7][690] = 16'b0000000000100111;
    assign weights1[7][691] = 16'b0000000000100110;
    assign weights1[7][692] = 16'b0000000000011001;
    assign weights1[7][693] = 16'b1111111111111010;
    assign weights1[7][694] = 16'b1111111111101110;
    assign weights1[7][695] = 16'b1111111111011001;
    assign weights1[7][696] = 16'b1111111111011001;
    assign weights1[7][697] = 16'b1111111111100010;
    assign weights1[7][698] = 16'b1111111111110000;
    assign weights1[7][699] = 16'b1111111111111001;
    assign weights1[7][700] = 16'b0000000000000011;
    assign weights1[7][701] = 16'b1111111111111011;
    assign weights1[7][702] = 16'b1111111111110101;
    assign weights1[7][703] = 16'b0000000000010101;
    assign weights1[7][704] = 16'b0000000000001011;
    assign weights1[7][705] = 16'b0000000000000011;
    assign weights1[7][706] = 16'b0000000000000100;
    assign weights1[7][707] = 16'b0000000000001001;
    assign weights1[7][708] = 16'b0000000000000001;
    assign weights1[7][709] = 16'b0000000000001110;
    assign weights1[7][710] = 16'b0000000000000011;
    assign weights1[7][711] = 16'b0000000000010010;
    assign weights1[7][712] = 16'b0000000000000001;
    assign weights1[7][713] = 16'b0000000000000011;
    assign weights1[7][714] = 16'b0000000000000100;
    assign weights1[7][715] = 16'b0000000000010010;
    assign weights1[7][716] = 16'b0000000000000010;
    assign weights1[7][717] = 16'b0000000000001000;
    assign weights1[7][718] = 16'b0000000000010010;
    assign weights1[7][719] = 16'b0000000000100010;
    assign weights1[7][720] = 16'b0000000000010000;
    assign weights1[7][721] = 16'b1111111111111101;
    assign weights1[7][722] = 16'b1111111111110011;
    assign weights1[7][723] = 16'b1111111111101011;
    assign weights1[7][724] = 16'b1111111111100110;
    assign weights1[7][725] = 16'b1111111111110110;
    assign weights1[7][726] = 16'b1111111111111101;
    assign weights1[7][727] = 16'b1111111111111101;
    assign weights1[7][728] = 16'b0000000000000000;
    assign weights1[7][729] = 16'b0000000000000001;
    assign weights1[7][730] = 16'b0000000000000010;
    assign weights1[7][731] = 16'b0000000000000110;
    assign weights1[7][732] = 16'b0000000000000100;
    assign weights1[7][733] = 16'b0000000000001000;
    assign weights1[7][734] = 16'b1111111111110101;
    assign weights1[7][735] = 16'b0000000000000011;
    assign weights1[7][736] = 16'b1111111111111100;
    assign weights1[7][737] = 16'b0000000000000000;
    assign weights1[7][738] = 16'b0000000000000111;
    assign weights1[7][739] = 16'b1111111111111100;
    assign weights1[7][740] = 16'b0000000000001000;
    assign weights1[7][741] = 16'b0000000000010101;
    assign weights1[7][742] = 16'b1111111111111100;
    assign weights1[7][743] = 16'b0000000000011111;
    assign weights1[7][744] = 16'b0000000000001110;
    assign weights1[7][745] = 16'b0000000000100110;
    assign weights1[7][746] = 16'b0000000000010010;
    assign weights1[7][747] = 16'b0000000000001001;
    assign weights1[7][748] = 16'b0000000000010011;
    assign weights1[7][749] = 16'b1111111111111101;
    assign weights1[7][750] = 16'b0000000000000100;
    assign weights1[7][751] = 16'b1111111111110110;
    assign weights1[7][752] = 16'b1111111111111010;
    assign weights1[7][753] = 16'b1111111111111110;
    assign weights1[7][754] = 16'b1111111111111110;
    assign weights1[7][755] = 16'b1111111111111111;
    assign weights1[7][756] = 16'b0000000000000010;
    assign weights1[7][757] = 16'b0000000000001011;
    assign weights1[7][758] = 16'b0000000000001111;
    assign weights1[7][759] = 16'b0000000000001110;
    assign weights1[7][760] = 16'b0000000000001011;
    assign weights1[7][761] = 16'b0000000000001001;
    assign weights1[7][762] = 16'b0000000000001101;
    assign weights1[7][763] = 16'b0000000000011100;
    assign weights1[7][764] = 16'b0000000000011100;
    assign weights1[7][765] = 16'b0000000000010001;
    assign weights1[7][766] = 16'b0000000000101001;
    assign weights1[7][767] = 16'b0000000000101101;
    assign weights1[7][768] = 16'b0000000000101000;
    assign weights1[7][769] = 16'b0000000000011010;
    assign weights1[7][770] = 16'b0000000000100100;
    assign weights1[7][771] = 16'b0000000000100100;
    assign weights1[7][772] = 16'b0000000000110001;
    assign weights1[7][773] = 16'b0000000000011011;
    assign weights1[7][774] = 16'b0000000000010001;
    assign weights1[7][775] = 16'b0000000000000110;
    assign weights1[7][776] = 16'b0000000000010100;
    assign weights1[7][777] = 16'b0000000000001011;
    assign weights1[7][778] = 16'b1111111111111101;
    assign weights1[7][779] = 16'b1111111111111010;
    assign weights1[7][780] = 16'b0000000000000000;
    assign weights1[7][781] = 16'b0000000000000000;
    assign weights1[7][782] = 16'b1111111111111110;
    assign weights1[7][783] = 16'b0000000000000000;
    assign weights1[8][0] = 16'b0000000000000000;
    assign weights1[8][1] = 16'b1111111111111110;
    assign weights1[8][2] = 16'b1111111111111110;
    assign weights1[8][3] = 16'b1111111111111110;
    assign weights1[8][4] = 16'b1111111111111011;
    assign weights1[8][5] = 16'b1111111111111100;
    assign weights1[8][6] = 16'b0000000000000001;
    assign weights1[8][7] = 16'b0000000000000101;
    assign weights1[8][8] = 16'b0000000000000111;
    assign weights1[8][9] = 16'b0000000000001001;
    assign weights1[8][10] = 16'b0000000000010010;
    assign weights1[8][11] = 16'b0000000000000010;
    assign weights1[8][12] = 16'b0000000000001010;
    assign weights1[8][13] = 16'b0000000000010000;
    assign weights1[8][14] = 16'b0000000000011110;
    assign weights1[8][15] = 16'b0000000000010011;
    assign weights1[8][16] = 16'b0000000000001011;
    assign weights1[8][17] = 16'b0000000000010010;
    assign weights1[8][18] = 16'b0000000000001010;
    assign weights1[8][19] = 16'b0000000000001010;
    assign weights1[8][20] = 16'b0000000000000000;
    assign weights1[8][21] = 16'b0000000000000000;
    assign weights1[8][22] = 16'b1111111111111111;
    assign weights1[8][23] = 16'b0000000000000001;
    assign weights1[8][24] = 16'b0000000000000001;
    assign weights1[8][25] = 16'b1111111111111111;
    assign weights1[8][26] = 16'b0000000000000000;
    assign weights1[8][27] = 16'b0000000000000011;
    assign weights1[8][28] = 16'b1111111111111111;
    assign weights1[8][29] = 16'b1111111111111110;
    assign weights1[8][30] = 16'b1111111111111100;
    assign weights1[8][31] = 16'b1111111111111000;
    assign weights1[8][32] = 16'b1111111111110110;
    assign weights1[8][33] = 16'b1111111111110100;
    assign weights1[8][34] = 16'b1111111111111000;
    assign weights1[8][35] = 16'b1111111111111010;
    assign weights1[8][36] = 16'b0000000000000101;
    assign weights1[8][37] = 16'b0000000000000100;
    assign weights1[8][38] = 16'b0000000000001011;
    assign weights1[8][39] = 16'b0000000000010110;
    assign weights1[8][40] = 16'b0000000000100000;
    assign weights1[8][41] = 16'b0000000000010101;
    assign weights1[8][42] = 16'b0000000000001011;
    assign weights1[8][43] = 16'b0000000000001100;
    assign weights1[8][44] = 16'b0000000000010101;
    assign weights1[8][45] = 16'b0000000000001110;
    assign weights1[8][46] = 16'b0000000000010111;
    assign weights1[8][47] = 16'b0000000000001000;
    assign weights1[8][48] = 16'b0000000000000110;
    assign weights1[8][49] = 16'b0000000000001010;
    assign weights1[8][50] = 16'b0000000000010111;
    assign weights1[8][51] = 16'b0000000000001101;
    assign weights1[8][52] = 16'b0000000000001101;
    assign weights1[8][53] = 16'b0000000000001101;
    assign weights1[8][54] = 16'b0000000000000111;
    assign weights1[8][55] = 16'b0000000000000010;
    assign weights1[8][56] = 16'b1111111111111111;
    assign weights1[8][57] = 16'b1111111111111100;
    assign weights1[8][58] = 16'b1111111111111010;
    assign weights1[8][59] = 16'b1111111111110111;
    assign weights1[8][60] = 16'b1111111111110001;
    assign weights1[8][61] = 16'b1111111111101111;
    assign weights1[8][62] = 16'b1111111111110010;
    assign weights1[8][63] = 16'b0000000000000010;
    assign weights1[8][64] = 16'b1111111111111010;
    assign weights1[8][65] = 16'b0000000000000000;
    assign weights1[8][66] = 16'b1111111111111111;
    assign weights1[8][67] = 16'b0000000000001010;
    assign weights1[8][68] = 16'b0000000000000001;
    assign weights1[8][69] = 16'b0000000000000001;
    assign weights1[8][70] = 16'b0000000000000100;
    assign weights1[8][71] = 16'b1111111111111001;
    assign weights1[8][72] = 16'b0000000000010000;
    assign weights1[8][73] = 16'b0000000000001001;
    assign weights1[8][74] = 16'b0000000000000010;
    assign weights1[8][75] = 16'b0000000000001110;
    assign weights1[8][76] = 16'b0000000000000110;
    assign weights1[8][77] = 16'b0000000000010000;
    assign weights1[8][78] = 16'b0000000000011010;
    assign weights1[8][79] = 16'b1111111111111111;
    assign weights1[8][80] = 16'b0000000000000101;
    assign weights1[8][81] = 16'b0000000000001110;
    assign weights1[8][82] = 16'b0000000000001010;
    assign weights1[8][83] = 16'b0000000000001100;
    assign weights1[8][84] = 16'b1111111111111111;
    assign weights1[8][85] = 16'b1111111111111111;
    assign weights1[8][86] = 16'b1111111111111011;
    assign weights1[8][87] = 16'b1111111111110001;
    assign weights1[8][88] = 16'b1111111111101011;
    assign weights1[8][89] = 16'b1111111111110000;
    assign weights1[8][90] = 16'b1111111111110111;
    assign weights1[8][91] = 16'b1111111111111111;
    assign weights1[8][92] = 16'b0000000000001100;
    assign weights1[8][93] = 16'b1111111111110011;
    assign weights1[8][94] = 16'b0000000000001011;
    assign weights1[8][95] = 16'b1111111111111000;
    assign weights1[8][96] = 16'b1111111111111111;
    assign weights1[8][97] = 16'b0000000000001001;
    assign weights1[8][98] = 16'b1111111111110001;
    assign weights1[8][99] = 16'b1111111111101010;
    assign weights1[8][100] = 16'b1111111111111011;
    assign weights1[8][101] = 16'b1111111111111001;
    assign weights1[8][102] = 16'b1111111111111101;
    assign weights1[8][103] = 16'b0000000000000111;
    assign weights1[8][104] = 16'b0000000000001001;
    assign weights1[8][105] = 16'b0000000000010001;
    assign weights1[8][106] = 16'b0000000000010110;
    assign weights1[8][107] = 16'b0000000000010101;
    assign weights1[8][108] = 16'b0000000000010111;
    assign weights1[8][109] = 16'b0000000000001010;
    assign weights1[8][110] = 16'b0000000000010000;
    assign weights1[8][111] = 16'b0000000000010000;
    assign weights1[8][112] = 16'b1111111111111011;
    assign weights1[8][113] = 16'b1111111111111001;
    assign weights1[8][114] = 16'b1111111111111000;
    assign weights1[8][115] = 16'b1111111111110010;
    assign weights1[8][116] = 16'b1111111111101100;
    assign weights1[8][117] = 16'b1111111111101001;
    assign weights1[8][118] = 16'b1111111111110110;
    assign weights1[8][119] = 16'b0000000000000011;
    assign weights1[8][120] = 16'b1111111111110010;
    assign weights1[8][121] = 16'b0000000000010010;
    assign weights1[8][122] = 16'b0000000000010110;
    assign weights1[8][123] = 16'b1111111111110101;
    assign weights1[8][124] = 16'b0000000000001111;
    assign weights1[8][125] = 16'b0000000000000110;
    assign weights1[8][126] = 16'b1111111111111000;
    assign weights1[8][127] = 16'b0000000000010001;
    assign weights1[8][128] = 16'b0000000000001100;
    assign weights1[8][129] = 16'b1111111111111010;
    assign weights1[8][130] = 16'b1111111111101111;
    assign weights1[8][131] = 16'b1111111111111011;
    assign weights1[8][132] = 16'b0000000000001101;
    assign weights1[8][133] = 16'b1111111111111001;
    assign weights1[8][134] = 16'b1111111111111100;
    assign weights1[8][135] = 16'b0000000000000111;
    assign weights1[8][136] = 16'b1111111111111000;
    assign weights1[8][137] = 16'b0000000000001000;
    assign weights1[8][138] = 16'b0000000000010000;
    assign weights1[8][139] = 16'b0000000000001011;
    assign weights1[8][140] = 16'b1111111111111100;
    assign weights1[8][141] = 16'b1111111111111000;
    assign weights1[8][142] = 16'b1111111111111010;
    assign weights1[8][143] = 16'b1111111111111100;
    assign weights1[8][144] = 16'b1111111111110111;
    assign weights1[8][145] = 16'b1111111111100101;
    assign weights1[8][146] = 16'b1111111111101101;
    assign weights1[8][147] = 16'b0000000000000101;
    assign weights1[8][148] = 16'b1111111111101110;
    assign weights1[8][149] = 16'b0000000000001001;
    assign weights1[8][150] = 16'b0000000000000110;
    assign weights1[8][151] = 16'b0000000000000100;
    assign weights1[8][152] = 16'b0000000000001010;
    assign weights1[8][153] = 16'b1111111111101011;
    assign weights1[8][154] = 16'b0000000000001110;
    assign weights1[8][155] = 16'b1111111111111001;
    assign weights1[8][156] = 16'b0000000000011101;
    assign weights1[8][157] = 16'b0000000000001110;
    assign weights1[8][158] = 16'b0000000000011101;
    assign weights1[8][159] = 16'b0000000000001001;
    assign weights1[8][160] = 16'b0000000000010111;
    assign weights1[8][161] = 16'b0000000000010110;
    assign weights1[8][162] = 16'b0000000000001010;
    assign weights1[8][163] = 16'b1111111111110110;
    assign weights1[8][164] = 16'b0000000000000111;
    assign weights1[8][165] = 16'b0000000000100001;
    assign weights1[8][166] = 16'b0000000000001110;
    assign weights1[8][167] = 16'b0000000000010001;
    assign weights1[8][168] = 16'b1111111111111001;
    assign weights1[8][169] = 16'b1111111111110000;
    assign weights1[8][170] = 16'b1111111111110001;
    assign weights1[8][171] = 16'b1111111111110110;
    assign weights1[8][172] = 16'b1111111111111000;
    assign weights1[8][173] = 16'b1111111111101000;
    assign weights1[8][174] = 16'b1111111111101010;
    assign weights1[8][175] = 16'b1111111111100101;
    assign weights1[8][176] = 16'b1111111111110001;
    assign weights1[8][177] = 16'b0000000000011001;
    assign weights1[8][178] = 16'b1111111111101111;
    assign weights1[8][179] = 16'b1111111111111110;
    assign weights1[8][180] = 16'b0000000000001110;
    assign weights1[8][181] = 16'b0000000000000010;
    assign weights1[8][182] = 16'b1111111111111100;
    assign weights1[8][183] = 16'b0000000000010000;
    assign weights1[8][184] = 16'b1111111111111001;
    assign weights1[8][185] = 16'b1111111111111010;
    assign weights1[8][186] = 16'b0000000000010111;
    assign weights1[8][187] = 16'b0000000000001010;
    assign weights1[8][188] = 16'b0000000000000000;
    assign weights1[8][189] = 16'b0000000000011000;
    assign weights1[8][190] = 16'b1111111111110000;
    assign weights1[8][191] = 16'b0000000000000110;
    assign weights1[8][192] = 16'b0000000000011111;
    assign weights1[8][193] = 16'b0000000000011001;
    assign weights1[8][194] = 16'b0000000000010110;
    assign weights1[8][195] = 16'b1111111111111111;
    assign weights1[8][196] = 16'b1111111111110101;
    assign weights1[8][197] = 16'b1111111111110100;
    assign weights1[8][198] = 16'b1111111111111111;
    assign weights1[8][199] = 16'b1111111111111010;
    assign weights1[8][200] = 16'b0000000000000011;
    assign weights1[8][201] = 16'b1111111111101101;
    assign weights1[8][202] = 16'b1111111111100101;
    assign weights1[8][203] = 16'b1111111111110011;
    assign weights1[8][204] = 16'b0000000000000000;
    assign weights1[8][205] = 16'b1111111111111000;
    assign weights1[8][206] = 16'b0000000000001111;
    assign weights1[8][207] = 16'b0000000000000110;
    assign weights1[8][208] = 16'b1111111111111100;
    assign weights1[8][209] = 16'b0000000000001000;
    assign weights1[8][210] = 16'b1111111111110001;
    assign weights1[8][211] = 16'b0000000000000001;
    assign weights1[8][212] = 16'b0000000000001001;
    assign weights1[8][213] = 16'b0000000000000110;
    assign weights1[8][214] = 16'b0000000000000110;
    assign weights1[8][215] = 16'b1111111111101110;
    assign weights1[8][216] = 16'b0000000000000011;
    assign weights1[8][217] = 16'b1111111111101101;
    assign weights1[8][218] = 16'b0000000000100000;
    assign weights1[8][219] = 16'b0000000000001110;
    assign weights1[8][220] = 16'b0000000000000000;
    assign weights1[8][221] = 16'b0000000000000110;
    assign weights1[8][222] = 16'b0000000000001100;
    assign weights1[8][223] = 16'b0000000000000011;
    assign weights1[8][224] = 16'b1111111111111010;
    assign weights1[8][225] = 16'b1111111111111011;
    assign weights1[8][226] = 16'b1111111111111110;
    assign weights1[8][227] = 16'b1111111111110011;
    assign weights1[8][228] = 16'b1111111111111111;
    assign weights1[8][229] = 16'b1111111111100110;
    assign weights1[8][230] = 16'b0000000000000010;
    assign weights1[8][231] = 16'b1111111111101000;
    assign weights1[8][232] = 16'b1111111111101111;
    assign weights1[8][233] = 16'b1111111111110010;
    assign weights1[8][234] = 16'b1111111111111010;
    assign weights1[8][235] = 16'b0000000000001111;
    assign weights1[8][236] = 16'b0000000000001001;
    assign weights1[8][237] = 16'b0000000000010011;
    assign weights1[8][238] = 16'b0000000000001110;
    assign weights1[8][239] = 16'b0000000000000100;
    assign weights1[8][240] = 16'b0000000000000111;
    assign weights1[8][241] = 16'b0000000000000110;
    assign weights1[8][242] = 16'b1111111111111110;
    assign weights1[8][243] = 16'b0000000000010001;
    assign weights1[8][244] = 16'b0000000000010001;
    assign weights1[8][245] = 16'b0000000000010010;
    assign weights1[8][246] = 16'b0000000000000110;
    assign weights1[8][247] = 16'b0000000000001001;
    assign weights1[8][248] = 16'b0000000000100010;
    assign weights1[8][249] = 16'b0000000000000000;
    assign weights1[8][250] = 16'b1111111111111000;
    assign weights1[8][251] = 16'b1111111111111000;
    assign weights1[8][252] = 16'b1111111111111101;
    assign weights1[8][253] = 16'b0000000000000010;
    assign weights1[8][254] = 16'b0000000000001000;
    assign weights1[8][255] = 16'b1111111111110110;
    assign weights1[8][256] = 16'b1111111111110001;
    assign weights1[8][257] = 16'b0000000000000110;
    assign weights1[8][258] = 16'b0000000000000010;
    assign weights1[8][259] = 16'b0000000000001000;
    assign weights1[8][260] = 16'b0000000000000010;
    assign weights1[8][261] = 16'b1111111111111001;
    assign weights1[8][262] = 16'b1111111111110110;
    assign weights1[8][263] = 16'b1111111111111110;
    assign weights1[8][264] = 16'b1111111111110111;
    assign weights1[8][265] = 16'b1111111111101110;
    assign weights1[8][266] = 16'b1111111111110011;
    assign weights1[8][267] = 16'b1111111111101111;
    assign weights1[8][268] = 16'b1111111111011110;
    assign weights1[8][269] = 16'b0000000000000101;
    assign weights1[8][270] = 16'b1111111111110000;
    assign weights1[8][271] = 16'b1111111111110111;
    assign weights1[8][272] = 16'b1111111111110111;
    assign weights1[8][273] = 16'b0000000000010000;
    assign weights1[8][274] = 16'b0000000000100010;
    assign weights1[8][275] = 16'b0000000000100101;
    assign weights1[8][276] = 16'b0000000000010011;
    assign weights1[8][277] = 16'b0000000000000001;
    assign weights1[8][278] = 16'b1111111111111000;
    assign weights1[8][279] = 16'b1111111111011010;
    assign weights1[8][280] = 16'b1111111111110100;
    assign weights1[8][281] = 16'b0000000000000101;
    assign weights1[8][282] = 16'b1111111111111100;
    assign weights1[8][283] = 16'b1111111111101110;
    assign weights1[8][284] = 16'b0000000000000111;
    assign weights1[8][285] = 16'b0000000000011011;
    assign weights1[8][286] = 16'b0000000000001010;
    assign weights1[8][287] = 16'b1111111111110011;
    assign weights1[8][288] = 16'b0000000000001101;
    assign weights1[8][289] = 16'b0000000000010001;
    assign weights1[8][290] = 16'b1111111111111010;
    assign weights1[8][291] = 16'b1111111111110011;
    assign weights1[8][292] = 16'b1111111111111101;
    assign weights1[8][293] = 16'b1111111111100110;
    assign weights1[8][294] = 16'b1111111111011011;
    assign weights1[8][295] = 16'b1111111111011100;
    assign weights1[8][296] = 16'b1111111111111101;
    assign weights1[8][297] = 16'b1111111111100011;
    assign weights1[8][298] = 16'b0000000000000111;
    assign weights1[8][299] = 16'b1111111111111011;
    assign weights1[8][300] = 16'b1111111111110001;
    assign weights1[8][301] = 16'b1111111111111110;
    assign weights1[8][302] = 16'b0000000000010101;
    assign weights1[8][303] = 16'b0000000000101100;
    assign weights1[8][304] = 16'b1111111111110011;
    assign weights1[8][305] = 16'b1111111111101111;
    assign weights1[8][306] = 16'b1111111111001100;
    assign weights1[8][307] = 16'b1111111111000010;
    assign weights1[8][308] = 16'b1111111111110011;
    assign weights1[8][309] = 16'b1111111111110111;
    assign weights1[8][310] = 16'b1111111111111000;
    assign weights1[8][311] = 16'b1111111111101110;
    assign weights1[8][312] = 16'b0000000000010111;
    assign weights1[8][313] = 16'b0000000000100010;
    assign weights1[8][314] = 16'b0000000000010110;
    assign weights1[8][315] = 16'b0000000000001100;
    assign weights1[8][316] = 16'b1111111111110000;
    assign weights1[8][317] = 16'b1111111111100011;
    assign weights1[8][318] = 16'b1111111111110010;
    assign weights1[8][319] = 16'b1111111111110000;
    assign weights1[8][320] = 16'b1111111111110110;
    assign weights1[8][321] = 16'b1111111111110010;
    assign weights1[8][322] = 16'b0000000000000110;
    assign weights1[8][323] = 16'b1111111111010011;
    assign weights1[8][324] = 16'b1111111111011001;
    assign weights1[8][325] = 16'b1111111111100000;
    assign weights1[8][326] = 16'b1111111111110111;
    assign weights1[8][327] = 16'b1111111111111101;
    assign weights1[8][328] = 16'b0000000000000010;
    assign weights1[8][329] = 16'b0000000000001100;
    assign weights1[8][330] = 16'b0000000000100010;
    assign weights1[8][331] = 16'b1111111111110111;
    assign weights1[8][332] = 16'b1111111111000010;
    assign weights1[8][333] = 16'b1111111111000101;
    assign weights1[8][334] = 16'b1111111110110110;
    assign weights1[8][335] = 16'b1111111110111100;
    assign weights1[8][336] = 16'b1111111111111100;
    assign weights1[8][337] = 16'b1111111111110010;
    assign weights1[8][338] = 16'b1111111111110010;
    assign weights1[8][339] = 16'b1111111111111101;
    assign weights1[8][340] = 16'b0000000000010001;
    assign weights1[8][341] = 16'b0000000000000101;
    assign weights1[8][342] = 16'b1111111111100001;
    assign weights1[8][343] = 16'b0000000000000001;
    assign weights1[8][344] = 16'b1111111111111011;
    assign weights1[8][345] = 16'b1111111111100001;
    assign weights1[8][346] = 16'b1111111111100111;
    assign weights1[8][347] = 16'b1111111111111010;
    assign weights1[8][348] = 16'b1111111111100101;
    assign weights1[8][349] = 16'b0000000000001101;
    assign weights1[8][350] = 16'b0000000000000010;
    assign weights1[8][351] = 16'b1111111111101000;
    assign weights1[8][352] = 16'b1111111111100001;
    assign weights1[8][353] = 16'b1111111111001101;
    assign weights1[8][354] = 16'b1111111111011101;
    assign weights1[8][355] = 16'b1111111111100100;
    assign weights1[8][356] = 16'b1111111111100100;
    assign weights1[8][357] = 16'b1111111111101001;
    assign weights1[8][358] = 16'b1111111111000010;
    assign weights1[8][359] = 16'b1111111110001101;
    assign weights1[8][360] = 16'b1111111110001000;
    assign weights1[8][361] = 16'b1111111110010111;
    assign weights1[8][362] = 16'b1111111110111000;
    assign weights1[8][363] = 16'b1111111110110101;
    assign weights1[8][364] = 16'b1111111111110010;
    assign weights1[8][365] = 16'b1111111111110001;
    assign weights1[8][366] = 16'b1111111111110001;
    assign weights1[8][367] = 16'b1111111111110100;
    assign weights1[8][368] = 16'b1111111111011000;
    assign weights1[8][369] = 16'b1111111111011010;
    assign weights1[8][370] = 16'b1111111111011111;
    assign weights1[8][371] = 16'b1111111111011001;
    assign weights1[8][372] = 16'b1111111111011001;
    assign weights1[8][373] = 16'b1111111111111010;
    assign weights1[8][374] = 16'b1111111111100001;
    assign weights1[8][375] = 16'b1111111111100110;
    assign weights1[8][376] = 16'b0000000000011111;
    assign weights1[8][377] = 16'b0000000000010111;
    assign weights1[8][378] = 16'b0000000000101111;
    assign weights1[8][379] = 16'b0000000000000001;
    assign weights1[8][380] = 16'b1111111111011000;
    assign weights1[8][381] = 16'b1111111111100101;
    assign weights1[8][382] = 16'b1111111111011000;
    assign weights1[8][383] = 16'b1111111111001101;
    assign weights1[8][384] = 16'b1111111110100010;
    assign weights1[8][385] = 16'b1111111101110000;
    assign weights1[8][386] = 16'b1111111101011010;
    assign weights1[8][387] = 16'b1111111101101010;
    assign weights1[8][388] = 16'b1111111101111001;
    assign weights1[8][389] = 16'b1111111110011111;
    assign weights1[8][390] = 16'b1111111110110000;
    assign weights1[8][391] = 16'b1111111110110111;
    assign weights1[8][392] = 16'b1111111111101101;
    assign weights1[8][393] = 16'b1111111111101101;
    assign weights1[8][394] = 16'b1111111111100001;
    assign weights1[8][395] = 16'b1111111111011100;
    assign weights1[8][396] = 16'b1111111111010100;
    assign weights1[8][397] = 16'b1111111110111110;
    assign weights1[8][398] = 16'b1111111111011011;
    assign weights1[8][399] = 16'b1111111111011000;
    assign weights1[8][400] = 16'b1111111111010111;
    assign weights1[8][401] = 16'b1111111111011101;
    assign weights1[8][402] = 16'b1111111111101111;
    assign weights1[8][403] = 16'b0000000000010011;
    assign weights1[8][404] = 16'b0000000000100101;
    assign weights1[8][405] = 16'b0000000000100100;
    assign weights1[8][406] = 16'b0000000000001101;
    assign weights1[8][407] = 16'b0000000000100011;
    assign weights1[8][408] = 16'b0000000000001000;
    assign weights1[8][409] = 16'b1111111111111000;
    assign weights1[8][410] = 16'b1111111111100110;
    assign weights1[8][411] = 16'b1111111111011100;
    assign weights1[8][412] = 16'b1111111110110000;
    assign weights1[8][413] = 16'b1111111110010011;
    assign weights1[8][414] = 16'b1111111101011001;
    assign weights1[8][415] = 16'b1111111101100100;
    assign weights1[8][416] = 16'b1111111101111011;
    assign weights1[8][417] = 16'b1111111110010101;
    assign weights1[8][418] = 16'b1111111110100101;
    assign weights1[8][419] = 16'b1111111110101111;
    assign weights1[8][420] = 16'b1111111111101111;
    assign weights1[8][421] = 16'b1111111111101001;
    assign weights1[8][422] = 16'b1111111111010110;
    assign weights1[8][423] = 16'b1111111111001100;
    assign weights1[8][424] = 16'b1111111111000110;
    assign weights1[8][425] = 16'b1111111111001101;
    assign weights1[8][426] = 16'b1111111110111101;
    assign weights1[8][427] = 16'b1111111111110011;
    assign weights1[8][428] = 16'b1111111111110000;
    assign weights1[8][429] = 16'b0000000000000000;
    assign weights1[8][430] = 16'b0000000000000100;
    assign weights1[8][431] = 16'b0000000000000010;
    assign weights1[8][432] = 16'b0000000000001111;
    assign weights1[8][433] = 16'b0000000000101000;
    assign weights1[8][434] = 16'b0000000000101010;
    assign weights1[8][435] = 16'b0000000000011100;
    assign weights1[8][436] = 16'b0000000000011011;
    assign weights1[8][437] = 16'b0000000000000000;
    assign weights1[8][438] = 16'b1111111111110110;
    assign weights1[8][439] = 16'b1111111111110100;
    assign weights1[8][440] = 16'b1111111111011101;
    assign weights1[8][441] = 16'b1111111111000010;
    assign weights1[8][442] = 16'b1111111110111111;
    assign weights1[8][443] = 16'b1111111110100000;
    assign weights1[8][444] = 16'b1111111110010100;
    assign weights1[8][445] = 16'b1111111110010011;
    assign weights1[8][446] = 16'b1111111110100101;
    assign weights1[8][447] = 16'b1111111110110000;
    assign weights1[8][448] = 16'b1111111111101110;
    assign weights1[8][449] = 16'b1111111111100110;
    assign weights1[8][450] = 16'b1111111111001110;
    assign weights1[8][451] = 16'b1111111111000011;
    assign weights1[8][452] = 16'b1111111111001001;
    assign weights1[8][453] = 16'b1111111111011011;
    assign weights1[8][454] = 16'b1111111111110101;
    assign weights1[8][455] = 16'b0000000000001010;
    assign weights1[8][456] = 16'b0000000000000011;
    assign weights1[8][457] = 16'b0000000000010010;
    assign weights1[8][458] = 16'b0000000000011101;
    assign weights1[8][459] = 16'b0000000000001010;
    assign weights1[8][460] = 16'b0000000000001110;
    assign weights1[8][461] = 16'b1111111111111111;
    assign weights1[8][462] = 16'b0000000000100100;
    assign weights1[8][463] = 16'b0000000000101001;
    assign weights1[8][464] = 16'b1111111111111101;
    assign weights1[8][465] = 16'b1111111111111100;
    assign weights1[8][466] = 16'b1111111111100110;
    assign weights1[8][467] = 16'b0000000000000000;
    assign weights1[8][468] = 16'b1111111111110010;
    assign weights1[8][469] = 16'b1111111111110011;
    assign weights1[8][470] = 16'b1111111111110010;
    assign weights1[8][471] = 16'b1111111111011110;
    assign weights1[8][472] = 16'b1111111111001010;
    assign weights1[8][473] = 16'b1111111110110010;
    assign weights1[8][474] = 16'b1111111110101101;
    assign weights1[8][475] = 16'b1111111111000100;
    assign weights1[8][476] = 16'b1111111111101111;
    assign weights1[8][477] = 16'b1111111111100101;
    assign weights1[8][478] = 16'b1111111111010011;
    assign weights1[8][479] = 16'b1111111111011010;
    assign weights1[8][480] = 16'b1111111111100101;
    assign weights1[8][481] = 16'b0000000000000001;
    assign weights1[8][482] = 16'b0000000000010010;
    assign weights1[8][483] = 16'b0000000000000110;
    assign weights1[8][484] = 16'b0000000000001110;
    assign weights1[8][485] = 16'b0000000000010011;
    assign weights1[8][486] = 16'b1111111111111101;
    assign weights1[8][487] = 16'b1111111111110101;
    assign weights1[8][488] = 16'b0000000000100001;
    assign weights1[8][489] = 16'b0000000000001010;
    assign weights1[8][490] = 16'b1111111111111101;
    assign weights1[8][491] = 16'b1111111111111111;
    assign weights1[8][492] = 16'b0000000000010011;
    assign weights1[8][493] = 16'b1111111111111000;
    assign weights1[8][494] = 16'b0000000000000111;
    assign weights1[8][495] = 16'b0000000000001011;
    assign weights1[8][496] = 16'b0000000000011100;
    assign weights1[8][497] = 16'b0000000000011011;
    assign weights1[8][498] = 16'b0000000000010111;
    assign weights1[8][499] = 16'b1111111111110011;
    assign weights1[8][500] = 16'b1111111111101111;
    assign weights1[8][501] = 16'b1111111111100000;
    assign weights1[8][502] = 16'b1111111111001100;
    assign weights1[8][503] = 16'b1111111111011100;
    assign weights1[8][504] = 16'b1111111111110010;
    assign weights1[8][505] = 16'b1111111111100010;
    assign weights1[8][506] = 16'b1111111111100010;
    assign weights1[8][507] = 16'b1111111111101111;
    assign weights1[8][508] = 16'b0000000000001101;
    assign weights1[8][509] = 16'b0000000000011001;
    assign weights1[8][510] = 16'b0000000000011101;
    assign weights1[8][511] = 16'b0000000000010100;
    assign weights1[8][512] = 16'b1111111111111101;
    assign weights1[8][513] = 16'b0000000000011110;
    assign weights1[8][514] = 16'b0000000000000110;
    assign weights1[8][515] = 16'b0000000000000110;
    assign weights1[8][516] = 16'b0000000000001111;
    assign weights1[8][517] = 16'b0000000000001100;
    assign weights1[8][518] = 16'b1111111111110011;
    assign weights1[8][519] = 16'b0000000000000110;
    assign weights1[8][520] = 16'b0000000000010110;
    assign weights1[8][521] = 16'b0000000000010010;
    assign weights1[8][522] = 16'b0000000000010001;
    assign weights1[8][523] = 16'b0000000000100010;
    assign weights1[8][524] = 16'b0000000000101001;
    assign weights1[8][525] = 16'b0000000000011000;
    assign weights1[8][526] = 16'b0000000000110000;
    assign weights1[8][527] = 16'b0000000000011100;
    assign weights1[8][528] = 16'b0000000000010010;
    assign weights1[8][529] = 16'b0000000000000100;
    assign weights1[8][530] = 16'b1111111111110000;
    assign weights1[8][531] = 16'b1111111111111011;
    assign weights1[8][532] = 16'b1111111111111011;
    assign weights1[8][533] = 16'b1111111111111100;
    assign weights1[8][534] = 16'b1111111111110111;
    assign weights1[8][535] = 16'b0000000000000101;
    assign weights1[8][536] = 16'b0000000000001011;
    assign weights1[8][537] = 16'b0000000000000011;
    assign weights1[8][538] = 16'b0000000000001001;
    assign weights1[8][539] = 16'b0000000000001011;
    assign weights1[8][540] = 16'b0000000000000001;
    assign weights1[8][541] = 16'b0000000000000101;
    assign weights1[8][542] = 16'b0000000000011001;
    assign weights1[8][543] = 16'b0000000000000000;
    assign weights1[8][544] = 16'b1111111111111101;
    assign weights1[8][545] = 16'b0000000000001010;
    assign weights1[8][546] = 16'b0000000000000001;
    assign weights1[8][547] = 16'b0000000000010110;
    assign weights1[8][548] = 16'b0000000000000010;
    assign weights1[8][549] = 16'b0000000000010110;
    assign weights1[8][550] = 16'b0000000000001001;
    assign weights1[8][551] = 16'b0000000000011101;
    assign weights1[8][552] = 16'b0000000000011101;
    assign weights1[8][553] = 16'b0000000001000001;
    assign weights1[8][554] = 16'b0000000001000110;
    assign weights1[8][555] = 16'b0000000001010101;
    assign weights1[8][556] = 16'b0000000000100001;
    assign weights1[8][557] = 16'b0000000000100110;
    assign weights1[8][558] = 16'b0000000000100011;
    assign weights1[8][559] = 16'b0000000000010101;
    assign weights1[8][560] = 16'b0000000000001011;
    assign weights1[8][561] = 16'b0000000000000111;
    assign weights1[8][562] = 16'b0000000000001100;
    assign weights1[8][563] = 16'b0000000000000011;
    assign weights1[8][564] = 16'b1111111111111101;
    assign weights1[8][565] = 16'b0000000000110101;
    assign weights1[8][566] = 16'b0000000000011010;
    assign weights1[8][567] = 16'b0000000000011101;
    assign weights1[8][568] = 16'b0000000000001100;
    assign weights1[8][569] = 16'b0000000000000010;
    assign weights1[8][570] = 16'b0000000000011010;
    assign weights1[8][571] = 16'b0000000000001010;
    assign weights1[8][572] = 16'b1111111111111010;
    assign weights1[8][573] = 16'b0000000000010011;
    assign weights1[8][574] = 16'b0000000000000001;
    assign weights1[8][575] = 16'b0000000000001001;
    assign weights1[8][576] = 16'b0000000000010011;
    assign weights1[8][577] = 16'b0000000000011011;
    assign weights1[8][578] = 16'b0000000000110110;
    assign weights1[8][579] = 16'b0000000000001110;
    assign weights1[8][580] = 16'b0000000000111001;
    assign weights1[8][581] = 16'b0000000000101110;
    assign weights1[8][582] = 16'b0000000000111000;
    assign weights1[8][583] = 16'b0000000001100001;
    assign weights1[8][584] = 16'b0000000000110110;
    assign weights1[8][585] = 16'b0000000000110111;
    assign weights1[8][586] = 16'b0000000000110100;
    assign weights1[8][587] = 16'b0000000000011010;
    assign weights1[8][588] = 16'b0000000000010001;
    assign weights1[8][589] = 16'b0000000000010101;
    assign weights1[8][590] = 16'b0000000000010010;
    assign weights1[8][591] = 16'b1111111111110110;
    assign weights1[8][592] = 16'b1111111111110111;
    assign weights1[8][593] = 16'b0000000000011011;
    assign weights1[8][594] = 16'b0000000000001010;
    assign weights1[8][595] = 16'b0000000000001001;
    assign weights1[8][596] = 16'b0000000000010001;
    assign weights1[8][597] = 16'b0000000000011000;
    assign weights1[8][598] = 16'b1111111111111010;
    assign weights1[8][599] = 16'b0000000000001011;
    assign weights1[8][600] = 16'b0000000000010100;
    assign weights1[8][601] = 16'b0000000000100111;
    assign weights1[8][602] = 16'b0000000000011100;
    assign weights1[8][603] = 16'b0000000000000111;
    assign weights1[8][604] = 16'b0000000000001110;
    assign weights1[8][605] = 16'b0000000000010111;
    assign weights1[8][606] = 16'b0000000000100110;
    assign weights1[8][607] = 16'b0000000000101101;
    assign weights1[8][608] = 16'b0000000000110100;
    assign weights1[8][609] = 16'b0000000000110011;
    assign weights1[8][610] = 16'b0000000000111000;
    assign weights1[8][611] = 16'b0000000001001100;
    assign weights1[8][612] = 16'b0000000000110111;
    assign weights1[8][613] = 16'b0000000001000110;
    assign weights1[8][614] = 16'b0000000000101110;
    assign weights1[8][615] = 16'b0000000000011100;
    assign weights1[8][616] = 16'b0000000000001101;
    assign weights1[8][617] = 16'b0000000000010001;
    assign weights1[8][618] = 16'b0000000000001010;
    assign weights1[8][619] = 16'b1111111111111011;
    assign weights1[8][620] = 16'b0000000000000111;
    assign weights1[8][621] = 16'b0000000000001101;
    assign weights1[8][622] = 16'b1111111111110111;
    assign weights1[8][623] = 16'b0000000000001100;
    assign weights1[8][624] = 16'b0000000000000010;
    assign weights1[8][625] = 16'b0000000000010100;
    assign weights1[8][626] = 16'b0000000000000010;
    assign weights1[8][627] = 16'b0000000000011111;
    assign weights1[8][628] = 16'b0000000000000110;
    assign weights1[8][629] = 16'b1111111111111110;
    assign weights1[8][630] = 16'b1111111111111101;
    assign weights1[8][631] = 16'b0000000000011001;
    assign weights1[8][632] = 16'b1111111111111000;
    assign weights1[8][633] = 16'b0000000000001110;
    assign weights1[8][634] = 16'b0000000000010101;
    assign weights1[8][635] = 16'b0000000000101010;
    assign weights1[8][636] = 16'b0000000000001111;
    assign weights1[8][637] = 16'b0000000000100100;
    assign weights1[8][638] = 16'b0000000000001111;
    assign weights1[8][639] = 16'b0000000000100010;
    assign weights1[8][640] = 16'b0000000000101111;
    assign weights1[8][641] = 16'b0000000000101110;
    assign weights1[8][642] = 16'b0000000000100010;
    assign weights1[8][643] = 16'b0000000000010100;
    assign weights1[8][644] = 16'b0000000000010001;
    assign weights1[8][645] = 16'b0000000000010110;
    assign weights1[8][646] = 16'b0000000000000111;
    assign weights1[8][647] = 16'b0000000000000010;
    assign weights1[8][648] = 16'b0000000000000111;
    assign weights1[8][649] = 16'b0000000000010101;
    assign weights1[8][650] = 16'b0000000000000001;
    assign weights1[8][651] = 16'b0000000000001100;
    assign weights1[8][652] = 16'b0000000000001100;
    assign weights1[8][653] = 16'b0000000000010000;
    assign weights1[8][654] = 16'b0000000000000110;
    assign weights1[8][655] = 16'b0000000000010111;
    assign weights1[8][656] = 16'b0000000000011000;
    assign weights1[8][657] = 16'b0000000000101011;
    assign weights1[8][658] = 16'b0000000000001010;
    assign weights1[8][659] = 16'b0000000000101001;
    assign weights1[8][660] = 16'b0000000000100000;
    assign weights1[8][661] = 16'b1111111111111110;
    assign weights1[8][662] = 16'b0000000000000010;
    assign weights1[8][663] = 16'b0000000000001001;
    assign weights1[8][664] = 16'b0000000000100111;
    assign weights1[8][665] = 16'b1111111111101011;
    assign weights1[8][666] = 16'b0000000000001100;
    assign weights1[8][667] = 16'b0000000000010000;
    assign weights1[8][668] = 16'b0000000000010010;
    assign weights1[8][669] = 16'b0000000000011010;
    assign weights1[8][670] = 16'b0000000000010001;
    assign weights1[8][671] = 16'b0000000000001010;
    assign weights1[8][672] = 16'b0000000000000110;
    assign weights1[8][673] = 16'b0000000000000100;
    assign weights1[8][674] = 16'b0000000000000011;
    assign weights1[8][675] = 16'b1111111111111100;
    assign weights1[8][676] = 16'b0000000000000101;
    assign weights1[8][677] = 16'b0000000000000010;
    assign weights1[8][678] = 16'b1111111111011011;
    assign weights1[8][679] = 16'b1111111111100010;
    assign weights1[8][680] = 16'b1111111111111110;
    assign weights1[8][681] = 16'b0000000000000010;
    assign weights1[8][682] = 16'b1111111111101001;
    assign weights1[8][683] = 16'b0000000000010100;
    assign weights1[8][684] = 16'b0000000000010010;
    assign weights1[8][685] = 16'b0000000000001001;
    assign weights1[8][686] = 16'b1111111111110100;
    assign weights1[8][687] = 16'b0000000000000101;
    assign weights1[8][688] = 16'b0000000000010010;
    assign weights1[8][689] = 16'b1111111111100010;
    assign weights1[8][690] = 16'b0000000000011010;
    assign weights1[8][691] = 16'b1111111111111100;
    assign weights1[8][692] = 16'b1111111111101101;
    assign weights1[8][693] = 16'b1111111111111000;
    assign weights1[8][694] = 16'b1111111111100111;
    assign weights1[8][695] = 16'b1111111111001010;
    assign weights1[8][696] = 16'b1111111111110010;
    assign weights1[8][697] = 16'b0000000000000010;
    assign weights1[8][698] = 16'b1111111111111111;
    assign weights1[8][699] = 16'b0000000000000000;
    assign weights1[8][700] = 16'b0000000000000011;
    assign weights1[8][701] = 16'b0000000000000111;
    assign weights1[8][702] = 16'b0000000000000001;
    assign weights1[8][703] = 16'b0000000000000111;
    assign weights1[8][704] = 16'b0000000000001010;
    assign weights1[8][705] = 16'b0000000000000100;
    assign weights1[8][706] = 16'b1111111111110010;
    assign weights1[8][707] = 16'b1111111111101110;
    assign weights1[8][708] = 16'b1111111111110101;
    assign weights1[8][709] = 16'b1111111111101100;
    assign weights1[8][710] = 16'b1111111111111110;
    assign weights1[8][711] = 16'b1111111111010011;
    assign weights1[8][712] = 16'b1111111111010001;
    assign weights1[8][713] = 16'b1111111111011101;
    assign weights1[8][714] = 16'b1111111111101111;
    assign weights1[8][715] = 16'b1111111111111001;
    assign weights1[8][716] = 16'b1111111111001001;
    assign weights1[8][717] = 16'b1111111111100110;
    assign weights1[8][718] = 16'b1111111111010110;
    assign weights1[8][719] = 16'b1111111111001011;
    assign weights1[8][720] = 16'b1111111111001001;
    assign weights1[8][721] = 16'b1111111110111100;
    assign weights1[8][722] = 16'b1111111110111101;
    assign weights1[8][723] = 16'b1111111111000111;
    assign weights1[8][724] = 16'b1111111111100111;
    assign weights1[8][725] = 16'b1111111111111001;
    assign weights1[8][726] = 16'b1111111111111011;
    assign weights1[8][727] = 16'b1111111111111011;
    assign weights1[8][728] = 16'b0000000000000000;
    assign weights1[8][729] = 16'b0000000000000000;
    assign weights1[8][730] = 16'b1111111111111011;
    assign weights1[8][731] = 16'b1111111111111001;
    assign weights1[8][732] = 16'b1111111111110101;
    assign weights1[8][733] = 16'b1111111111110000;
    assign weights1[8][734] = 16'b1111111111011101;
    assign weights1[8][735] = 16'b1111111111100010;
    assign weights1[8][736] = 16'b1111111111100001;
    assign weights1[8][737] = 16'b1111111111011101;
    assign weights1[8][738] = 16'b1111111111001110;
    assign weights1[8][739] = 16'b1111111111010100;
    assign weights1[8][740] = 16'b1111111111001111;
    assign weights1[8][741] = 16'b1111111111000110;
    assign weights1[8][742] = 16'b1111111111001001;
    assign weights1[8][743] = 16'b1111111110101011;
    assign weights1[8][744] = 16'b1111111111001110;
    assign weights1[8][745] = 16'b1111111110111101;
    assign weights1[8][746] = 16'b1111111110111000;
    assign weights1[8][747] = 16'b1111111110101101;
    assign weights1[8][748] = 16'b1111111110110100;
    assign weights1[8][749] = 16'b1111111111000010;
    assign weights1[8][750] = 16'b1111111111010101;
    assign weights1[8][751] = 16'b1111111111011000;
    assign weights1[8][752] = 16'b1111111111100100;
    assign weights1[8][753] = 16'b1111111111110100;
    assign weights1[8][754] = 16'b1111111111111010;
    assign weights1[8][755] = 16'b1111111111111100;
    assign weights1[8][756] = 16'b1111111111111110;
    assign weights1[8][757] = 16'b0000000000000000;
    assign weights1[8][758] = 16'b1111111111111111;
    assign weights1[8][759] = 16'b1111111111111000;
    assign weights1[8][760] = 16'b1111111111110011;
    assign weights1[8][761] = 16'b1111111111101111;
    assign weights1[8][762] = 16'b1111111111100101;
    assign weights1[8][763] = 16'b1111111111001110;
    assign weights1[8][764] = 16'b1111111111001100;
    assign weights1[8][765] = 16'b1111111111001101;
    assign weights1[8][766] = 16'b1111111110111000;
    assign weights1[8][767] = 16'b1111111111000111;
    assign weights1[8][768] = 16'b1111111111000011;
    assign weights1[8][769] = 16'b1111111110110110;
    assign weights1[8][770] = 16'b1111111110101110;
    assign weights1[8][771] = 16'b1111111110110101;
    assign weights1[8][772] = 16'b1111111111000001;
    assign weights1[8][773] = 16'b1111111111000001;
    assign weights1[8][774] = 16'b1111111111001101;
    assign weights1[8][775] = 16'b1111111111010010;
    assign weights1[8][776] = 16'b1111111111010110;
    assign weights1[8][777] = 16'b1111111111010110;
    assign weights1[8][778] = 16'b1111111111101000;
    assign weights1[8][779] = 16'b1111111111101101;
    assign weights1[8][780] = 16'b1111111111101110;
    assign weights1[8][781] = 16'b1111111111111010;
    assign weights1[8][782] = 16'b1111111111111101;
    assign weights1[8][783] = 16'b1111111111111110;
    assign weights1[9][0] = 16'b0000000000000000;
    assign weights1[9][1] = 16'b0000000000000000;
    assign weights1[9][2] = 16'b1111111111111111;
    assign weights1[9][3] = 16'b1111111111111111;
    assign weights1[9][4] = 16'b1111111111111111;
    assign weights1[9][5] = 16'b1111111111111101;
    assign weights1[9][6] = 16'b1111111111111100;
    assign weights1[9][7] = 16'b1111111111111100;
    assign weights1[9][8] = 16'b1111111111110101;
    assign weights1[9][9] = 16'b1111111111110101;
    assign weights1[9][10] = 16'b1111111111110111;
    assign weights1[9][11] = 16'b1111111111110111;
    assign weights1[9][12] = 16'b1111111111110010;
    assign weights1[9][13] = 16'b1111111111110100;
    assign weights1[9][14] = 16'b1111111111101110;
    assign weights1[9][15] = 16'b1111111111101100;
    assign weights1[9][16] = 16'b1111111111101001;
    assign weights1[9][17] = 16'b1111111111101011;
    assign weights1[9][18] = 16'b1111111111101101;
    assign weights1[9][19] = 16'b1111111111101111;
    assign weights1[9][20] = 16'b1111111111101110;
    assign weights1[9][21] = 16'b1111111111101010;
    assign weights1[9][22] = 16'b1111111111110010;
    assign weights1[9][23] = 16'b1111111111110110;
    assign weights1[9][24] = 16'b1111111111110110;
    assign weights1[9][25] = 16'b1111111111111000;
    assign weights1[9][26] = 16'b1111111111111111;
    assign weights1[9][27] = 16'b0000000000000000;
    assign weights1[9][28] = 16'b1111111111111110;
    assign weights1[9][29] = 16'b1111111111111111;
    assign weights1[9][30] = 16'b1111111111111110;
    assign weights1[9][31] = 16'b1111111111111010;
    assign weights1[9][32] = 16'b1111111111111011;
    assign weights1[9][33] = 16'b1111111111111010;
    assign weights1[9][34] = 16'b1111111111111000;
    assign weights1[9][35] = 16'b0000000000000000;
    assign weights1[9][36] = 16'b1111111111110101;
    assign weights1[9][37] = 16'b1111111111111000;
    assign weights1[9][38] = 16'b1111111111110111;
    assign weights1[9][39] = 16'b1111111111110110;
    assign weights1[9][40] = 16'b0000000000000001;
    assign weights1[9][41] = 16'b1111111111101000;
    assign weights1[9][42] = 16'b1111111111011111;
    assign weights1[9][43] = 16'b1111111111110001;
    assign weights1[9][44] = 16'b1111111111110000;
    assign weights1[9][45] = 16'b1111111111110010;
    assign weights1[9][46] = 16'b1111111111110000;
    assign weights1[9][47] = 16'b1111111111110001;
    assign weights1[9][48] = 16'b1111111111110001;
    assign weights1[9][49] = 16'b1111111111110100;
    assign weights1[9][50] = 16'b1111111111100110;
    assign weights1[9][51] = 16'b1111111111101000;
    assign weights1[9][52] = 16'b1111111111101111;
    assign weights1[9][53] = 16'b1111111111111010;
    assign weights1[9][54] = 16'b1111111111110111;
    assign weights1[9][55] = 16'b1111111111111110;
    assign weights1[9][56] = 16'b1111111111111100;
    assign weights1[9][57] = 16'b1111111111111010;
    assign weights1[9][58] = 16'b1111111111111100;
    assign weights1[9][59] = 16'b1111111111110111;
    assign weights1[9][60] = 16'b1111111111110110;
    assign weights1[9][61] = 16'b1111111111111001;
    assign weights1[9][62] = 16'b0000000000000000;
    assign weights1[9][63] = 16'b0000000000000100;
    assign weights1[9][64] = 16'b0000000000000000;
    assign weights1[9][65] = 16'b0000000000000000;
    assign weights1[9][66] = 16'b1111111111111001;
    assign weights1[9][67] = 16'b1111111111110100;
    assign weights1[9][68] = 16'b1111111111110101;
    assign weights1[9][69] = 16'b1111111111100011;
    assign weights1[9][70] = 16'b1111111111111011;
    assign weights1[9][71] = 16'b1111111111101111;
    assign weights1[9][72] = 16'b1111111111111000;
    assign weights1[9][73] = 16'b1111111111100110;
    assign weights1[9][74] = 16'b1111111111110001;
    assign weights1[9][75] = 16'b1111111111110100;
    assign weights1[9][76] = 16'b1111111111100001;
    assign weights1[9][77] = 16'b1111111111110001;
    assign weights1[9][78] = 16'b1111111111110111;
    assign weights1[9][79] = 16'b1111111111101110;
    assign weights1[9][80] = 16'b1111111111110101;
    assign weights1[9][81] = 16'b1111111111111001;
    assign weights1[9][82] = 16'b1111111111110011;
    assign weights1[9][83] = 16'b1111111111110101;
    assign weights1[9][84] = 16'b1111111111111100;
    assign weights1[9][85] = 16'b1111111111111110;
    assign weights1[9][86] = 16'b1111111111111001;
    assign weights1[9][87] = 16'b1111111111110100;
    assign weights1[9][88] = 16'b1111111111110110;
    assign weights1[9][89] = 16'b1111111111110101;
    assign weights1[9][90] = 16'b1111111111110110;
    assign weights1[9][91] = 16'b1111111111111011;
    assign weights1[9][92] = 16'b1111111111110110;
    assign weights1[9][93] = 16'b1111111111111010;
    assign weights1[9][94] = 16'b1111111111110011;
    assign weights1[9][95] = 16'b1111111111111100;
    assign weights1[9][96] = 16'b1111111111111010;
    assign weights1[9][97] = 16'b0000000000000000;
    assign weights1[9][98] = 16'b1111111111110100;
    assign weights1[9][99] = 16'b1111111111111111;
    assign weights1[9][100] = 16'b0000000000001001;
    assign weights1[9][101] = 16'b1111111111111010;
    assign weights1[9][102] = 16'b1111111111101110;
    assign weights1[9][103] = 16'b0000000000000001;
    assign weights1[9][104] = 16'b1111111111110111;
    assign weights1[9][105] = 16'b1111111111110011;
    assign weights1[9][106] = 16'b1111111111111100;
    assign weights1[9][107] = 16'b1111111111110100;
    assign weights1[9][108] = 16'b1111111111110100;
    assign weights1[9][109] = 16'b1111111111111001;
    assign weights1[9][110] = 16'b1111111111110100;
    assign weights1[9][111] = 16'b1111111111111011;
    assign weights1[9][112] = 16'b1111111111111101;
    assign weights1[9][113] = 16'b1111111111111110;
    assign weights1[9][114] = 16'b1111111111110101;
    assign weights1[9][115] = 16'b1111111111110110;
    assign weights1[9][116] = 16'b1111111111110011;
    assign weights1[9][117] = 16'b1111111111110100;
    assign weights1[9][118] = 16'b1111111111100110;
    assign weights1[9][119] = 16'b1111111111100101;
    assign weights1[9][120] = 16'b1111111111110110;
    assign weights1[9][121] = 16'b1111111111110011;
    assign weights1[9][122] = 16'b1111111111101111;
    assign weights1[9][123] = 16'b1111111111111111;
    assign weights1[9][124] = 16'b1111111111111011;
    assign weights1[9][125] = 16'b1111111111101010;
    assign weights1[9][126] = 16'b1111111111111001;
    assign weights1[9][127] = 16'b1111111111110111;
    assign weights1[9][128] = 16'b1111111111011001;
    assign weights1[9][129] = 16'b0000000000000110;
    assign weights1[9][130] = 16'b1111111111101110;
    assign weights1[9][131] = 16'b1111111111101100;
    assign weights1[9][132] = 16'b0000000000000111;
    assign weights1[9][133] = 16'b1111111111110110;
    assign weights1[9][134] = 16'b0000000000001011;
    assign weights1[9][135] = 16'b1111111111110000;
    assign weights1[9][136] = 16'b0000000000010101;
    assign weights1[9][137] = 16'b0000000000000000;
    assign weights1[9][138] = 16'b1111111111110111;
    assign weights1[9][139] = 16'b1111111111111001;
    assign weights1[9][140] = 16'b1111111111111111;
    assign weights1[9][141] = 16'b1111111111111100;
    assign weights1[9][142] = 16'b0000000000000011;
    assign weights1[9][143] = 16'b1111111111111001;
    assign weights1[9][144] = 16'b1111111111110001;
    assign weights1[9][145] = 16'b1111111111110000;
    assign weights1[9][146] = 16'b0000000000000010;
    assign weights1[9][147] = 16'b1111111111101111;
    assign weights1[9][148] = 16'b1111111111110101;
    assign weights1[9][149] = 16'b1111111111111111;
    assign weights1[9][150] = 16'b1111111111111111;
    assign weights1[9][151] = 16'b1111111111101110;
    assign weights1[9][152] = 16'b1111111111110000;
    assign weights1[9][153] = 16'b0000000000000001;
    assign weights1[9][154] = 16'b1111111111111000;
    assign weights1[9][155] = 16'b1111111111100010;
    assign weights1[9][156] = 16'b0000000000000101;
    assign weights1[9][157] = 16'b1111111111110010;
    assign weights1[9][158] = 16'b1111111111111101;
    assign weights1[9][159] = 16'b0000000000000010;
    assign weights1[9][160] = 16'b1111111111101111;
    assign weights1[9][161] = 16'b1111111111100010;
    assign weights1[9][162] = 16'b0000000000001000;
    assign weights1[9][163] = 16'b0000000000011001;
    assign weights1[9][164] = 16'b0000000000000101;
    assign weights1[9][165] = 16'b1111111111101111;
    assign weights1[9][166] = 16'b1111111111111000;
    assign weights1[9][167] = 16'b1111111111110101;
    assign weights1[9][168] = 16'b1111111111111111;
    assign weights1[9][169] = 16'b0000000000000010;
    assign weights1[9][170] = 16'b1111111111111111;
    assign weights1[9][171] = 16'b1111111111110000;
    assign weights1[9][172] = 16'b1111111111110101;
    assign weights1[9][173] = 16'b0000000000000101;
    assign weights1[9][174] = 16'b1111111111011011;
    assign weights1[9][175] = 16'b1111111111110110;
    assign weights1[9][176] = 16'b1111111111011011;
    assign weights1[9][177] = 16'b1111111111011010;
    assign weights1[9][178] = 16'b1111111111111010;
    assign weights1[9][179] = 16'b1111111111100101;
    assign weights1[9][180] = 16'b1111111111110110;
    assign weights1[9][181] = 16'b1111111111110011;
    assign weights1[9][182] = 16'b1111111111111100;
    assign weights1[9][183] = 16'b1111111111101100;
    assign weights1[9][184] = 16'b1111111111111110;
    assign weights1[9][185] = 16'b1111111111111110;
    assign weights1[9][186] = 16'b1111111111111001;
    assign weights1[9][187] = 16'b1111111111111001;
    assign weights1[9][188] = 16'b0000000000000111;
    assign weights1[9][189] = 16'b0000000000000100;
    assign weights1[9][190] = 16'b1111111111010100;
    assign weights1[9][191] = 16'b1111111111101001;
    assign weights1[9][192] = 16'b0000000000001011;
    assign weights1[9][193] = 16'b1111111111110111;
    assign weights1[9][194] = 16'b1111111111110110;
    assign weights1[9][195] = 16'b1111111111110110;
    assign weights1[9][196] = 16'b0000000000000100;
    assign weights1[9][197] = 16'b0000000000000010;
    assign weights1[9][198] = 16'b0000000000000101;
    assign weights1[9][199] = 16'b1111111111110111;
    assign weights1[9][200] = 16'b1111111111110111;
    assign weights1[9][201] = 16'b1111111111100000;
    assign weights1[9][202] = 16'b1111111111100010;
    assign weights1[9][203] = 16'b1111111111100001;
    assign weights1[9][204] = 16'b1111111111111100;
    assign weights1[9][205] = 16'b1111111111101110;
    assign weights1[9][206] = 16'b1111111111100011;
    assign weights1[9][207] = 16'b1111111111100011;
    assign weights1[9][208] = 16'b1111111111011101;
    assign weights1[9][209] = 16'b1111111111110001;
    assign weights1[9][210] = 16'b1111111111101101;
    assign weights1[9][211] = 16'b0000000000000001;
    assign weights1[9][212] = 16'b1111111111101110;
    assign weights1[9][213] = 16'b0000000000001000;
    assign weights1[9][214] = 16'b1111111111101100;
    assign weights1[9][215] = 16'b1111111111101110;
    assign weights1[9][216] = 16'b1111111111011100;
    assign weights1[9][217] = 16'b1111111111100001;
    assign weights1[9][218] = 16'b1111111111111100;
    assign weights1[9][219] = 16'b1111111111011001;
    assign weights1[9][220] = 16'b1111111111101011;
    assign weights1[9][221] = 16'b1111111111101000;
    assign weights1[9][222] = 16'b1111111111110001;
    assign weights1[9][223] = 16'b1111111111100110;
    assign weights1[9][224] = 16'b0000000000000010;
    assign weights1[9][225] = 16'b0000000000000100;
    assign weights1[9][226] = 16'b0000000000001011;
    assign weights1[9][227] = 16'b1111111111111101;
    assign weights1[9][228] = 16'b1111111111110111;
    assign weights1[9][229] = 16'b1111111111010100;
    assign weights1[9][230] = 16'b1111111111011010;
    assign weights1[9][231] = 16'b1111111111110000;
    assign weights1[9][232] = 16'b1111111111011011;
    assign weights1[9][233] = 16'b1111111111001100;
    assign weights1[9][234] = 16'b1111111111100101;
    assign weights1[9][235] = 16'b1111111111011000;
    assign weights1[9][236] = 16'b1111111111111001;
    assign weights1[9][237] = 16'b1111111111011011;
    assign weights1[9][238] = 16'b1111111111100111;
    assign weights1[9][239] = 16'b1111111111100000;
    assign weights1[9][240] = 16'b1111111111110001;
    assign weights1[9][241] = 16'b1111111111100001;
    assign weights1[9][242] = 16'b1111111111110000;
    assign weights1[9][243] = 16'b1111111111100001;
    assign weights1[9][244] = 16'b0000000000000101;
    assign weights1[9][245] = 16'b1111111111110001;
    assign weights1[9][246] = 16'b1111111111111100;
    assign weights1[9][247] = 16'b1111111111101000;
    assign weights1[9][248] = 16'b1111111111001111;
    assign weights1[9][249] = 16'b1111111111011000;
    assign weights1[9][250] = 16'b1111111111110100;
    assign weights1[9][251] = 16'b1111111111100000;
    assign weights1[9][252] = 16'b0000000000000001;
    assign weights1[9][253] = 16'b0000000000000010;
    assign weights1[9][254] = 16'b0000000000001000;
    assign weights1[9][255] = 16'b0000000000000011;
    assign weights1[9][256] = 16'b1111111111110111;
    assign weights1[9][257] = 16'b1111111111100001;
    assign weights1[9][258] = 16'b1111111111100110;
    assign weights1[9][259] = 16'b1111111111101000;
    assign weights1[9][260] = 16'b1111111111010100;
    assign weights1[9][261] = 16'b1111111111110010;
    assign weights1[9][262] = 16'b1111111111100010;
    assign weights1[9][263] = 16'b1111111111100011;
    assign weights1[9][264] = 16'b1111111111100011;
    assign weights1[9][265] = 16'b1111111111101010;
    assign weights1[9][266] = 16'b1111111111101011;
    assign weights1[9][267] = 16'b1111111111011000;
    assign weights1[9][268] = 16'b1111111111101101;
    assign weights1[9][269] = 16'b1111111111011000;
    assign weights1[9][270] = 16'b1111111111101000;
    assign weights1[9][271] = 16'b1111111111100000;
    assign weights1[9][272] = 16'b1111111111010100;
    assign weights1[9][273] = 16'b1111111111011011;
    assign weights1[9][274] = 16'b1111111111100001;
    assign weights1[9][275] = 16'b1111111111011010;
    assign weights1[9][276] = 16'b1111111111100100;
    assign weights1[9][277] = 16'b1111111111100000;
    assign weights1[9][278] = 16'b1111111111011110;
    assign weights1[9][279] = 16'b1111111111011011;
    assign weights1[9][280] = 16'b0000000000000011;
    assign weights1[9][281] = 16'b1111111111111101;
    assign weights1[9][282] = 16'b1111111111111011;
    assign weights1[9][283] = 16'b1111111111101111;
    assign weights1[9][284] = 16'b1111111111011111;
    assign weights1[9][285] = 16'b1111111111101000;
    assign weights1[9][286] = 16'b1111111111111001;
    assign weights1[9][287] = 16'b1111111111110000;
    assign weights1[9][288] = 16'b1111111111010010;
    assign weights1[9][289] = 16'b1111111111100001;
    assign weights1[9][290] = 16'b1111111111101001;
    assign weights1[9][291] = 16'b1111111111011001;
    assign weights1[9][292] = 16'b1111111111100010;
    assign weights1[9][293] = 16'b1111111111100100;
    assign weights1[9][294] = 16'b1111111111011110;
    assign weights1[9][295] = 16'b1111111111011000;
    assign weights1[9][296] = 16'b1111111111010111;
    assign weights1[9][297] = 16'b1111111111100010;
    assign weights1[9][298] = 16'b1111111111011011;
    assign weights1[9][299] = 16'b1111111111011000;
    assign weights1[9][300] = 16'b1111111111100001;
    assign weights1[9][301] = 16'b1111111111011011;
    assign weights1[9][302] = 16'b1111111111011010;
    assign weights1[9][303] = 16'b1111111111011110;
    assign weights1[9][304] = 16'b1111111111001101;
    assign weights1[9][305] = 16'b1111111111100001;
    assign weights1[9][306] = 16'b1111111111011001;
    assign weights1[9][307] = 16'b1111111111011011;
    assign weights1[9][308] = 16'b1111111111111111;
    assign weights1[9][309] = 16'b1111111111111100;
    assign weights1[9][310] = 16'b0000000000000100;
    assign weights1[9][311] = 16'b1111111111110110;
    assign weights1[9][312] = 16'b1111111111110111;
    assign weights1[9][313] = 16'b1111111111110001;
    assign weights1[9][314] = 16'b1111111111111100;
    assign weights1[9][315] = 16'b1111111111111001;
    assign weights1[9][316] = 16'b1111111111110100;
    assign weights1[9][317] = 16'b1111111111111001;
    assign weights1[9][318] = 16'b1111111111110011;
    assign weights1[9][319] = 16'b1111111111010010;
    assign weights1[9][320] = 16'b1111111111100111;
    assign weights1[9][321] = 16'b1111111111011100;
    assign weights1[9][322] = 16'b1111111111010111;
    assign weights1[9][323] = 16'b1111111111101000;
    assign weights1[9][324] = 16'b1111111111100110;
    assign weights1[9][325] = 16'b1111111111011101;
    assign weights1[9][326] = 16'b1111111111100010;
    assign weights1[9][327] = 16'b1111111111111000;
    assign weights1[9][328] = 16'b1111111111011100;
    assign weights1[9][329] = 16'b1111111111100111;
    assign weights1[9][330] = 16'b1111111111010011;
    assign weights1[9][331] = 16'b1111111111010101;
    assign weights1[9][332] = 16'b1111111111000110;
    assign weights1[9][333] = 16'b1111111111011000;
    assign weights1[9][334] = 16'b1111111111011001;
    assign weights1[9][335] = 16'b1111111111100110;
    assign weights1[9][336] = 16'b0000000000000000;
    assign weights1[9][337] = 16'b0000000000000011;
    assign weights1[9][338] = 16'b1111111111111110;
    assign weights1[9][339] = 16'b0000000000001110;
    assign weights1[9][340] = 16'b0000000000000000;
    assign weights1[9][341] = 16'b0000000000000111;
    assign weights1[9][342] = 16'b1111111111110100;
    assign weights1[9][343] = 16'b1111111111110000;
    assign weights1[9][344] = 16'b0000000000000000;
    assign weights1[9][345] = 16'b1111111111011100;
    assign weights1[9][346] = 16'b1111111111101010;
    assign weights1[9][347] = 16'b1111111111010100;
    assign weights1[9][348] = 16'b1111111111110011;
    assign weights1[9][349] = 16'b1111111111011010;
    assign weights1[9][350] = 16'b1111111111110000;
    assign weights1[9][351] = 16'b1111111111110011;
    assign weights1[9][352] = 16'b1111111111010110;
    assign weights1[9][353] = 16'b1111111111100101;
    assign weights1[9][354] = 16'b1111111111100101;
    assign weights1[9][355] = 16'b1111111111100010;
    assign weights1[9][356] = 16'b1111111111001100;
    assign weights1[9][357] = 16'b1111111111101010;
    assign weights1[9][358] = 16'b1111111111011111;
    assign weights1[9][359] = 16'b1111111111010111;
    assign weights1[9][360] = 16'b1111111111000001;
    assign weights1[9][361] = 16'b1111111111011111;
    assign weights1[9][362] = 16'b1111111111101001;
    assign weights1[9][363] = 16'b1111111111100101;
    assign weights1[9][364] = 16'b1111111111111101;
    assign weights1[9][365] = 16'b0000000000001110;
    assign weights1[9][366] = 16'b0000000000000101;
    assign weights1[9][367] = 16'b0000000000110010;
    assign weights1[9][368] = 16'b0000000000010100;
    assign weights1[9][369] = 16'b0000000000000000;
    assign weights1[9][370] = 16'b0000000000100110;
    assign weights1[9][371] = 16'b1111111111101101;
    assign weights1[9][372] = 16'b1111111111111000;
    assign weights1[9][373] = 16'b1111111111111010;
    assign weights1[9][374] = 16'b0000000000001011;
    assign weights1[9][375] = 16'b1111111111101110;
    assign weights1[9][376] = 16'b1111111111011100;
    assign weights1[9][377] = 16'b1111111111101010;
    assign weights1[9][378] = 16'b1111111111110101;
    assign weights1[9][379] = 16'b1111111111010111;
    assign weights1[9][380] = 16'b1111111111100101;
    assign weights1[9][381] = 16'b1111111111111011;
    assign weights1[9][382] = 16'b1111111111100101;
    assign weights1[9][383] = 16'b1111111110111101;
    assign weights1[9][384] = 16'b1111111111100000;
    assign weights1[9][385] = 16'b1111111111100111;
    assign weights1[9][386] = 16'b1111111111101000;
    assign weights1[9][387] = 16'b1111111111101011;
    assign weights1[9][388] = 16'b1111111111101110;
    assign weights1[9][389] = 16'b1111111111100010;
    assign weights1[9][390] = 16'b1111111111110010;
    assign weights1[9][391] = 16'b1111111111101111;
    assign weights1[9][392] = 16'b1111111111111111;
    assign weights1[9][393] = 16'b0000000000010101;
    assign weights1[9][394] = 16'b0000000000110000;
    assign weights1[9][395] = 16'b0000000000110111;
    assign weights1[9][396] = 16'b0000000000111010;
    assign weights1[9][397] = 16'b0000000000010100;
    assign weights1[9][398] = 16'b0000000000011011;
    assign weights1[9][399] = 16'b0000000000011111;
    assign weights1[9][400] = 16'b1111111111110111;
    assign weights1[9][401] = 16'b0000000000000100;
    assign weights1[9][402] = 16'b1111111111001101;
    assign weights1[9][403] = 16'b1111111111100000;
    assign weights1[9][404] = 16'b1111111111101100;
    assign weights1[9][405] = 16'b1111111111100101;
    assign weights1[9][406] = 16'b1111111111100011;
    assign weights1[9][407] = 16'b1111111111100100;
    assign weights1[9][408] = 16'b1111111111110100;
    assign weights1[9][409] = 16'b1111111111111111;
    assign weights1[9][410] = 16'b1111111111110001;
    assign weights1[9][411] = 16'b1111111111101110;
    assign weights1[9][412] = 16'b0000000000001001;
    assign weights1[9][413] = 16'b0000000000001000;
    assign weights1[9][414] = 16'b1111111111111010;
    assign weights1[9][415] = 16'b0000000000001000;
    assign weights1[9][416] = 16'b0000000000001001;
    assign weights1[9][417] = 16'b0000000000011000;
    assign weights1[9][418] = 16'b0000000000000000;
    assign weights1[9][419] = 16'b1111111111111111;
    assign weights1[9][420] = 16'b0000000000010100;
    assign weights1[9][421] = 16'b0000000000011011;
    assign weights1[9][422] = 16'b0000000000111011;
    assign weights1[9][423] = 16'b0000000000110011;
    assign weights1[9][424] = 16'b0000000001000010;
    assign weights1[9][425] = 16'b0000000000101010;
    assign weights1[9][426] = 16'b0000000000110100;
    assign weights1[9][427] = 16'b0000000000100110;
    assign weights1[9][428] = 16'b0000000000100101;
    assign weights1[9][429] = 16'b0000000000100001;
    assign weights1[9][430] = 16'b0000000000001111;
    assign weights1[9][431] = 16'b1111111111101001;
    assign weights1[9][432] = 16'b1111111111111110;
    assign weights1[9][433] = 16'b0000000000000001;
    assign weights1[9][434] = 16'b1111111111110010;
    assign weights1[9][435] = 16'b1111111111101101;
    assign weights1[9][436] = 16'b1111111111101111;
    assign weights1[9][437] = 16'b0000000000000110;
    assign weights1[9][438] = 16'b1111111111111011;
    assign weights1[9][439] = 16'b0000000000011011;
    assign weights1[9][440] = 16'b0000000000010111;
    assign weights1[9][441] = 16'b0000000000001110;
    assign weights1[9][442] = 16'b0000000000001010;
    assign weights1[9][443] = 16'b1111111111101000;
    assign weights1[9][444] = 16'b0000000000010001;
    assign weights1[9][445] = 16'b0000000000100111;
    assign weights1[9][446] = 16'b0000000000100001;
    assign weights1[9][447] = 16'b0000000000011000;
    assign weights1[9][448] = 16'b0000000000011010;
    assign weights1[9][449] = 16'b0000000000011110;
    assign weights1[9][450] = 16'b0000000000101000;
    assign weights1[9][451] = 16'b0000000000110001;
    assign weights1[9][452] = 16'b0000000000111001;
    assign weights1[9][453] = 16'b0000000001001010;
    assign weights1[9][454] = 16'b0000000000110110;
    assign weights1[9][455] = 16'b0000000001000110;
    assign weights1[9][456] = 16'b0000000001000100;
    assign weights1[9][457] = 16'b0000000001000010;
    assign weights1[9][458] = 16'b0000000001001101;
    assign weights1[9][459] = 16'b0000000000100100;
    assign weights1[9][460] = 16'b0000000000101010;
    assign weights1[9][461] = 16'b0000000000100110;
    assign weights1[9][462] = 16'b0000000000011011;
    assign weights1[9][463] = 16'b0000000000010111;
    assign weights1[9][464] = 16'b0000000000001110;
    assign weights1[9][465] = 16'b0000000000011010;
    assign weights1[9][466] = 16'b0000000000010010;
    assign weights1[9][467] = 16'b0000000000010001;
    assign weights1[9][468] = 16'b0000000000101001;
    assign weights1[9][469] = 16'b0000000000110001;
    assign weights1[9][470] = 16'b0000000000100001;
    assign weights1[9][471] = 16'b0000000000010010;
    assign weights1[9][472] = 16'b0000000000101001;
    assign weights1[9][473] = 16'b0000000000111100;
    assign weights1[9][474] = 16'b0000000000101111;
    assign weights1[9][475] = 16'b0000000000011100;
    assign weights1[9][476] = 16'b0000000000011000;
    assign weights1[9][477] = 16'b0000000000100011;
    assign weights1[9][478] = 16'b0000000000101101;
    assign weights1[9][479] = 16'b0000000000011011;
    assign weights1[9][480] = 16'b0000000000011110;
    assign weights1[9][481] = 16'b0000000000101001;
    assign weights1[9][482] = 16'b0000000000100110;
    assign weights1[9][483] = 16'b0000000000110000;
    assign weights1[9][484] = 16'b0000000001010100;
    assign weights1[9][485] = 16'b0000000000111100;
    assign weights1[9][486] = 16'b0000000000110110;
    assign weights1[9][487] = 16'b0000000000111101;
    assign weights1[9][488] = 16'b0000000000101101;
    assign weights1[9][489] = 16'b0000000001000001;
    assign weights1[9][490] = 16'b0000000000101111;
    assign weights1[9][491] = 16'b0000000000100110;
    assign weights1[9][492] = 16'b0000000000110110;
    assign weights1[9][493] = 16'b0000000000100101;
    assign weights1[9][494] = 16'b0000000000101111;
    assign weights1[9][495] = 16'b0000000000101001;
    assign weights1[9][496] = 16'b0000000000111011;
    assign weights1[9][497] = 16'b0000000001000000;
    assign weights1[9][498] = 16'b0000000001010001;
    assign weights1[9][499] = 16'b0000000000101010;
    assign weights1[9][500] = 16'b0000000000110111;
    assign weights1[9][501] = 16'b0000000001010000;
    assign weights1[9][502] = 16'b0000000000101110;
    assign weights1[9][503] = 16'b0000000000101110;
    assign weights1[9][504] = 16'b0000000000001001;
    assign weights1[9][505] = 16'b0000000000010101;
    assign weights1[9][506] = 16'b0000000000011101;
    assign weights1[9][507] = 16'b0000000000011011;
    assign weights1[9][508] = 16'b0000000000100110;
    assign weights1[9][509] = 16'b0000000000100011;
    assign weights1[9][510] = 16'b0000000000101010;
    assign weights1[9][511] = 16'b0000000000110010;
    assign weights1[9][512] = 16'b0000000000101000;
    assign weights1[9][513] = 16'b0000000000100110;
    assign weights1[9][514] = 16'b0000000001000111;
    assign weights1[9][515] = 16'b0000000000101000;
    assign weights1[9][516] = 16'b0000000001001111;
    assign weights1[9][517] = 16'b0000000000110100;
    assign weights1[9][518] = 16'b0000000001010000;
    assign weights1[9][519] = 16'b0000000000101011;
    assign weights1[9][520] = 16'b0000000000111010;
    assign weights1[9][521] = 16'b0000000000110101;
    assign weights1[9][522] = 16'b0000000000101001;
    assign weights1[9][523] = 16'b0000000000110100;
    assign weights1[9][524] = 16'b0000000000111010;
    assign weights1[9][525] = 16'b0000000000111010;
    assign weights1[9][526] = 16'b0000000000111000;
    assign weights1[9][527] = 16'b0000000000100111;
    assign weights1[9][528] = 16'b0000000001010010;
    assign weights1[9][529] = 16'b0000000001000001;
    assign weights1[9][530] = 16'b0000000000110100;
    assign weights1[9][531] = 16'b0000000000101010;
    assign weights1[9][532] = 16'b0000000000001001;
    assign weights1[9][533] = 16'b0000000000001011;
    assign weights1[9][534] = 16'b0000000000001010;
    assign weights1[9][535] = 16'b0000000000001101;
    assign weights1[9][536] = 16'b0000000000010010;
    assign weights1[9][537] = 16'b0000000000001010;
    assign weights1[9][538] = 16'b0000000000011001;
    assign weights1[9][539] = 16'b0000000000100000;
    assign weights1[9][540] = 16'b0000000000110000;
    assign weights1[9][541] = 16'b0000000000110110;
    assign weights1[9][542] = 16'b0000000000101101;
    assign weights1[9][543] = 16'b0000000000101110;
    assign weights1[9][544] = 16'b0000000000110110;
    assign weights1[9][545] = 16'b0000000000111011;
    assign weights1[9][546] = 16'b0000000000110011;
    assign weights1[9][547] = 16'b0000000000110101;
    assign weights1[9][548] = 16'b0000000000101010;
    assign weights1[9][549] = 16'b0000000000110100;
    assign weights1[9][550] = 16'b0000000000111000;
    assign weights1[9][551] = 16'b0000000000111010;
    assign weights1[9][552] = 16'b0000000000101110;
    assign weights1[9][553] = 16'b0000000001000110;
    assign weights1[9][554] = 16'b0000000000111110;
    assign weights1[9][555] = 16'b0000000000111000;
    assign weights1[9][556] = 16'b0000000000101100;
    assign weights1[9][557] = 16'b0000000000100101;
    assign weights1[9][558] = 16'b0000000000101110;
    assign weights1[9][559] = 16'b0000000000100100;
    assign weights1[9][560] = 16'b0000000000001000;
    assign weights1[9][561] = 16'b0000000000000010;
    assign weights1[9][562] = 16'b1111111111111111;
    assign weights1[9][563] = 16'b0000000000000101;
    assign weights1[9][564] = 16'b0000000000010001;
    assign weights1[9][565] = 16'b0000000000001100;
    assign weights1[9][566] = 16'b1111111111110100;
    assign weights1[9][567] = 16'b0000000000011001;
    assign weights1[9][568] = 16'b0000000000000110;
    assign weights1[9][569] = 16'b0000000000000100;
    assign weights1[9][570] = 16'b0000000000010100;
    assign weights1[9][571] = 16'b0000000000101011;
    assign weights1[9][572] = 16'b0000000000011010;
    assign weights1[9][573] = 16'b0000000000001101;
    assign weights1[9][574] = 16'b0000000000011101;
    assign weights1[9][575] = 16'b0000000000110101;
    assign weights1[9][576] = 16'b0000000000100111;
    assign weights1[9][577] = 16'b0000000000101110;
    assign weights1[9][578] = 16'b0000000001000111;
    assign weights1[9][579] = 16'b0000000000110101;
    assign weights1[9][580] = 16'b0000000000110100;
    assign weights1[9][581] = 16'b1111111111111001;
    assign weights1[9][582] = 16'b0000000000101100;
    assign weights1[9][583] = 16'b0000000000011000;
    assign weights1[9][584] = 16'b0000000000010010;
    assign weights1[9][585] = 16'b0000000000010001;
    assign weights1[9][586] = 16'b0000000000100011;
    assign weights1[9][587] = 16'b0000000000100000;
    assign weights1[9][588] = 16'b0000000000000000;
    assign weights1[9][589] = 16'b1111111111111011;
    assign weights1[9][590] = 16'b1111111111110110;
    assign weights1[9][591] = 16'b1111111111110101;
    assign weights1[9][592] = 16'b0000000000001001;
    assign weights1[9][593] = 16'b0000000000010100;
    assign weights1[9][594] = 16'b0000000000010101;
    assign weights1[9][595] = 16'b0000000000000000;
    assign weights1[9][596] = 16'b1111111111110110;
    assign weights1[9][597] = 16'b0000000000001010;
    assign weights1[9][598] = 16'b0000000000000111;
    assign weights1[9][599] = 16'b1111111111111010;
    assign weights1[9][600] = 16'b0000000000001011;
    assign weights1[9][601] = 16'b0000000000011001;
    assign weights1[9][602] = 16'b0000000000011101;
    assign weights1[9][603] = 16'b1111111111111000;
    assign weights1[9][604] = 16'b0000000000100000;
    assign weights1[9][605] = 16'b0000000000010001;
    assign weights1[9][606] = 16'b0000000000001000;
    assign weights1[9][607] = 16'b0000000000000100;
    assign weights1[9][608] = 16'b0000000000011110;
    assign weights1[9][609] = 16'b0000000000011110;
    assign weights1[9][610] = 16'b0000000000100101;
    assign weights1[9][611] = 16'b0000000000010111;
    assign weights1[9][612] = 16'b0000000000010000;
    assign weights1[9][613] = 16'b0000000000001110;
    assign weights1[9][614] = 16'b0000000000010100;
    assign weights1[9][615] = 16'b0000000000001010;
    assign weights1[9][616] = 16'b0000000000000000;
    assign weights1[9][617] = 16'b1111111111110100;
    assign weights1[9][618] = 16'b1111111111100111;
    assign weights1[9][619] = 16'b1111111111111110;
    assign weights1[9][620] = 16'b1111111111111110;
    assign weights1[9][621] = 16'b0000000000001011;
    assign weights1[9][622] = 16'b1111111111110110;
    assign weights1[9][623] = 16'b0000000000001100;
    assign weights1[9][624] = 16'b1111111111101111;
    assign weights1[9][625] = 16'b0000000000001101;
    assign weights1[9][626] = 16'b1111111111111011;
    assign weights1[9][627] = 16'b0000000000010001;
    assign weights1[9][628] = 16'b1111111111111111;
    assign weights1[9][629] = 16'b0000000000000000;
    assign weights1[9][630] = 16'b1111111111110000;
    assign weights1[9][631] = 16'b1111111111111010;
    assign weights1[9][632] = 16'b1111111111110101;
    assign weights1[9][633] = 16'b0000000000000111;
    assign weights1[9][634] = 16'b0000000000001001;
    assign weights1[9][635] = 16'b0000000000001100;
    assign weights1[9][636] = 16'b0000000000010100;
    assign weights1[9][637] = 16'b0000000000010001;
    assign weights1[9][638] = 16'b0000000000001101;
    assign weights1[9][639] = 16'b0000000000000010;
    assign weights1[9][640] = 16'b0000000000010001;
    assign weights1[9][641] = 16'b0000000000001100;
    assign weights1[9][642] = 16'b1111111111111110;
    assign weights1[9][643] = 16'b0000000000000110;
    assign weights1[9][644] = 16'b1111111111111010;
    assign weights1[9][645] = 16'b1111111111101100;
    assign weights1[9][646] = 16'b1111111111100000;
    assign weights1[9][647] = 16'b1111111111110001;
    assign weights1[9][648] = 16'b1111111111101011;
    assign weights1[9][649] = 16'b1111111111101001;
    assign weights1[9][650] = 16'b1111111111100111;
    assign weights1[9][651] = 16'b1111111111110110;
    assign weights1[9][652] = 16'b1111111111101001;
    assign weights1[9][653] = 16'b1111111111110011;
    assign weights1[9][654] = 16'b1111111111110100;
    assign weights1[9][655] = 16'b1111111111100110;
    assign weights1[9][656] = 16'b1111111111100010;
    assign weights1[9][657] = 16'b1111111111011110;
    assign weights1[9][658] = 16'b1111111111101100;
    assign weights1[9][659] = 16'b0000000000011101;
    assign weights1[9][660] = 16'b1111111111011010;
    assign weights1[9][661] = 16'b1111111111101101;
    assign weights1[9][662] = 16'b0000000000001001;
    assign weights1[9][663] = 16'b0000000000000001;
    assign weights1[9][664] = 16'b1111111111111110;
    assign weights1[9][665] = 16'b1111111111110101;
    assign weights1[9][666] = 16'b1111111111111111;
    assign weights1[9][667] = 16'b1111111111110110;
    assign weights1[9][668] = 16'b1111111111111111;
    assign weights1[9][669] = 16'b1111111111111011;
    assign weights1[9][670] = 16'b1111111111111101;
    assign weights1[9][671] = 16'b1111111111111110;
    assign weights1[9][672] = 16'b1111111111111100;
    assign weights1[9][673] = 16'b1111111111111011;
    assign weights1[9][674] = 16'b1111111111101010;
    assign weights1[9][675] = 16'b1111111111011111;
    assign weights1[9][676] = 16'b1111111111001111;
    assign weights1[9][677] = 16'b1111111111001111;
    assign weights1[9][678] = 16'b1111111111010011;
    assign weights1[9][679] = 16'b1111111111011000;
    assign weights1[9][680] = 16'b1111111111010000;
    assign weights1[9][681] = 16'b1111111111111101;
    assign weights1[9][682] = 16'b1111111111101011;
    assign weights1[9][683] = 16'b1111111111111110;
    assign weights1[9][684] = 16'b1111111111111001;
    assign weights1[9][685] = 16'b0000000000001000;
    assign weights1[9][686] = 16'b1111111111100001;
    assign weights1[9][687] = 16'b0000000000000111;
    assign weights1[9][688] = 16'b1111111111111010;
    assign weights1[9][689] = 16'b0000000000001001;
    assign weights1[9][690] = 16'b1111111111110011;
    assign weights1[9][691] = 16'b1111111111011111;
    assign weights1[9][692] = 16'b1111111111110000;
    assign weights1[9][693] = 16'b1111111111110101;
    assign weights1[9][694] = 16'b1111111111110010;
    assign weights1[9][695] = 16'b1111111111101101;
    assign weights1[9][696] = 16'b1111111111111001;
    assign weights1[9][697] = 16'b0000000000000110;
    assign weights1[9][698] = 16'b0000000000000111;
    assign weights1[9][699] = 16'b0000000000000010;
    assign weights1[9][700] = 16'b1111111111111100;
    assign weights1[9][701] = 16'b0000000000000011;
    assign weights1[9][702] = 16'b1111111111111001;
    assign weights1[9][703] = 16'b1111111111100001;
    assign weights1[9][704] = 16'b1111111111010000;
    assign weights1[9][705] = 16'b1111111111010110;
    assign weights1[9][706] = 16'b1111111111001101;
    assign weights1[9][707] = 16'b1111111111001110;
    assign weights1[9][708] = 16'b1111111111000101;
    assign weights1[9][709] = 16'b1111111111001011;
    assign weights1[9][710] = 16'b1111111111001011;
    assign weights1[9][711] = 16'b1111111111010110;
    assign weights1[9][712] = 16'b1111111111011111;
    assign weights1[9][713] = 16'b1111111111011000;
    assign weights1[9][714] = 16'b1111111111011000;
    assign weights1[9][715] = 16'b1111111111011101;
    assign weights1[9][716] = 16'b1111111111011010;
    assign weights1[9][717] = 16'b1111111111010111;
    assign weights1[9][718] = 16'b1111111111100101;
    assign weights1[9][719] = 16'b1111111111100100;
    assign weights1[9][720] = 16'b1111111111011000;
    assign weights1[9][721] = 16'b1111111111101000;
    assign weights1[9][722] = 16'b1111111111011110;
    assign weights1[9][723] = 16'b1111111111100011;
    assign weights1[9][724] = 16'b1111111111111000;
    assign weights1[9][725] = 16'b1111111111111111;
    assign weights1[9][726] = 16'b1111111111111110;
    assign weights1[9][727] = 16'b0000000000000000;
    assign weights1[9][728] = 16'b1111111111111110;
    assign weights1[9][729] = 16'b0000000000000000;
    assign weights1[9][730] = 16'b1111111111111011;
    assign weights1[9][731] = 16'b1111111111101110;
    assign weights1[9][732] = 16'b1111111111101110;
    assign weights1[9][733] = 16'b1111111111101011;
    assign weights1[9][734] = 16'b1111111111110100;
    assign weights1[9][735] = 16'b1111111111101100;
    assign weights1[9][736] = 16'b1111111111100011;
    assign weights1[9][737] = 16'b1111111111011100;
    assign weights1[9][738] = 16'b1111111111001000;
    assign weights1[9][739] = 16'b1111111111011101;
    assign weights1[9][740] = 16'b1111111111100111;
    assign weights1[9][741] = 16'b1111111111011011;
    assign weights1[9][742] = 16'b1111111111010011;
    assign weights1[9][743] = 16'b1111111111001011;
    assign weights1[9][744] = 16'b1111111111010111;
    assign weights1[9][745] = 16'b1111111111100011;
    assign weights1[9][746] = 16'b1111111111100010;
    assign weights1[9][747] = 16'b1111111111110001;
    assign weights1[9][748] = 16'b1111111111100011;
    assign weights1[9][749] = 16'b1111111111011111;
    assign weights1[9][750] = 16'b1111111111011111;
    assign weights1[9][751] = 16'b1111111111101110;
    assign weights1[9][752] = 16'b1111111111111100;
    assign weights1[9][753] = 16'b0000000000000010;
    assign weights1[9][754] = 16'b1111111111111110;
    assign weights1[9][755] = 16'b0000000000000000;
    assign weights1[9][756] = 16'b0000000000000010;
    assign weights1[9][757] = 16'b0000000000000011;
    assign weights1[9][758] = 16'b0000000000000011;
    assign weights1[9][759] = 16'b1111111111111110;
    assign weights1[9][760] = 16'b1111111111111010;
    assign weights1[9][761] = 16'b1111111111111111;
    assign weights1[9][762] = 16'b1111111111111100;
    assign weights1[9][763] = 16'b1111111111110110;
    assign weights1[9][764] = 16'b1111111111100001;
    assign weights1[9][765] = 16'b1111111111011111;
    assign weights1[9][766] = 16'b1111111111011111;
    assign weights1[9][767] = 16'b1111111111101110;
    assign weights1[9][768] = 16'b1111111111011110;
    assign weights1[9][769] = 16'b1111111111100101;
    assign weights1[9][770] = 16'b1111111111100000;
    assign weights1[9][771] = 16'b1111111111110001;
    assign weights1[9][772] = 16'b1111111111011111;
    assign weights1[9][773] = 16'b1111111111101001;
    assign weights1[9][774] = 16'b1111111111100000;
    assign weights1[9][775] = 16'b1111111111011011;
    assign weights1[9][776] = 16'b1111111111011000;
    assign weights1[9][777] = 16'b1111111111100011;
    assign weights1[9][778] = 16'b1111111111100100;
    assign weights1[9][779] = 16'b1111111111110001;
    assign weights1[9][780] = 16'b1111111111110011;
    assign weights1[9][781] = 16'b1111111111111101;
    assign weights1[9][782] = 16'b0000000000000001;
    assign weights1[9][783] = 16'b0000000000000010;
    assign weights1[10][0] = 16'b0000000000000000;
    assign weights1[10][1] = 16'b0000000000000000;
    assign weights1[10][2] = 16'b0000000000000000;
    assign weights1[10][3] = 16'b0000000000000000;
    assign weights1[10][4] = 16'b1111111111111110;
    assign weights1[10][5] = 16'b1111111111111111;
    assign weights1[10][6] = 16'b1111111111111111;
    assign weights1[10][7] = 16'b0000000000000001;
    assign weights1[10][8] = 16'b0000000000001011;
    assign weights1[10][9] = 16'b0000000000001011;
    assign weights1[10][10] = 16'b0000000000010101;
    assign weights1[10][11] = 16'b0000000000010001;
    assign weights1[10][12] = 16'b0000000000011111;
    assign weights1[10][13] = 16'b0000000000100110;
    assign weights1[10][14] = 16'b0000000000101010;
    assign weights1[10][15] = 16'b0000000000011010;
    assign weights1[10][16] = 16'b0000000000100001;
    assign weights1[10][17] = 16'b0000000000010001;
    assign weights1[10][18] = 16'b0000000000000011;
    assign weights1[10][19] = 16'b0000000000011111;
    assign weights1[10][20] = 16'b0000000000010100;
    assign weights1[10][21] = 16'b0000000000000110;
    assign weights1[10][22] = 16'b0000000000001111;
    assign weights1[10][23] = 16'b0000000000011011;
    assign weights1[10][24] = 16'b0000000000001101;
    assign weights1[10][25] = 16'b0000000000000101;
    assign weights1[10][26] = 16'b0000000000000010;
    assign weights1[10][27] = 16'b0000000000000000;
    assign weights1[10][28] = 16'b0000000000000000;
    assign weights1[10][29] = 16'b0000000000000000;
    assign weights1[10][30] = 16'b1111111111111111;
    assign weights1[10][31] = 16'b1111111111111011;
    assign weights1[10][32] = 16'b1111111111111010;
    assign weights1[10][33] = 16'b1111111111111111;
    assign weights1[10][34] = 16'b0000000000001001;
    assign weights1[10][35] = 16'b0000000000000100;
    assign weights1[10][36] = 16'b1111111111111010;
    assign weights1[10][37] = 16'b0000000000000011;
    assign weights1[10][38] = 16'b0000000000001000;
    assign weights1[10][39] = 16'b0000000000100001;
    assign weights1[10][40] = 16'b0000000000100010;
    assign weights1[10][41] = 16'b0000000000011010;
    assign weights1[10][42] = 16'b0000000000101100;
    assign weights1[10][43] = 16'b0000000000011010;
    assign weights1[10][44] = 16'b0000000000010010;
    assign weights1[10][45] = 16'b0000000000010100;
    assign weights1[10][46] = 16'b0000000000011101;
    assign weights1[10][47] = 16'b0000000000001000;
    assign weights1[10][48] = 16'b0000000000011110;
    assign weights1[10][49] = 16'b0000000000010000;
    assign weights1[10][50] = 16'b0000000000011100;
    assign weights1[10][51] = 16'b0000000000000111;
    assign weights1[10][52] = 16'b0000000000000010;
    assign weights1[10][53] = 16'b0000000000001110;
    assign weights1[10][54] = 16'b0000000000001010;
    assign weights1[10][55] = 16'b0000000000000011;
    assign weights1[10][56] = 16'b0000000000000000;
    assign weights1[10][57] = 16'b0000000000000001;
    assign weights1[10][58] = 16'b1111111111111110;
    assign weights1[10][59] = 16'b1111111111111100;
    assign weights1[10][60] = 16'b1111111111111001;
    assign weights1[10][61] = 16'b1111111111111101;
    assign weights1[10][62] = 16'b0000000000001010;
    assign weights1[10][63] = 16'b0000000000000100;
    assign weights1[10][64] = 16'b1111111111111101;
    assign weights1[10][65] = 16'b0000000000000001;
    assign weights1[10][66] = 16'b0000000000010011;
    assign weights1[10][67] = 16'b0000000000010100;
    assign weights1[10][68] = 16'b0000000000011100;
    assign weights1[10][69] = 16'b0000000000100101;
    assign weights1[10][70] = 16'b0000000000100010;
    assign weights1[10][71] = 16'b0000000000011010;
    assign weights1[10][72] = 16'b0000000000011100;
    assign weights1[10][73] = 16'b0000000000001100;
    assign weights1[10][74] = 16'b1111111111111111;
    assign weights1[10][75] = 16'b0000000000001100;
    assign weights1[10][76] = 16'b0000000000010000;
    assign weights1[10][77] = 16'b0000000000001101;
    assign weights1[10][78] = 16'b0000000000000111;
    assign weights1[10][79] = 16'b0000000000000101;
    assign weights1[10][80] = 16'b1111111111111110;
    assign weights1[10][81] = 16'b0000000000010000;
    assign weights1[10][82] = 16'b0000000000001000;
    assign weights1[10][83] = 16'b0000000000010101;
    assign weights1[10][84] = 16'b0000000000000001;
    assign weights1[10][85] = 16'b1111111111111111;
    assign weights1[10][86] = 16'b1111111111111100;
    assign weights1[10][87] = 16'b1111111111110101;
    assign weights1[10][88] = 16'b1111111111110110;
    assign weights1[10][89] = 16'b1111111111111100;
    assign weights1[10][90] = 16'b0000000000000101;
    assign weights1[10][91] = 16'b0000000000000010;
    assign weights1[10][92] = 16'b1111111111111010;
    assign weights1[10][93] = 16'b0000000000000011;
    assign weights1[10][94] = 16'b0000000000000010;
    assign weights1[10][95] = 16'b1111111111111001;
    assign weights1[10][96] = 16'b0000000000011011;
    assign weights1[10][97] = 16'b0000000000010110;
    assign weights1[10][98] = 16'b0000000000010110;
    assign weights1[10][99] = 16'b0000000000010101;
    assign weights1[10][100] = 16'b0000000000010011;
    assign weights1[10][101] = 16'b0000000000010011;
    assign weights1[10][102] = 16'b0000000000011010;
    assign weights1[10][103] = 16'b0000000000010001;
    assign weights1[10][104] = 16'b0000000000010111;
    assign weights1[10][105] = 16'b1111111111111001;
    assign weights1[10][106] = 16'b0000000000000010;
    assign weights1[10][107] = 16'b0000000000001000;
    assign weights1[10][108] = 16'b0000000000001110;
    assign weights1[10][109] = 16'b0000000000011000;
    assign weights1[10][110] = 16'b0000000000011011;
    assign weights1[10][111] = 16'b0000000000011100;
    assign weights1[10][112] = 16'b0000000000000000;
    assign weights1[10][113] = 16'b1111111111111101;
    assign weights1[10][114] = 16'b1111111111110111;
    assign weights1[10][115] = 16'b1111111111110000;
    assign weights1[10][116] = 16'b1111111111101100;
    assign weights1[10][117] = 16'b1111111111110000;
    assign weights1[10][118] = 16'b1111111111110000;
    assign weights1[10][119] = 16'b1111111111101100;
    assign weights1[10][120] = 16'b1111111111110000;
    assign weights1[10][121] = 16'b1111111111110110;
    assign weights1[10][122] = 16'b1111111111110001;
    assign weights1[10][123] = 16'b1111111111110000;
    assign weights1[10][124] = 16'b0000000000000001;
    assign weights1[10][125] = 16'b0000000000000011;
    assign weights1[10][126] = 16'b0000000000010100;
    assign weights1[10][127] = 16'b0000000000010110;
    assign weights1[10][128] = 16'b0000000000001011;
    assign weights1[10][129] = 16'b0000000000011001;
    assign weights1[10][130] = 16'b0000000000011000;
    assign weights1[10][131] = 16'b0000000000010000;
    assign weights1[10][132] = 16'b0000000000001111;
    assign weights1[10][133] = 16'b0000000000010101;
    assign weights1[10][134] = 16'b0000000000000111;
    assign weights1[10][135] = 16'b0000000000010010;
    assign weights1[10][136] = 16'b0000000000010011;
    assign weights1[10][137] = 16'b0000000000100010;
    assign weights1[10][138] = 16'b0000000000100100;
    assign weights1[10][139] = 16'b0000000000011000;
    assign weights1[10][140] = 16'b0000000000000000;
    assign weights1[10][141] = 16'b1111111111111101;
    assign weights1[10][142] = 16'b1111111111110001;
    assign weights1[10][143] = 16'b1111111111101011;
    assign weights1[10][144] = 16'b1111111111101110;
    assign weights1[10][145] = 16'b1111111111110000;
    assign weights1[10][146] = 16'b1111111111100000;
    assign weights1[10][147] = 16'b1111111111011001;
    assign weights1[10][148] = 16'b1111111111100010;
    assign weights1[10][149] = 16'b1111111111110011;
    assign weights1[10][150] = 16'b1111111111110100;
    assign weights1[10][151] = 16'b0000000000001011;
    assign weights1[10][152] = 16'b0000000000000000;
    assign weights1[10][153] = 16'b1111111111101000;
    assign weights1[10][154] = 16'b0000000000011101;
    assign weights1[10][155] = 16'b0000000000100111;
    assign weights1[10][156] = 16'b0000000000000001;
    assign weights1[10][157] = 16'b0000000000011001;
    assign weights1[10][158] = 16'b0000000000001111;
    assign weights1[10][159] = 16'b0000000000010010;
    assign weights1[10][160] = 16'b0000000000010011;
    assign weights1[10][161] = 16'b0000000000001010;
    assign weights1[10][162] = 16'b0000000000010011;
    assign weights1[10][163] = 16'b0000000000010110;
    assign weights1[10][164] = 16'b0000000000000110;
    assign weights1[10][165] = 16'b0000000000011011;
    assign weights1[10][166] = 16'b0000000000011100;
    assign weights1[10][167] = 16'b0000000000100000;
    assign weights1[10][168] = 16'b0000000000000000;
    assign weights1[10][169] = 16'b1111111111111011;
    assign weights1[10][170] = 16'b1111111111101010;
    assign weights1[10][171] = 16'b1111111111101000;
    assign weights1[10][172] = 16'b1111111111100100;
    assign weights1[10][173] = 16'b1111111111011101;
    assign weights1[10][174] = 16'b1111111111011010;
    assign weights1[10][175] = 16'b1111111111110100;
    assign weights1[10][176] = 16'b1111111111101101;
    assign weights1[10][177] = 16'b1111111111111000;
    assign weights1[10][178] = 16'b1111111111110011;
    assign weights1[10][179] = 16'b1111111111111011;
    assign weights1[10][180] = 16'b0000000000000110;
    assign weights1[10][181] = 16'b0000000000001001;
    assign weights1[10][182] = 16'b0000000000010010;
    assign weights1[10][183] = 16'b0000000000010101;
    assign weights1[10][184] = 16'b0000000000000100;
    assign weights1[10][185] = 16'b0000000000010000;
    assign weights1[10][186] = 16'b1111111111111010;
    assign weights1[10][187] = 16'b1111111111110100;
    assign weights1[10][188] = 16'b0000000000010001;
    assign weights1[10][189] = 16'b0000000000000101;
    assign weights1[10][190] = 16'b0000000000001000;
    assign weights1[10][191] = 16'b0000000000001011;
    assign weights1[10][192] = 16'b0000000000001010;
    assign weights1[10][193] = 16'b0000000000001100;
    assign weights1[10][194] = 16'b0000000000001101;
    assign weights1[10][195] = 16'b0000000000010101;
    assign weights1[10][196] = 16'b1111111111111100;
    assign weights1[10][197] = 16'b1111111111110010;
    assign weights1[10][198] = 16'b1111111111101000;
    assign weights1[10][199] = 16'b1111111111100010;
    assign weights1[10][200] = 16'b1111111111011101;
    assign weights1[10][201] = 16'b1111111111011000;
    assign weights1[10][202] = 16'b1111111111101010;
    assign weights1[10][203] = 16'b1111111111101010;
    assign weights1[10][204] = 16'b1111111111011101;
    assign weights1[10][205] = 16'b1111111111101000;
    assign weights1[10][206] = 16'b1111111111110011;
    assign weights1[10][207] = 16'b1111111111101110;
    assign weights1[10][208] = 16'b0000000000000110;
    assign weights1[10][209] = 16'b0000000000000111;
    assign weights1[10][210] = 16'b0000000000001001;
    assign weights1[10][211] = 16'b0000000000011001;
    assign weights1[10][212] = 16'b0000000000000101;
    assign weights1[10][213] = 16'b0000000000010000;
    assign weights1[10][214] = 16'b0000000000001111;
    assign weights1[10][215] = 16'b0000000000011110;
    assign weights1[10][216] = 16'b0000000000000111;
    assign weights1[10][217] = 16'b0000000000000110;
    assign weights1[10][218] = 16'b1111111111111011;
    assign weights1[10][219] = 16'b0000000000000110;
    assign weights1[10][220] = 16'b0000000000000111;
    assign weights1[10][221] = 16'b0000000000001000;
    assign weights1[10][222] = 16'b0000000000000100;
    assign weights1[10][223] = 16'b0000000000010111;
    assign weights1[10][224] = 16'b1111111111111110;
    assign weights1[10][225] = 16'b1111111111101101;
    assign weights1[10][226] = 16'b1111111111100110;
    assign weights1[10][227] = 16'b1111111111010010;
    assign weights1[10][228] = 16'b1111111111010010;
    assign weights1[10][229] = 16'b1111111111001011;
    assign weights1[10][230] = 16'b1111111111010101;
    assign weights1[10][231] = 16'b1111111111101111;
    assign weights1[10][232] = 16'b1111111111011011;
    assign weights1[10][233] = 16'b1111111111110001;
    assign weights1[10][234] = 16'b0000000000010001;
    assign weights1[10][235] = 16'b0000000000010000;
    assign weights1[10][236] = 16'b0000000000001001;
    assign weights1[10][237] = 16'b0000000000100000;
    assign weights1[10][238] = 16'b0000000000101001;
    assign weights1[10][239] = 16'b0000000000101100;
    assign weights1[10][240] = 16'b0000000000100101;
    assign weights1[10][241] = 16'b0000000000101100;
    assign weights1[10][242] = 16'b0000000000011010;
    assign weights1[10][243] = 16'b0000000000001100;
    assign weights1[10][244] = 16'b0000000000000110;
    assign weights1[10][245] = 16'b0000000000000111;
    assign weights1[10][246] = 16'b1111111111111101;
    assign weights1[10][247] = 16'b0000000000000101;
    assign weights1[10][248] = 16'b0000000000001001;
    assign weights1[10][249] = 16'b0000000000001110;
    assign weights1[10][250] = 16'b0000000000001010;
    assign weights1[10][251] = 16'b0000000000010000;
    assign weights1[10][252] = 16'b1111111111111001;
    assign weights1[10][253] = 16'b1111111111101110;
    assign weights1[10][254] = 16'b1111111111100010;
    assign weights1[10][255] = 16'b1111111111100000;
    assign weights1[10][256] = 16'b1111111111001101;
    assign weights1[10][257] = 16'b1111111111000001;
    assign weights1[10][258] = 16'b1111111110111101;
    assign weights1[10][259] = 16'b1111111110111101;
    assign weights1[10][260] = 16'b1111111111010111;
    assign weights1[10][261] = 16'b1111111111100111;
    assign weights1[10][262] = 16'b1111111111110111;
    assign weights1[10][263] = 16'b1111111111110111;
    assign weights1[10][264] = 16'b0000000000010001;
    assign weights1[10][265] = 16'b0000000000000111;
    assign weights1[10][266] = 16'b0000000000111100;
    assign weights1[10][267] = 16'b0000000001000110;
    assign weights1[10][268] = 16'b0000000001010000;
    assign weights1[10][269] = 16'b0000000000110001;
    assign weights1[10][270] = 16'b0000000000101101;
    assign weights1[10][271] = 16'b0000000000100001;
    assign weights1[10][272] = 16'b0000000000010110;
    assign weights1[10][273] = 16'b0000000000001101;
    assign weights1[10][274] = 16'b0000000000001111;
    assign weights1[10][275] = 16'b0000000000001101;
    assign weights1[10][276] = 16'b1111111111111101;
    assign weights1[10][277] = 16'b1111111111111111;
    assign weights1[10][278] = 16'b0000000000001101;
    assign weights1[10][279] = 16'b0000000000010001;
    assign weights1[10][280] = 16'b1111111111111010;
    assign weights1[10][281] = 16'b1111111111101000;
    assign weights1[10][282] = 16'b1111111111011110;
    assign weights1[10][283] = 16'b1111111111100100;
    assign weights1[10][284] = 16'b1111111111010001;
    assign weights1[10][285] = 16'b1111111111000001;
    assign weights1[10][286] = 16'b1111111110101011;
    assign weights1[10][287] = 16'b1111111110111000;
    assign weights1[10][288] = 16'b1111111110101110;
    assign weights1[10][289] = 16'b1111111110110101;
    assign weights1[10][290] = 16'b1111111111001011;
    assign weights1[10][291] = 16'b1111111111010111;
    assign weights1[10][292] = 16'b1111111111110101;
    assign weights1[10][293] = 16'b0000000000001111;
    assign weights1[10][294] = 16'b0000000000001110;
    assign weights1[10][295] = 16'b0000000000010110;
    assign weights1[10][296] = 16'b0000000001000000;
    assign weights1[10][297] = 16'b0000000000101110;
    assign weights1[10][298] = 16'b0000000000010111;
    assign weights1[10][299] = 16'b0000000000100101;
    assign weights1[10][300] = 16'b0000000000011100;
    assign weights1[10][301] = 16'b0000000000011001;
    assign weights1[10][302] = 16'b1111111111111100;
    assign weights1[10][303] = 16'b0000000000010111;
    assign weights1[10][304] = 16'b0000000000000011;
    assign weights1[10][305] = 16'b0000000000010001;
    assign weights1[10][306] = 16'b0000000000010101;
    assign weights1[10][307] = 16'b0000000000011010;
    assign weights1[10][308] = 16'b1111111111111101;
    assign weights1[10][309] = 16'b1111111111101111;
    assign weights1[10][310] = 16'b1111111111101101;
    assign weights1[10][311] = 16'b1111111111110011;
    assign weights1[10][312] = 16'b1111111111001011;
    assign weights1[10][313] = 16'b1111111111010011;
    assign weights1[10][314] = 16'b1111111111000110;
    assign weights1[10][315] = 16'b1111111110101101;
    assign weights1[10][316] = 16'b1111111110001110;
    assign weights1[10][317] = 16'b1111111110001000;
    assign weights1[10][318] = 16'b1111111110100110;
    assign weights1[10][319] = 16'b1111111111000111;
    assign weights1[10][320] = 16'b1111111111100000;
    assign weights1[10][321] = 16'b1111111111100101;
    assign weights1[10][322] = 16'b0000000000000111;
    assign weights1[10][323] = 16'b0000000000101011;
    assign weights1[10][324] = 16'b0000000000101111;
    assign weights1[10][325] = 16'b0000000000100010;
    assign weights1[10][326] = 16'b0000000000010000;
    assign weights1[10][327] = 16'b0000000000001010;
    assign weights1[10][328] = 16'b0000000000001110;
    assign weights1[10][329] = 16'b0000000000001110;
    assign weights1[10][330] = 16'b0000000000010110;
    assign weights1[10][331] = 16'b0000000000011100;
    assign weights1[10][332] = 16'b0000000000001010;
    assign weights1[10][333] = 16'b1111111111111001;
    assign weights1[10][334] = 16'b0000000000010000;
    assign weights1[10][335] = 16'b0000000000010111;
    assign weights1[10][336] = 16'b1111111111111010;
    assign weights1[10][337] = 16'b1111111111110101;
    assign weights1[10][338] = 16'b1111111111111010;
    assign weights1[10][339] = 16'b0000000000000001;
    assign weights1[10][340] = 16'b1111111111110011;
    assign weights1[10][341] = 16'b1111111111100100;
    assign weights1[10][342] = 16'b1111111111011111;
    assign weights1[10][343] = 16'b1111111110111111;
    assign weights1[10][344] = 16'b1111111110011011;
    assign weights1[10][345] = 16'b1111111110000001;
    assign weights1[10][346] = 16'b1111111110000110;
    assign weights1[10][347] = 16'b1111111101111110;
    assign weights1[10][348] = 16'b1111111110100001;
    assign weights1[10][349] = 16'b1111111111000111;
    assign weights1[10][350] = 16'b1111111111100111;
    assign weights1[10][351] = 16'b0000000000011001;
    assign weights1[10][352] = 16'b0000000000111101;
    assign weights1[10][353] = 16'b0000000000010000;
    assign weights1[10][354] = 16'b0000000000010001;
    assign weights1[10][355] = 16'b0000000000010011;
    assign weights1[10][356] = 16'b0000000000001101;
    assign weights1[10][357] = 16'b0000000000000011;
    assign weights1[10][358] = 16'b0000000000001010;
    assign weights1[10][359] = 16'b1111111111111111;
    assign weights1[10][360] = 16'b1111111111111000;
    assign weights1[10][361] = 16'b1111111111111011;
    assign weights1[10][362] = 16'b0000000000000101;
    assign weights1[10][363] = 16'b0000000000000000;
    assign weights1[10][364] = 16'b0000000000000100;
    assign weights1[10][365] = 16'b1111111111111111;
    assign weights1[10][366] = 16'b1111111111111011;
    assign weights1[10][367] = 16'b0000000000001001;
    assign weights1[10][368] = 16'b0000000000001000;
    assign weights1[10][369] = 16'b0000000000001011;
    assign weights1[10][370] = 16'b0000000000000000;
    assign weights1[10][371] = 16'b0000000000000000;
    assign weights1[10][372] = 16'b1111111111011111;
    assign weights1[10][373] = 16'b1111111110110001;
    assign weights1[10][374] = 16'b1111111110011000;
    assign weights1[10][375] = 16'b1111111110010000;
    assign weights1[10][376] = 16'b1111111101110011;
    assign weights1[10][377] = 16'b1111111110010000;
    assign weights1[10][378] = 16'b1111111110110001;
    assign weights1[10][379] = 16'b0000000000011100;
    assign weights1[10][380] = 16'b0000000000111101;
    assign weights1[10][381] = 16'b0000000000110100;
    assign weights1[10][382] = 16'b0000000000001001;
    assign weights1[10][383] = 16'b0000000000000111;
    assign weights1[10][384] = 16'b0000000000100000;
    assign weights1[10][385] = 16'b1111111111111000;
    assign weights1[10][386] = 16'b1111111111111110;
    assign weights1[10][387] = 16'b1111111111110111;
    assign weights1[10][388] = 16'b1111111111111101;
    assign weights1[10][389] = 16'b1111111111110111;
    assign weights1[10][390] = 16'b1111111111110010;
    assign weights1[10][391] = 16'b1111111111110000;
    assign weights1[10][392] = 16'b0000000000001001;
    assign weights1[10][393] = 16'b0000000000000011;
    assign weights1[10][394] = 16'b0000000000001010;
    assign weights1[10][395] = 16'b0000000000010010;
    assign weights1[10][396] = 16'b0000000000011011;
    assign weights1[10][397] = 16'b0000000000010110;
    assign weights1[10][398] = 16'b0000000000011000;
    assign weights1[10][399] = 16'b0000000000101010;
    assign weights1[10][400] = 16'b0000000000001101;
    assign weights1[10][401] = 16'b0000000000001000;
    assign weights1[10][402] = 16'b1111111111100100;
    assign weights1[10][403] = 16'b1111111110111011;
    assign weights1[10][404] = 16'b1111111110001110;
    assign weights1[10][405] = 16'b1111111110000110;
    assign weights1[10][406] = 16'b1111111110001111;
    assign weights1[10][407] = 16'b1111111111010001;
    assign weights1[10][408] = 16'b0000000000100011;
    assign weights1[10][409] = 16'b0000000000010000;
    assign weights1[10][410] = 16'b0000000000011100;
    assign weights1[10][411] = 16'b0000000000001110;
    assign weights1[10][412] = 16'b0000000000000110;
    assign weights1[10][413] = 16'b0000000000000101;
    assign weights1[10][414] = 16'b0000000000001000;
    assign weights1[10][415] = 16'b0000000000000111;
    assign weights1[10][416] = 16'b0000000000000011;
    assign weights1[10][417] = 16'b1111111111111001;
    assign weights1[10][418] = 16'b1111111111101101;
    assign weights1[10][419] = 16'b1111111111100001;
    assign weights1[10][420] = 16'b0000000000000101;
    assign weights1[10][421] = 16'b0000000000000111;
    assign weights1[10][422] = 16'b0000000000001110;
    assign weights1[10][423] = 16'b0000000000001001;
    assign weights1[10][424] = 16'b0000000000101000;
    assign weights1[10][425] = 16'b0000000000100011;
    assign weights1[10][426] = 16'b0000000000101101;
    assign weights1[10][427] = 16'b0000000000111101;
    assign weights1[10][428] = 16'b0000000000110110;
    assign weights1[10][429] = 16'b0000000000111000;
    assign weights1[10][430] = 16'b0000000000010001;
    assign weights1[10][431] = 16'b1111111111111001;
    assign weights1[10][432] = 16'b1111111111011011;
    assign weights1[10][433] = 16'b1111111110010100;
    assign weights1[10][434] = 16'b1111111110000100;
    assign weights1[10][435] = 16'b1111111110111111;
    assign weights1[10][436] = 16'b0000000000000000;
    assign weights1[10][437] = 16'b0000000000010110;
    assign weights1[10][438] = 16'b0000000000011100;
    assign weights1[10][439] = 16'b0000000000000001;
    assign weights1[10][440] = 16'b0000000000000010;
    assign weights1[10][441] = 16'b0000000000100001;
    assign weights1[10][442] = 16'b0000000000010101;
    assign weights1[10][443] = 16'b1111111111110101;
    assign weights1[10][444] = 16'b1111111111110101;
    assign weights1[10][445] = 16'b0000000000000010;
    assign weights1[10][446] = 16'b1111111111100111;
    assign weights1[10][447] = 16'b1111111111101010;
    assign weights1[10][448] = 16'b1111111111111111;
    assign weights1[10][449] = 16'b1111111111111111;
    assign weights1[10][450] = 16'b0000000000001011;
    assign weights1[10][451] = 16'b0000000000000011;
    assign weights1[10][452] = 16'b0000000000100111;
    assign weights1[10][453] = 16'b1111111111110000;
    assign weights1[10][454] = 16'b0000000000001100;
    assign weights1[10][455] = 16'b1111111111110100;
    assign weights1[10][456] = 16'b0000000000001011;
    assign weights1[10][457] = 16'b0000000000011111;
    assign weights1[10][458] = 16'b0000000000001100;
    assign weights1[10][459] = 16'b0000000000001011;
    assign weights1[10][460] = 16'b1111111111111011;
    assign weights1[10][461] = 16'b1111111111000100;
    assign weights1[10][462] = 16'b1111111110011000;
    assign weights1[10][463] = 16'b1111111110110001;
    assign weights1[10][464] = 16'b1111111111011111;
    assign weights1[10][465] = 16'b0000000000011010;
    assign weights1[10][466] = 16'b0000000000001110;
    assign weights1[10][467] = 16'b1111111111111101;
    assign weights1[10][468] = 16'b0000000000010010;
    assign weights1[10][469] = 16'b1111111111111101;
    assign weights1[10][470] = 16'b0000000000011000;
    assign weights1[10][471] = 16'b0000000000001101;
    assign weights1[10][472] = 16'b1111111111111000;
    assign weights1[10][473] = 16'b1111111111111111;
    assign weights1[10][474] = 16'b1111111111101111;
    assign weights1[10][475] = 16'b1111111111100100;
    assign weights1[10][476] = 16'b1111111111111001;
    assign weights1[10][477] = 16'b1111111111101101;
    assign weights1[10][478] = 16'b1111111111101100;
    assign weights1[10][479] = 16'b1111111111100111;
    assign weights1[10][480] = 16'b0000000000001011;
    assign weights1[10][481] = 16'b0000000000000100;
    assign weights1[10][482] = 16'b1111111111100110;
    assign weights1[10][483] = 16'b1111111111111110;
    assign weights1[10][484] = 16'b0000000000000001;
    assign weights1[10][485] = 16'b0000000000000000;
    assign weights1[10][486] = 16'b1111111111111000;
    assign weights1[10][487] = 16'b0000000000010000;
    assign weights1[10][488] = 16'b1111111111111111;
    assign weights1[10][489] = 16'b1111111111100000;
    assign weights1[10][490] = 16'b1111111110110100;
    assign weights1[10][491] = 16'b1111111110111101;
    assign weights1[10][492] = 16'b1111111111011110;
    assign weights1[10][493] = 16'b0000000000000011;
    assign weights1[10][494] = 16'b0000000000001010;
    assign weights1[10][495] = 16'b0000000000010000;
    assign weights1[10][496] = 16'b0000000000001100;
    assign weights1[10][497] = 16'b0000000000000101;
    assign weights1[10][498] = 16'b0000000000000000;
    assign weights1[10][499] = 16'b0000000000000100;
    assign weights1[10][500] = 16'b0000000000010000;
    assign weights1[10][501] = 16'b1111111111110111;
    assign weights1[10][502] = 16'b1111111111100111;
    assign weights1[10][503] = 16'b1111111111101000;
    assign weights1[10][504] = 16'b1111111111111000;
    assign weights1[10][505] = 16'b1111111111110001;
    assign weights1[10][506] = 16'b1111111111100100;
    assign weights1[10][507] = 16'b1111111111011111;
    assign weights1[10][508] = 16'b1111111111110011;
    assign weights1[10][509] = 16'b1111111111010110;
    assign weights1[10][510] = 16'b1111111111100110;
    assign weights1[10][511] = 16'b1111111111111010;
    assign weights1[10][512] = 16'b1111111111101111;
    assign weights1[10][513] = 16'b1111111111111101;
    assign weights1[10][514] = 16'b1111111111101000;
    assign weights1[10][515] = 16'b1111111111111011;
    assign weights1[10][516] = 16'b0000000000001001;
    assign weights1[10][517] = 16'b1111111111110010;
    assign weights1[10][518] = 16'b1111111111100000;
    assign weights1[10][519] = 16'b1111111111001110;
    assign weights1[10][520] = 16'b1111111111010110;
    assign weights1[10][521] = 16'b0000000000000100;
    assign weights1[10][522] = 16'b0000000000000101;
    assign weights1[10][523] = 16'b0000000000001111;
    assign weights1[10][524] = 16'b0000000000010011;
    assign weights1[10][525] = 16'b0000000000010011;
    assign weights1[10][526] = 16'b0000000000001111;
    assign weights1[10][527] = 16'b0000000000011100;
    assign weights1[10][528] = 16'b0000000000010001;
    assign weights1[10][529] = 16'b1111111111110011;
    assign weights1[10][530] = 16'b1111111111101100;
    assign weights1[10][531] = 16'b1111111111011101;
    assign weights1[10][532] = 16'b1111111111111010;
    assign weights1[10][533] = 16'b1111111111110111;
    assign weights1[10][534] = 16'b1111111111101101;
    assign weights1[10][535] = 16'b1111111111101000;
    assign weights1[10][536] = 16'b1111111111100110;
    assign weights1[10][537] = 16'b1111111111011100;
    assign weights1[10][538] = 16'b1111111111110101;
    assign weights1[10][539] = 16'b1111111111111110;
    assign weights1[10][540] = 16'b1111111111110001;
    assign weights1[10][541] = 16'b0000000000000001;
    assign weights1[10][542] = 16'b1111111111110001;
    assign weights1[10][543] = 16'b1111111111110100;
    assign weights1[10][544] = 16'b1111111111110110;
    assign weights1[10][545] = 16'b1111111111110100;
    assign weights1[10][546] = 16'b1111111111110100;
    assign weights1[10][547] = 16'b1111111111101111;
    assign weights1[10][548] = 16'b1111111111110111;
    assign weights1[10][549] = 16'b1111111111101100;
    assign weights1[10][550] = 16'b1111111111110101;
    assign weights1[10][551] = 16'b0000000000001110;
    assign weights1[10][552] = 16'b0000000000010100;
    assign weights1[10][553] = 16'b0000000000010110;
    assign weights1[10][554] = 16'b0000000000011000;
    assign weights1[10][555] = 16'b0000000000010000;
    assign weights1[10][556] = 16'b0000000000000101;
    assign weights1[10][557] = 16'b1111111111101100;
    assign weights1[10][558] = 16'b1111111111011101;
    assign weights1[10][559] = 16'b1111111111010110;
    assign weights1[10][560] = 16'b1111111111111100;
    assign weights1[10][561] = 16'b1111111111111000;
    assign weights1[10][562] = 16'b1111111111110010;
    assign weights1[10][563] = 16'b1111111111100000;
    assign weights1[10][564] = 16'b1111111111001110;
    assign weights1[10][565] = 16'b1111111111111011;
    assign weights1[10][566] = 16'b1111111111110011;
    assign weights1[10][567] = 16'b1111111111111000;
    assign weights1[10][568] = 16'b1111111111101011;
    assign weights1[10][569] = 16'b1111111111110110;
    assign weights1[10][570] = 16'b1111111111111011;
    assign weights1[10][571] = 16'b1111111111101110;
    assign weights1[10][572] = 16'b1111111111111111;
    assign weights1[10][573] = 16'b1111111111101100;
    assign weights1[10][574] = 16'b1111111111101101;
    assign weights1[10][575] = 16'b1111111111011010;
    assign weights1[10][576] = 16'b1111111111011111;
    assign weights1[10][577] = 16'b1111111111011111;
    assign weights1[10][578] = 16'b1111111111111001;
    assign weights1[10][579] = 16'b0000000000001001;
    assign weights1[10][580] = 16'b0000000000011001;
    assign weights1[10][581] = 16'b1111111111111010;
    assign weights1[10][582] = 16'b0000000000001111;
    assign weights1[10][583] = 16'b0000000000000100;
    assign weights1[10][584] = 16'b1111111111110101;
    assign weights1[10][585] = 16'b1111111111101101;
    assign weights1[10][586] = 16'b1111111111100001;
    assign weights1[10][587] = 16'b1111111111100001;
    assign weights1[10][588] = 16'b1111111111111100;
    assign weights1[10][589] = 16'b1111111111110101;
    assign weights1[10][590] = 16'b1111111111110000;
    assign weights1[10][591] = 16'b1111111111100100;
    assign weights1[10][592] = 16'b1111111111101100;
    assign weights1[10][593] = 16'b1111111111111110;
    assign weights1[10][594] = 16'b1111111111111010;
    assign weights1[10][595] = 16'b1111111111101010;
    assign weights1[10][596] = 16'b1111111111101110;
    assign weights1[10][597] = 16'b1111111111111000;
    assign weights1[10][598] = 16'b1111111111110111;
    assign weights1[10][599] = 16'b0000000000010000;
    assign weights1[10][600] = 16'b1111111111110001;
    assign weights1[10][601] = 16'b1111111111100111;
    assign weights1[10][602] = 16'b1111111111100100;
    assign weights1[10][603] = 16'b1111111111010101;
    assign weights1[10][604] = 16'b1111111111100101;
    assign weights1[10][605] = 16'b1111111111101010;
    assign weights1[10][606] = 16'b1111111111101110;
    assign weights1[10][607] = 16'b0000000000000011;
    assign weights1[10][608] = 16'b0000000000000100;
    assign weights1[10][609] = 16'b0000000000010000;
    assign weights1[10][610] = 16'b0000000000001110;
    assign weights1[10][611] = 16'b0000000000011011;
    assign weights1[10][612] = 16'b1111111111101100;
    assign weights1[10][613] = 16'b1111111111111111;
    assign weights1[10][614] = 16'b1111111111100101;
    assign weights1[10][615] = 16'b1111111111101011;
    assign weights1[10][616] = 16'b1111111111111101;
    assign weights1[10][617] = 16'b1111111111111010;
    assign weights1[10][618] = 16'b1111111111110011;
    assign weights1[10][619] = 16'b1111111111110111;
    assign weights1[10][620] = 16'b0000000000000100;
    assign weights1[10][621] = 16'b1111111111110001;
    assign weights1[10][622] = 16'b1111111111111100;
    assign weights1[10][623] = 16'b1111111111110100;
    assign weights1[10][624] = 16'b1111111111001010;
    assign weights1[10][625] = 16'b0000000000000001;
    assign weights1[10][626] = 16'b1111111111110000;
    assign weights1[10][627] = 16'b0000000000000011;
    assign weights1[10][628] = 16'b1111111111110001;
    assign weights1[10][629] = 16'b1111111111101111;
    assign weights1[10][630] = 16'b0000000000000000;
    assign weights1[10][631] = 16'b1111111111111111;
    assign weights1[10][632] = 16'b1111111111101001;
    assign weights1[10][633] = 16'b1111111111101111;
    assign weights1[10][634] = 16'b1111111111100001;
    assign weights1[10][635] = 16'b1111111111111010;
    assign weights1[10][636] = 16'b0000000000000001;
    assign weights1[10][637] = 16'b0000000000010011;
    assign weights1[10][638] = 16'b0000000000010101;
    assign weights1[10][639] = 16'b0000000000001001;
    assign weights1[10][640] = 16'b1111111111110111;
    assign weights1[10][641] = 16'b1111111111101011;
    assign weights1[10][642] = 16'b1111111111101010;
    assign weights1[10][643] = 16'b1111111111110100;
    assign weights1[10][644] = 16'b0000000000000000;
    assign weights1[10][645] = 16'b1111111111111011;
    assign weights1[10][646] = 16'b1111111111111110;
    assign weights1[10][647] = 16'b0000000000000001;
    assign weights1[10][648] = 16'b0000000000001101;
    assign weights1[10][649] = 16'b1111111111111110;
    assign weights1[10][650] = 16'b1111111111110000;
    assign weights1[10][651] = 16'b1111111111111011;
    assign weights1[10][652] = 16'b1111111111110011;
    assign weights1[10][653] = 16'b0000000000000110;
    assign weights1[10][654] = 16'b1111111111101101;
    assign weights1[10][655] = 16'b1111111111110000;
    assign weights1[10][656] = 16'b1111111111110111;
    assign weights1[10][657] = 16'b1111111111011101;
    assign weights1[10][658] = 16'b1111111111101100;
    assign weights1[10][659] = 16'b1111111111011101;
    assign weights1[10][660] = 16'b1111111111101111;
    assign weights1[10][661] = 16'b0000000000001101;
    assign weights1[10][662] = 16'b1111111111111110;
    assign weights1[10][663] = 16'b0000000000000001;
    assign weights1[10][664] = 16'b0000000000000010;
    assign weights1[10][665] = 16'b0000000000001001;
    assign weights1[10][666] = 16'b0000000000011010;
    assign weights1[10][667] = 16'b1111111111110010;
    assign weights1[10][668] = 16'b1111111111110100;
    assign weights1[10][669] = 16'b1111111111100101;
    assign weights1[10][670] = 16'b1111111111100101;
    assign weights1[10][671] = 16'b1111111111110010;
    assign weights1[10][672] = 16'b0000000000000000;
    assign weights1[10][673] = 16'b1111111111111101;
    assign weights1[10][674] = 16'b1111111111111011;
    assign weights1[10][675] = 16'b1111111111111100;
    assign weights1[10][676] = 16'b1111111111111110;
    assign weights1[10][677] = 16'b1111111111110101;
    assign weights1[10][678] = 16'b1111111111100111;
    assign weights1[10][679] = 16'b1111111111101011;
    assign weights1[10][680] = 16'b1111111111100010;
    assign weights1[10][681] = 16'b1111111111011101;
    assign weights1[10][682] = 16'b1111111111100101;
    assign weights1[10][683] = 16'b1111111111110100;
    assign weights1[10][684] = 16'b1111111111101100;
    assign weights1[10][685] = 16'b1111111111100000;
    assign weights1[10][686] = 16'b0000000000000001;
    assign weights1[10][687] = 16'b1111111111100110;
    assign weights1[10][688] = 16'b0000000000000011;
    assign weights1[10][689] = 16'b0000000000000111;
    assign weights1[10][690] = 16'b0000000000001001;
    assign weights1[10][691] = 16'b0000000000000011;
    assign weights1[10][692] = 16'b0000000000010000;
    assign weights1[10][693] = 16'b0000000000000000;
    assign weights1[10][694] = 16'b0000000000011000;
    assign weights1[10][695] = 16'b1111111111111101;
    assign weights1[10][696] = 16'b1111111111110001;
    assign weights1[10][697] = 16'b1111111111100010;
    assign weights1[10][698] = 16'b1111111111101100;
    assign weights1[10][699] = 16'b1111111111110111;
    assign weights1[10][700] = 16'b0000000000000000;
    assign weights1[10][701] = 16'b1111111111111111;
    assign weights1[10][702] = 16'b1111111111111011;
    assign weights1[10][703] = 16'b1111111111111001;
    assign weights1[10][704] = 16'b1111111111111100;
    assign weights1[10][705] = 16'b1111111111111100;
    assign weights1[10][706] = 16'b1111111111101110;
    assign weights1[10][707] = 16'b1111111111101001;
    assign weights1[10][708] = 16'b1111111111101100;
    assign weights1[10][709] = 16'b1111111111101000;
    assign weights1[10][710] = 16'b1111111111110001;
    assign weights1[10][711] = 16'b1111111111111110;
    assign weights1[10][712] = 16'b1111111111110101;
    assign weights1[10][713] = 16'b1111111111101100;
    assign weights1[10][714] = 16'b1111111111111100;
    assign weights1[10][715] = 16'b1111111111111000;
    assign weights1[10][716] = 16'b1111111111111011;
    assign weights1[10][717] = 16'b1111111111111001;
    assign weights1[10][718] = 16'b1111111111110110;
    assign weights1[10][719] = 16'b1111111111110110;
    assign weights1[10][720] = 16'b0000000000000011;
    assign weights1[10][721] = 16'b0000000000001100;
    assign weights1[10][722] = 16'b0000000000000110;
    assign weights1[10][723] = 16'b1111111111101110;
    assign weights1[10][724] = 16'b1111111111110001;
    assign weights1[10][725] = 16'b1111111111101010;
    assign weights1[10][726] = 16'b1111111111101111;
    assign weights1[10][727] = 16'b1111111111111110;
    assign weights1[10][728] = 16'b0000000000000000;
    assign weights1[10][729] = 16'b0000000000000000;
    assign weights1[10][730] = 16'b1111111111111100;
    assign weights1[10][731] = 16'b1111111111111011;
    assign weights1[10][732] = 16'b1111111111111010;
    assign weights1[10][733] = 16'b1111111111110001;
    assign weights1[10][734] = 16'b1111111111110110;
    assign weights1[10][735] = 16'b1111111111110110;
    assign weights1[10][736] = 16'b1111111111110101;
    assign weights1[10][737] = 16'b1111111111101111;
    assign weights1[10][738] = 16'b1111111111110011;
    assign weights1[10][739] = 16'b1111111111110000;
    assign weights1[10][740] = 16'b1111111111101011;
    assign weights1[10][741] = 16'b1111111111111010;
    assign weights1[10][742] = 16'b1111111111110100;
    assign weights1[10][743] = 16'b1111111111101001;
    assign weights1[10][744] = 16'b1111111111110110;
    assign weights1[10][745] = 16'b1111111111110001;
    assign weights1[10][746] = 16'b1111111111111000;
    assign weights1[10][747] = 16'b1111111111101101;
    assign weights1[10][748] = 16'b1111111111111110;
    assign weights1[10][749] = 16'b0000000000001010;
    assign weights1[10][750] = 16'b0000000000000000;
    assign weights1[10][751] = 16'b1111111111101100;
    assign weights1[10][752] = 16'b1111111111110000;
    assign weights1[10][753] = 16'b1111111111110110;
    assign weights1[10][754] = 16'b1111111111111010;
    assign weights1[10][755] = 16'b1111111111111111;
    assign weights1[10][756] = 16'b0000000000000000;
    assign weights1[10][757] = 16'b1111111111111110;
    assign weights1[10][758] = 16'b1111111111111110;
    assign weights1[10][759] = 16'b1111111111111100;
    assign weights1[10][760] = 16'b1111111111111010;
    assign weights1[10][761] = 16'b1111111111111001;
    assign weights1[10][762] = 16'b1111111111110101;
    assign weights1[10][763] = 16'b1111111111111000;
    assign weights1[10][764] = 16'b1111111111110110;
    assign weights1[10][765] = 16'b1111111111110111;
    assign weights1[10][766] = 16'b1111111111111010;
    assign weights1[10][767] = 16'b1111111111101100;
    assign weights1[10][768] = 16'b1111111111110101;
    assign weights1[10][769] = 16'b1111111111101111;
    assign weights1[10][770] = 16'b1111111111100010;
    assign weights1[10][771] = 16'b1111111111111100;
    assign weights1[10][772] = 16'b1111111111110000;
    assign weights1[10][773] = 16'b1111111111110110;
    assign weights1[10][774] = 16'b0000000000001011;
    assign weights1[10][775] = 16'b0000000000010010;
    assign weights1[10][776] = 16'b0000000000000111;
    assign weights1[10][777] = 16'b0000000000001111;
    assign weights1[10][778] = 16'b0000000000000000;
    assign weights1[10][779] = 16'b1111111111111111;
    assign weights1[10][780] = 16'b1111111111111100;
    assign weights1[10][781] = 16'b1111111111111101;
    assign weights1[10][782] = 16'b1111111111111101;
    assign weights1[10][783] = 16'b1111111111111111;
    assign weights1[11][0] = 16'b0000000000000000;
    assign weights1[11][1] = 16'b0000000000000000;
    assign weights1[11][2] = 16'b0000000000000000;
    assign weights1[11][3] = 16'b1111111111111110;
    assign weights1[11][4] = 16'b0000000000000010;
    assign weights1[11][5] = 16'b0000000000000011;
    assign weights1[11][6] = 16'b1111111111111110;
    assign weights1[11][7] = 16'b1111111111111101;
    assign weights1[11][8] = 16'b1111111111111010;
    assign weights1[11][9] = 16'b1111111111110101;
    assign weights1[11][10] = 16'b1111111111110000;
    assign weights1[11][11] = 16'b1111111111101011;
    assign weights1[11][12] = 16'b0000000000000011;
    assign weights1[11][13] = 16'b1111111111110100;
    assign weights1[11][14] = 16'b1111111111101111;
    assign weights1[11][15] = 16'b1111111111111011;
    assign weights1[11][16] = 16'b1111111111110111;
    assign weights1[11][17] = 16'b0000000000001000;
    assign weights1[11][18] = 16'b0000000000000001;
    assign weights1[11][19] = 16'b0000000000000011;
    assign weights1[11][20] = 16'b0000000000000101;
    assign weights1[11][21] = 16'b1111111111111111;
    assign weights1[11][22] = 16'b1111111111110110;
    assign weights1[11][23] = 16'b1111111111101101;
    assign weights1[11][24] = 16'b1111111111101110;
    assign weights1[11][25] = 16'b1111111111110100;
    assign weights1[11][26] = 16'b1111111111111001;
    assign weights1[11][27] = 16'b1111111111111100;
    assign weights1[11][28] = 16'b0000000000000000;
    assign weights1[11][29] = 16'b0000000000000001;
    assign weights1[11][30] = 16'b0000000000000100;
    assign weights1[11][31] = 16'b0000000000000100;
    assign weights1[11][32] = 16'b0000000000000111;
    assign weights1[11][33] = 16'b0000000000000100;
    assign weights1[11][34] = 16'b1111111111111010;
    assign weights1[11][35] = 16'b1111111111111101;
    assign weights1[11][36] = 16'b0000000000000110;
    assign weights1[11][37] = 16'b1111111111111011;
    assign weights1[11][38] = 16'b0000000000000110;
    assign weights1[11][39] = 16'b1111111111111111;
    assign weights1[11][40] = 16'b1111111111110110;
    assign weights1[11][41] = 16'b1111111111111011;
    assign weights1[11][42] = 16'b0000000000000010;
    assign weights1[11][43] = 16'b1111111111110111;
    assign weights1[11][44] = 16'b1111111111111010;
    assign weights1[11][45] = 16'b1111111111110111;
    assign weights1[11][46] = 16'b0000000000001100;
    assign weights1[11][47] = 16'b1111111111111110;
    assign weights1[11][48] = 16'b1111111111111001;
    assign weights1[11][49] = 16'b0000000000000011;
    assign weights1[11][50] = 16'b1111111111111000;
    assign weights1[11][51] = 16'b1111111111111011;
    assign weights1[11][52] = 16'b1111111111101100;
    assign weights1[11][53] = 16'b1111111111110111;
    assign weights1[11][54] = 16'b1111111111110111;
    assign weights1[11][55] = 16'b1111111111111110;
    assign weights1[11][56] = 16'b0000000000000001;
    assign weights1[11][57] = 16'b0000000000000100;
    assign weights1[11][58] = 16'b0000000000000111;
    assign weights1[11][59] = 16'b0000000000000110;
    assign weights1[11][60] = 16'b0000000000000111;
    assign weights1[11][61] = 16'b0000000000000010;
    assign weights1[11][62] = 16'b0000000000001000;
    assign weights1[11][63] = 16'b1111111111110000;
    assign weights1[11][64] = 16'b1111111111111101;
    assign weights1[11][65] = 16'b1111111111110111;
    assign weights1[11][66] = 16'b1111111111111101;
    assign weights1[11][67] = 16'b0000000000000001;
    assign weights1[11][68] = 16'b0000000000000000;
    assign weights1[11][69] = 16'b0000000000000110;
    assign weights1[11][70] = 16'b0000000000010010;
    assign weights1[11][71] = 16'b1111111111111000;
    assign weights1[11][72] = 16'b1111111111111010;
    assign weights1[11][73] = 16'b1111111111101110;
    assign weights1[11][74] = 16'b1111111111101110;
    assign weights1[11][75] = 16'b1111111111101100;
    assign weights1[11][76] = 16'b1111111111111111;
    assign weights1[11][77] = 16'b1111111111111001;
    assign weights1[11][78] = 16'b1111111111110110;
    assign weights1[11][79] = 16'b1111111111111101;
    assign weights1[11][80] = 16'b1111111111111011;
    assign weights1[11][81] = 16'b0000000000000000;
    assign weights1[11][82] = 16'b0000000000001000;
    assign weights1[11][83] = 16'b1111111111111111;
    assign weights1[11][84] = 16'b0000000000000100;
    assign weights1[11][85] = 16'b0000000000000111;
    assign weights1[11][86] = 16'b0000000000000001;
    assign weights1[11][87] = 16'b1111111111111001;
    assign weights1[11][88] = 16'b0000000000000001;
    assign weights1[11][89] = 16'b0000000000000000;
    assign weights1[11][90] = 16'b0000000000001000;
    assign weights1[11][91] = 16'b1111111111111100;
    assign weights1[11][92] = 16'b0000000000001000;
    assign weights1[11][93] = 16'b0000000000010000;
    assign weights1[11][94] = 16'b0000000000001101;
    assign weights1[11][95] = 16'b0000000000010000;
    assign weights1[11][96] = 16'b1111111111111100;
    assign weights1[11][97] = 16'b1111111111100010;
    assign weights1[11][98] = 16'b1111111111101100;
    assign weights1[11][99] = 16'b1111111111101011;
    assign weights1[11][100] = 16'b0000000000000011;
    assign weights1[11][101] = 16'b0000000000100000;
    assign weights1[11][102] = 16'b1111111111111100;
    assign weights1[11][103] = 16'b1111111111111111;
    assign weights1[11][104] = 16'b1111111111111010;
    assign weights1[11][105] = 16'b0000000000000000;
    assign weights1[11][106] = 16'b0000000000000001;
    assign weights1[11][107] = 16'b1111111111110100;
    assign weights1[11][108] = 16'b1111111111111110;
    assign weights1[11][109] = 16'b1111111111110111;
    assign weights1[11][110] = 16'b0000000000000000;
    assign weights1[11][111] = 16'b1111111111111100;
    assign weights1[11][112] = 16'b0000000000000110;
    assign weights1[11][113] = 16'b0000000000001010;
    assign weights1[11][114] = 16'b1111111111111100;
    assign weights1[11][115] = 16'b1111111111110100;
    assign weights1[11][116] = 16'b0000000000000010;
    assign weights1[11][117] = 16'b0000000000011000;
    assign weights1[11][118] = 16'b0000000000010010;
    assign weights1[11][119] = 16'b0000000000001011;
    assign weights1[11][120] = 16'b0000000000001000;
    assign weights1[11][121] = 16'b1111111111110101;
    assign weights1[11][122] = 16'b1111111111110111;
    assign weights1[11][123] = 16'b0000000000000001;
    assign weights1[11][124] = 16'b0000000000000011;
    assign weights1[11][125] = 16'b1111111111111011;
    assign weights1[11][126] = 16'b0000000000010001;
    assign weights1[11][127] = 16'b0000000000011010;
    assign weights1[11][128] = 16'b1111111111111101;
    assign weights1[11][129] = 16'b1111111111111001;
    assign weights1[11][130] = 16'b0000000000010111;
    assign weights1[11][131] = 16'b1111111111110011;
    assign weights1[11][132] = 16'b0000000000011101;
    assign weights1[11][133] = 16'b1111111111110000;
    assign weights1[11][134] = 16'b0000000000001111;
    assign weights1[11][135] = 16'b0000000000001010;
    assign weights1[11][136] = 16'b1111111111101011;
    assign weights1[11][137] = 16'b1111111111111001;
    assign weights1[11][138] = 16'b1111111111111111;
    assign weights1[11][139] = 16'b1111111111111011;
    assign weights1[11][140] = 16'b0000000000000011;
    assign weights1[11][141] = 16'b0000000000000110;
    assign weights1[11][142] = 16'b1111111111111101;
    assign weights1[11][143] = 16'b1111111111111011;
    assign weights1[11][144] = 16'b0000000000010010;
    assign weights1[11][145] = 16'b1111111111111011;
    assign weights1[11][146] = 16'b0000000000001111;
    assign weights1[11][147] = 16'b0000000000001100;
    assign weights1[11][148] = 16'b1111111111111110;
    assign weights1[11][149] = 16'b1111111111110111;
    assign weights1[11][150] = 16'b0000000000001100;
    assign weights1[11][151] = 16'b0000000000001110;
    assign weights1[11][152] = 16'b0000000000000110;
    assign weights1[11][153] = 16'b1111111111111110;
    assign weights1[11][154] = 16'b1111111111110001;
    assign weights1[11][155] = 16'b1111111111111010;
    assign weights1[11][156] = 16'b0000000000000000;
    assign weights1[11][157] = 16'b0000000000000000;
    assign weights1[11][158] = 16'b1111111111111101;
    assign weights1[11][159] = 16'b0000000000010100;
    assign weights1[11][160] = 16'b0000000000001110;
    assign weights1[11][161] = 16'b0000000000000010;
    assign weights1[11][162] = 16'b1111111111111001;
    assign weights1[11][163] = 16'b0000000000001001;
    assign weights1[11][164] = 16'b1111111111111110;
    assign weights1[11][165] = 16'b1111111111111110;
    assign weights1[11][166] = 16'b1111111111111010;
    assign weights1[11][167] = 16'b1111111111110110;
    assign weights1[11][168] = 16'b0000000000000001;
    assign weights1[11][169] = 16'b0000000000000101;
    assign weights1[11][170] = 16'b0000000000001001;
    assign weights1[11][171] = 16'b0000000000000110;
    assign weights1[11][172] = 16'b0000000000010010;
    assign weights1[11][173] = 16'b0000000000000000;
    assign weights1[11][174] = 16'b0000000000010101;
    assign weights1[11][175] = 16'b0000000000000001;
    assign weights1[11][176] = 16'b1111111111110001;
    assign weights1[11][177] = 16'b0000000000010011;
    assign weights1[11][178] = 16'b0000000000011101;
    assign weights1[11][179] = 16'b0000000000000111;
    assign weights1[11][180] = 16'b0000000000001010;
    assign weights1[11][181] = 16'b1111111111111011;
    assign weights1[11][182] = 16'b0000000000010111;
    assign weights1[11][183] = 16'b1111111111111101;
    assign weights1[11][184] = 16'b0000000000000110;
    assign weights1[11][185] = 16'b1111111111111010;
    assign weights1[11][186] = 16'b0000000000000001;
    assign weights1[11][187] = 16'b0000000000000000;
    assign weights1[11][188] = 16'b1111111111110010;
    assign weights1[11][189] = 16'b1111111111110110;
    assign weights1[11][190] = 16'b1111111111111001;
    assign weights1[11][191] = 16'b1111111111110110;
    assign weights1[11][192] = 16'b0000000000000100;
    assign weights1[11][193] = 16'b1111111111110111;
    assign weights1[11][194] = 16'b1111111111111111;
    assign weights1[11][195] = 16'b1111111111101110;
    assign weights1[11][196] = 16'b0000000000000110;
    assign weights1[11][197] = 16'b0000000000000000;
    assign weights1[11][198] = 16'b0000000000010010;
    assign weights1[11][199] = 16'b0000000000001100;
    assign weights1[11][200] = 16'b1111111111110110;
    assign weights1[11][201] = 16'b1111111111111101;
    assign weights1[11][202] = 16'b0000000000011001;
    assign weights1[11][203] = 16'b0000000000001101;
    assign weights1[11][204] = 16'b0000000000011110;
    assign weights1[11][205] = 16'b0000000000011111;
    assign weights1[11][206] = 16'b0000000000010100;
    assign weights1[11][207] = 16'b1111111111111100;
    assign weights1[11][208] = 16'b0000000000000111;
    assign weights1[11][209] = 16'b0000000000010111;
    assign weights1[11][210] = 16'b0000000000000101;
    assign weights1[11][211] = 16'b0000000000001111;
    assign weights1[11][212] = 16'b0000000000001111;
    assign weights1[11][213] = 16'b0000000000001110;
    assign weights1[11][214] = 16'b0000000000000000;
    assign weights1[11][215] = 16'b0000000000000100;
    assign weights1[11][216] = 16'b0000000000010011;
    assign weights1[11][217] = 16'b1111111111111101;
    assign weights1[11][218] = 16'b0000000000001010;
    assign weights1[11][219] = 16'b1111111111111011;
    assign weights1[11][220] = 16'b1111111111111100;
    assign weights1[11][221] = 16'b1111111111110111;
    assign weights1[11][222] = 16'b1111111111111010;
    assign weights1[11][223] = 16'b1111111111110011;
    assign weights1[11][224] = 16'b0000000000001100;
    assign weights1[11][225] = 16'b0000000000001001;
    assign weights1[11][226] = 16'b0000000000010101;
    assign weights1[11][227] = 16'b0000000000001111;
    assign weights1[11][228] = 16'b0000000000100100;
    assign weights1[11][229] = 16'b0000000000000011;
    assign weights1[11][230] = 16'b0000000000000111;
    assign weights1[11][231] = 16'b0000000000011100;
    assign weights1[11][232] = 16'b0000000000101010;
    assign weights1[11][233] = 16'b0000000000001110;
    assign weights1[11][234] = 16'b1111111111110110;
    assign weights1[11][235] = 16'b0000000000101110;
    assign weights1[11][236] = 16'b0000000000001010;
    assign weights1[11][237] = 16'b0000000000000000;
    assign weights1[11][238] = 16'b0000000000100100;
    assign weights1[11][239] = 16'b0000000000001101;
    assign weights1[11][240] = 16'b0000000000010001;
    assign weights1[11][241] = 16'b1111111111111110;
    assign weights1[11][242] = 16'b1111111111110010;
    assign weights1[11][243] = 16'b0000000000000100;
    assign weights1[11][244] = 16'b0000000000000101;
    assign weights1[11][245] = 16'b1111111111110111;
    assign weights1[11][246] = 16'b0000000000000101;
    assign weights1[11][247] = 16'b0000000000000111;
    assign weights1[11][248] = 16'b0000000000000100;
    assign weights1[11][249] = 16'b0000000000000111;
    assign weights1[11][250] = 16'b0000000000000100;
    assign weights1[11][251] = 16'b1111111111110001;
    assign weights1[11][252] = 16'b0000000000001011;
    assign weights1[11][253] = 16'b0000000000001100;
    assign weights1[11][254] = 16'b0000000000011001;
    assign weights1[11][255] = 16'b0000000000100100;
    assign weights1[11][256] = 16'b0000000000110000;
    assign weights1[11][257] = 16'b0000000000101011;
    assign weights1[11][258] = 16'b0000000000100011;
    assign weights1[11][259] = 16'b0000000000010111;
    assign weights1[11][260] = 16'b0000000000101000;
    assign weights1[11][261] = 16'b0000000000101101;
    assign weights1[11][262] = 16'b0000000000101011;
    assign weights1[11][263] = 16'b0000000000110111;
    assign weights1[11][264] = 16'b0000000000101110;
    assign weights1[11][265] = 16'b0000000000101011;
    assign weights1[11][266] = 16'b0000000000010100;
    assign weights1[11][267] = 16'b0000000000000111;
    assign weights1[11][268] = 16'b0000000000001101;
    assign weights1[11][269] = 16'b0000000000001100;
    assign weights1[11][270] = 16'b0000000000001110;
    assign weights1[11][271] = 16'b0000000000000111;
    assign weights1[11][272] = 16'b0000000000001100;
    assign weights1[11][273] = 16'b0000000000000111;
    assign weights1[11][274] = 16'b1111111111111100;
    assign weights1[11][275] = 16'b1111111111110000;
    assign weights1[11][276] = 16'b0000000000001001;
    assign weights1[11][277] = 16'b1111111111101101;
    assign weights1[11][278] = 16'b1111111111111110;
    assign weights1[11][279] = 16'b1111111111100111;
    assign weights1[11][280] = 16'b0000000000001100;
    assign weights1[11][281] = 16'b0000000000010111;
    assign weights1[11][282] = 16'b0000000000100110;
    assign weights1[11][283] = 16'b0000000000101011;
    assign weights1[11][284] = 16'b0000000000110001;
    assign weights1[11][285] = 16'b0000000001001111;
    assign weights1[11][286] = 16'b0000000000100100;
    assign weights1[11][287] = 16'b0000000000111110;
    assign weights1[11][288] = 16'b0000000001001101;
    assign weights1[11][289] = 16'b0000000001010100;
    assign weights1[11][290] = 16'b0000000000110110;
    assign weights1[11][291] = 16'b0000000000101110;
    assign weights1[11][292] = 16'b0000000000011110;
    assign weights1[11][293] = 16'b0000000000010011;
    assign weights1[11][294] = 16'b0000000000000010;
    assign weights1[11][295] = 16'b0000000000001000;
    assign weights1[11][296] = 16'b0000000000001110;
    assign weights1[11][297] = 16'b1111111111111111;
    assign weights1[11][298] = 16'b0000000000000010;
    assign weights1[11][299] = 16'b0000000000000001;
    assign weights1[11][300] = 16'b1111111111111010;
    assign weights1[11][301] = 16'b1111111111110001;
    assign weights1[11][302] = 16'b1111111111111010;
    assign weights1[11][303] = 16'b1111111111100110;
    assign weights1[11][304] = 16'b0000000000000000;
    assign weights1[11][305] = 16'b1111111111110010;
    assign weights1[11][306] = 16'b1111111111111011;
    assign weights1[11][307] = 16'b1111111111110100;
    assign weights1[11][308] = 16'b1111111111111101;
    assign weights1[11][309] = 16'b1111111111111101;
    assign weights1[11][310] = 16'b0000000000010100;
    assign weights1[11][311] = 16'b0000000000010001;
    assign weights1[11][312] = 16'b0000000000010000;
    assign weights1[11][313] = 16'b0000000000100110;
    assign weights1[11][314] = 16'b0000000000100100;
    assign weights1[11][315] = 16'b0000000000110001;
    assign weights1[11][316] = 16'b0000000000010000;
    assign weights1[11][317] = 16'b0000000000000010;
    assign weights1[11][318] = 16'b1111111111011011;
    assign weights1[11][319] = 16'b1111111111100111;
    assign weights1[11][320] = 16'b1111111111011111;
    assign weights1[11][321] = 16'b1111111111010110;
    assign weights1[11][322] = 16'b1111111111100010;
    assign weights1[11][323] = 16'b1111111111100010;
    assign weights1[11][324] = 16'b1111111111101000;
    assign weights1[11][325] = 16'b1111111111110101;
    assign weights1[11][326] = 16'b1111111111101101;
    assign weights1[11][327] = 16'b0000000000000101;
    assign weights1[11][328] = 16'b1111111111111001;
    assign weights1[11][329] = 16'b1111111111111001;
    assign weights1[11][330] = 16'b1111111111110010;
    assign weights1[11][331] = 16'b0000000000000001;
    assign weights1[11][332] = 16'b1111111111110001;
    assign weights1[11][333] = 16'b1111111111110011;
    assign weights1[11][334] = 16'b1111111111111000;
    assign weights1[11][335] = 16'b1111111111111111;
    assign weights1[11][336] = 16'b1111111111101101;
    assign weights1[11][337] = 16'b1111111111101000;
    assign weights1[11][338] = 16'b1111111111100101;
    assign weights1[11][339] = 16'b1111111111110100;
    assign weights1[11][340] = 16'b1111111111101011;
    assign weights1[11][341] = 16'b1111111111100101;
    assign weights1[11][342] = 16'b1111111111011010;
    assign weights1[11][343] = 16'b1111111110101111;
    assign weights1[11][344] = 16'b1111111110011001;
    assign weights1[11][345] = 16'b1111111101011001;
    assign weights1[11][346] = 16'b1111111101101001;
    assign weights1[11][347] = 16'b1111111101000110;
    assign weights1[11][348] = 16'b1111111101100011;
    assign weights1[11][349] = 16'b1111111110011101;
    assign weights1[11][350] = 16'b1111111110100011;
    assign weights1[11][351] = 16'b1111111111010010;
    assign weights1[11][352] = 16'b1111111111100010;
    assign weights1[11][353] = 16'b1111111111011100;
    assign weights1[11][354] = 16'b1111111111100001;
    assign weights1[11][355] = 16'b1111111111101111;
    assign weights1[11][356] = 16'b1111111111110110;
    assign weights1[11][357] = 16'b1111111111111110;
    assign weights1[11][358] = 16'b1111111111110000;
    assign weights1[11][359] = 16'b1111111111101111;
    assign weights1[11][360] = 16'b1111111111111000;
    assign weights1[11][361] = 16'b1111111111111101;
    assign weights1[11][362] = 16'b1111111111111010;
    assign weights1[11][363] = 16'b0000000000001011;
    assign weights1[11][364] = 16'b1111111111010100;
    assign weights1[11][365] = 16'b1111111110111000;
    assign weights1[11][366] = 16'b1111111110111000;
    assign weights1[11][367] = 16'b1111111110011101;
    assign weights1[11][368] = 16'b1111111110010000;
    assign weights1[11][369] = 16'b1111111110000010;
    assign weights1[11][370] = 16'b1111111101100011;
    assign weights1[11][371] = 16'b1111111011110011;
    assign weights1[11][372] = 16'b1111111010111001;
    assign weights1[11][373] = 16'b1111111011011110;
    assign weights1[11][374] = 16'b1111111100110100;
    assign weights1[11][375] = 16'b1111111110011011;
    assign weights1[11][376] = 16'b1111111111001100;
    assign weights1[11][377] = 16'b1111111111100010;
    assign weights1[11][378] = 16'b1111111111100010;
    assign weights1[11][379] = 16'b1111111111011001;
    assign weights1[11][380] = 16'b1111111111101111;
    assign weights1[11][381] = 16'b1111111111110100;
    assign weights1[11][382] = 16'b1111111111110101;
    assign weights1[11][383] = 16'b1111111111101000;
    assign weights1[11][384] = 16'b1111111111110001;
    assign weights1[11][385] = 16'b0000000000000100;
    assign weights1[11][386] = 16'b1111111111111011;
    assign weights1[11][387] = 16'b0000000000000111;
    assign weights1[11][388] = 16'b0000000000001111;
    assign weights1[11][389] = 16'b1111111111111001;
    assign weights1[11][390] = 16'b0000000000001011;
    assign weights1[11][391] = 16'b0000000000001011;
    assign weights1[11][392] = 16'b1111111110111100;
    assign weights1[11][393] = 16'b1111111110010110;
    assign weights1[11][394] = 16'b1111111110010000;
    assign weights1[11][395] = 16'b1111111101101100;
    assign weights1[11][396] = 16'b1111111101001011;
    assign weights1[11][397] = 16'b1111111100011111;
    assign weights1[11][398] = 16'b1111111100010010;
    assign weights1[11][399] = 16'b1111111100001000;
    assign weights1[11][400] = 16'b1111111101110111;
    assign weights1[11][401] = 16'b1111111111110010;
    assign weights1[11][402] = 16'b0000000000001111;
    assign weights1[11][403] = 16'b0000000000001011;
    assign weights1[11][404] = 16'b0000000000010001;
    assign weights1[11][405] = 16'b1111111111111001;
    assign weights1[11][406] = 16'b1111111111111111;
    assign weights1[11][407] = 16'b0000000000000010;
    assign weights1[11][408] = 16'b0000000000000110;
    assign weights1[11][409] = 16'b0000000000000000;
    assign weights1[11][410] = 16'b0000000000001001;
    assign weights1[11][411] = 16'b0000000000001011;
    assign weights1[11][412] = 16'b0000000000000100;
    assign weights1[11][413] = 16'b0000000000010011;
    assign weights1[11][414] = 16'b0000000000001111;
    assign weights1[11][415] = 16'b0000000000001011;
    assign weights1[11][416] = 16'b0000000000010010;
    assign weights1[11][417] = 16'b0000000000000101;
    assign weights1[11][418] = 16'b0000000000010110;
    assign weights1[11][419] = 16'b0000000000001101;
    assign weights1[11][420] = 16'b1111111110111011;
    assign weights1[11][421] = 16'b1111111110010010;
    assign weights1[11][422] = 16'b1111111110010001;
    assign weights1[11][423] = 16'b1111111101100001;
    assign weights1[11][424] = 16'b1111111101000111;
    assign weights1[11][425] = 16'b1111111101100011;
    assign weights1[11][426] = 16'b1111111110001011;
    assign weights1[11][427] = 16'b1111111111101110;
    assign weights1[11][428] = 16'b0000000000110000;
    assign weights1[11][429] = 16'b0000000000110100;
    assign weights1[11][430] = 16'b0000000001000011;
    assign weights1[11][431] = 16'b0000000000101011;
    assign weights1[11][432] = 16'b0000000000010110;
    assign weights1[11][433] = 16'b0000000000011110;
    assign weights1[11][434] = 16'b0000000000001101;
    assign weights1[11][435] = 16'b0000000000001001;
    assign weights1[11][436] = 16'b0000000000000010;
    assign weights1[11][437] = 16'b0000000000000011;
    assign weights1[11][438] = 16'b0000000000000000;
    assign weights1[11][439] = 16'b0000000000001101;
    assign weights1[11][440] = 16'b0000000000000110;
    assign weights1[11][441] = 16'b0000000000000000;
    assign weights1[11][442] = 16'b1111111111111011;
    assign weights1[11][443] = 16'b0000000000001110;
    assign weights1[11][444] = 16'b1111111111111111;
    assign weights1[11][445] = 16'b0000000000000101;
    assign weights1[11][446] = 16'b1111111111111110;
    assign weights1[11][447] = 16'b1111111111111110;
    assign weights1[11][448] = 16'b1111111111000011;
    assign weights1[11][449] = 16'b1111111110101100;
    assign weights1[11][450] = 16'b1111111110101111;
    assign weights1[11][451] = 16'b1111111110011101;
    assign weights1[11][452] = 16'b1111111110101011;
    assign weights1[11][453] = 16'b1111111111100000;
    assign weights1[11][454] = 16'b0000000000010101;
    assign weights1[11][455] = 16'b0000000001000100;
    assign weights1[11][456] = 16'b0000000000110111;
    assign weights1[11][457] = 16'b0000000000011010;
    assign weights1[11][458] = 16'b0000000000010110;
    assign weights1[11][459] = 16'b0000000000000101;
    assign weights1[11][460] = 16'b0000000000000011;
    assign weights1[11][461] = 16'b0000000000001001;
    assign weights1[11][462] = 16'b0000000000010000;
    assign weights1[11][463] = 16'b1111111111111101;
    assign weights1[11][464] = 16'b0000000000000011;
    assign weights1[11][465] = 16'b0000000000000110;
    assign weights1[11][466] = 16'b0000000000010001;
    assign weights1[11][467] = 16'b1111111111111010;
    assign weights1[11][468] = 16'b1111111111111101;
    assign weights1[11][469] = 16'b0000000000001100;
    assign weights1[11][470] = 16'b0000000000000110;
    assign weights1[11][471] = 16'b0000000000010101;
    assign weights1[11][472] = 16'b0000000000000000;
    assign weights1[11][473] = 16'b0000000000001010;
    assign weights1[11][474] = 16'b1111111111111111;
    assign weights1[11][475] = 16'b1111111111111111;
    assign weights1[11][476] = 16'b1111111111010000;
    assign weights1[11][477] = 16'b1111111111000110;
    assign weights1[11][478] = 16'b1111111111001100;
    assign weights1[11][479] = 16'b1111111111101010;
    assign weights1[11][480] = 16'b0000000000010010;
    assign weights1[11][481] = 16'b0000000000111010;
    assign weights1[11][482] = 16'b0000000001000110;
    assign weights1[11][483] = 16'b0000000000001000;
    assign weights1[11][484] = 16'b0000000000011010;
    assign weights1[11][485] = 16'b0000000000001111;
    assign weights1[11][486] = 16'b1111111111111001;
    assign weights1[11][487] = 16'b1111111111111011;
    assign weights1[11][488] = 16'b0000000000001001;
    assign weights1[11][489] = 16'b0000000000000010;
    assign weights1[11][490] = 16'b0000000000000010;
    assign weights1[11][491] = 16'b0000000000001010;
    assign weights1[11][492] = 16'b0000000000000111;
    assign weights1[11][493] = 16'b0000000000000110;
    assign weights1[11][494] = 16'b1111111111110111;
    assign weights1[11][495] = 16'b0000000000000111;
    assign weights1[11][496] = 16'b0000000000001111;
    assign weights1[11][497] = 16'b0000000000010011;
    assign weights1[11][498] = 16'b1111111111111010;
    assign weights1[11][499] = 16'b0000000000000101;
    assign weights1[11][500] = 16'b1111111111110000;
    assign weights1[11][501] = 16'b1111111111101111;
    assign weights1[11][502] = 16'b1111111111111010;
    assign weights1[11][503] = 16'b1111111111111101;
    assign weights1[11][504] = 16'b1111111111100011;
    assign weights1[11][505] = 16'b1111111111100000;
    assign weights1[11][506] = 16'b1111111111110011;
    assign weights1[11][507] = 16'b0000000000010001;
    assign weights1[11][508] = 16'b0000000000101001;
    assign weights1[11][509] = 16'b0000000000111010;
    assign weights1[11][510] = 16'b0000000000001101;
    assign weights1[11][511] = 16'b1111111111110101;
    assign weights1[11][512] = 16'b1111111111101100;
    assign weights1[11][513] = 16'b1111111111110001;
    assign weights1[11][514] = 16'b0000000000010011;
    assign weights1[11][515] = 16'b1111111111111001;
    assign weights1[11][516] = 16'b0000000000010000;
    assign weights1[11][517] = 16'b1111111111111110;
    assign weights1[11][518] = 16'b0000000000000001;
    assign weights1[11][519] = 16'b1111111111111001;
    assign weights1[11][520] = 16'b1111111111110001;
    assign weights1[11][521] = 16'b0000000000000110;
    assign weights1[11][522] = 16'b0000000000000100;
    assign weights1[11][523] = 16'b0000000000000101;
    assign weights1[11][524] = 16'b1111111111110100;
    assign weights1[11][525] = 16'b1111111111110001;
    assign weights1[11][526] = 16'b1111111111110000;
    assign weights1[11][527] = 16'b1111111111101001;
    assign weights1[11][528] = 16'b0000000000010011;
    assign weights1[11][529] = 16'b1111111111111110;
    assign weights1[11][530] = 16'b1111111111110110;
    assign weights1[11][531] = 16'b0000000000000011;
    assign weights1[11][532] = 16'b1111111111111100;
    assign weights1[11][533] = 16'b0000000000000100;
    assign weights1[11][534] = 16'b0000000000001011;
    assign weights1[11][535] = 16'b0000000000010110;
    assign weights1[11][536] = 16'b0000000000001100;
    assign weights1[11][537] = 16'b1111111111110110;
    assign weights1[11][538] = 16'b1111111111110000;
    assign weights1[11][539] = 16'b0000000000011001;
    assign weights1[11][540] = 16'b0000000000001100;
    assign weights1[11][541] = 16'b0000000000010001;
    assign weights1[11][542] = 16'b1111111111111111;
    assign weights1[11][543] = 16'b0000000000001010;
    assign weights1[11][544] = 16'b0000000000000011;
    assign weights1[11][545] = 16'b1111111111111111;
    assign weights1[11][546] = 16'b0000000000000001;
    assign weights1[11][547] = 16'b1111111111111010;
    assign weights1[11][548] = 16'b1111111111111111;
    assign weights1[11][549] = 16'b1111111111111100;
    assign weights1[11][550] = 16'b1111111111101000;
    assign weights1[11][551] = 16'b1111111111111011;
    assign weights1[11][552] = 16'b0000000000001000;
    assign weights1[11][553] = 16'b1111111111110010;
    assign weights1[11][554] = 16'b0000000000010111;
    assign weights1[11][555] = 16'b1111111111111011;
    assign weights1[11][556] = 16'b1111111111101011;
    assign weights1[11][557] = 16'b1111111111111011;
    assign weights1[11][558] = 16'b1111111111110011;
    assign weights1[11][559] = 16'b0000000000001001;
    assign weights1[11][560] = 16'b0000000000010101;
    assign weights1[11][561] = 16'b0000000000011101;
    assign weights1[11][562] = 16'b1111111111111111;
    assign weights1[11][563] = 16'b0000000000001010;
    assign weights1[11][564] = 16'b0000000000001100;
    assign weights1[11][565] = 16'b1111111111111010;
    assign weights1[11][566] = 16'b0000000000001110;
    assign weights1[11][567] = 16'b0000000000001100;
    assign weights1[11][568] = 16'b0000000000001010;
    assign weights1[11][569] = 16'b0000000000001110;
    assign weights1[11][570] = 16'b1111111111101010;
    assign weights1[11][571] = 16'b1111111111111110;
    assign weights1[11][572] = 16'b1111111111111110;
    assign weights1[11][573] = 16'b0000000000001001;
    assign weights1[11][574] = 16'b1111111111101101;
    assign weights1[11][575] = 16'b0000000000000100;
    assign weights1[11][576] = 16'b0000000000000000;
    assign weights1[11][577] = 16'b1111111111110101;
    assign weights1[11][578] = 16'b0000000000000100;
    assign weights1[11][579] = 16'b1111111111110001;
    assign weights1[11][580] = 16'b0000000000000001;
    assign weights1[11][581] = 16'b1111111111111000;
    assign weights1[11][582] = 16'b0000000000000100;
    assign weights1[11][583] = 16'b1111111111110001;
    assign weights1[11][584] = 16'b0000000000010000;
    assign weights1[11][585] = 16'b1111111111110001;
    assign weights1[11][586] = 16'b1111111111101101;
    assign weights1[11][587] = 16'b1111111111111100;
    assign weights1[11][588] = 16'b0000000000010010;
    assign weights1[11][589] = 16'b0000000000010001;
    assign weights1[11][590] = 16'b0000000000000001;
    assign weights1[11][591] = 16'b0000000000001100;
    assign weights1[11][592] = 16'b1111111111110111;
    assign weights1[11][593] = 16'b0000000000010010;
    assign weights1[11][594] = 16'b1111111111111100;
    assign weights1[11][595] = 16'b0000000000000100;
    assign weights1[11][596] = 16'b1111111111111000;
    assign weights1[11][597] = 16'b0000000000001001;
    assign weights1[11][598] = 16'b0000000000001001;
    assign weights1[11][599] = 16'b0000000000000000;
    assign weights1[11][600] = 16'b0000000000001010;
    assign weights1[11][601] = 16'b1111111111101001;
    assign weights1[11][602] = 16'b0000000000001011;
    assign weights1[11][603] = 16'b0000000000000100;
    assign weights1[11][604] = 16'b1111111111110110;
    assign weights1[11][605] = 16'b1111111111111100;
    assign weights1[11][606] = 16'b0000000000001000;
    assign weights1[11][607] = 16'b1111111111111001;
    assign weights1[11][608] = 16'b1111111111111100;
    assign weights1[11][609] = 16'b0000000000001101;
    assign weights1[11][610] = 16'b0000000000000111;
    assign weights1[11][611] = 16'b0000000000010001;
    assign weights1[11][612] = 16'b1111111111111101;
    assign weights1[11][613] = 16'b1111111111111100;
    assign weights1[11][614] = 16'b1111111111111001;
    assign weights1[11][615] = 16'b0000000000001000;
    assign weights1[11][616] = 16'b0000000000000101;
    assign weights1[11][617] = 16'b0000000000001110;
    assign weights1[11][618] = 16'b0000000000000110;
    assign weights1[11][619] = 16'b0000000000010011;
    assign weights1[11][620] = 16'b0000000000000111;
    assign weights1[11][621] = 16'b1111111111111100;
    assign weights1[11][622] = 16'b1111111111111010;
    assign weights1[11][623] = 16'b1111111111111100;
    assign weights1[11][624] = 16'b0000000000001010;
    assign weights1[11][625] = 16'b1111111111111100;
    assign weights1[11][626] = 16'b0000000000000111;
    assign weights1[11][627] = 16'b1111111111111110;
    assign weights1[11][628] = 16'b1111111111111111;
    assign weights1[11][629] = 16'b0000000000000100;
    assign weights1[11][630] = 16'b0000000000000001;
    assign weights1[11][631] = 16'b0000000000000001;
    assign weights1[11][632] = 16'b0000000000011100;
    assign weights1[11][633] = 16'b0000000000000001;
    assign weights1[11][634] = 16'b1111111111110110;
    assign weights1[11][635] = 16'b1111111111110111;
    assign weights1[11][636] = 16'b0000000000010101;
    assign weights1[11][637] = 16'b1111111111110110;
    assign weights1[11][638] = 16'b1111111111110110;
    assign weights1[11][639] = 16'b0000000000000001;
    assign weights1[11][640] = 16'b0000000000000100;
    assign weights1[11][641] = 16'b1111111111111100;
    assign weights1[11][642] = 16'b0000000000000000;
    assign weights1[11][643] = 16'b0000000000000110;
    assign weights1[11][644] = 16'b1111111111111110;
    assign weights1[11][645] = 16'b0000000000001011;
    assign weights1[11][646] = 16'b0000000000001000;
    assign weights1[11][647] = 16'b1111111111110111;
    assign weights1[11][648] = 16'b1111111111110110;
    assign weights1[11][649] = 16'b0000000000000110;
    assign weights1[11][650] = 16'b0000000000000011;
    assign weights1[11][651] = 16'b0000000000000000;
    assign weights1[11][652] = 16'b1111111111111101;
    assign weights1[11][653] = 16'b0000000000000110;
    assign weights1[11][654] = 16'b1111111111111101;
    assign weights1[11][655] = 16'b0000000000001101;
    assign weights1[11][656] = 16'b1111111111110110;
    assign weights1[11][657] = 16'b1111111111111101;
    assign weights1[11][658] = 16'b0000000000001010;
    assign weights1[11][659] = 16'b1111111111110001;
    assign weights1[11][660] = 16'b1111111111110111;
    assign weights1[11][661] = 16'b0000000000000110;
    assign weights1[11][662] = 16'b0000000000011101;
    assign weights1[11][663] = 16'b1111111111111100;
    assign weights1[11][664] = 16'b1111111111110001;
    assign weights1[11][665] = 16'b1111111111110010;
    assign weights1[11][666] = 16'b1111111111101011;
    assign weights1[11][667] = 16'b0000000000001000;
    assign weights1[11][668] = 16'b0000000000010101;
    assign weights1[11][669] = 16'b1111111111111101;
    assign weights1[11][670] = 16'b1111111111111110;
    assign weights1[11][671] = 16'b0000000000001010;
    assign weights1[11][672] = 16'b0000000000001011;
    assign weights1[11][673] = 16'b0000000000000010;
    assign weights1[11][674] = 16'b0000000000001010;
    assign weights1[11][675] = 16'b1111111111111111;
    assign weights1[11][676] = 16'b0000000000000100;
    assign weights1[11][677] = 16'b0000000000000100;
    assign weights1[11][678] = 16'b0000000000001110;
    assign weights1[11][679] = 16'b1111111111111000;
    assign weights1[11][680] = 16'b0000000000000010;
    assign weights1[11][681] = 16'b0000000000001010;
    assign weights1[11][682] = 16'b1111111111110010;
    assign weights1[11][683] = 16'b1111111111111001;
    assign weights1[11][684] = 16'b1111111111110010;
    assign weights1[11][685] = 16'b0000000000000010;
    assign weights1[11][686] = 16'b1111111111111100;
    assign weights1[11][687] = 16'b0000000000010001;
    assign weights1[11][688] = 16'b1111111111111110;
    assign weights1[11][689] = 16'b0000000000000100;
    assign weights1[11][690] = 16'b0000000000000011;
    assign weights1[11][691] = 16'b0000000000010000;
    assign weights1[11][692] = 16'b0000000000001000;
    assign weights1[11][693] = 16'b0000000000001000;
    assign weights1[11][694] = 16'b0000000000000000;
    assign weights1[11][695] = 16'b1111111111101110;
    assign weights1[11][696] = 16'b0000000000001101;
    assign weights1[11][697] = 16'b0000000000000100;
    assign weights1[11][698] = 16'b0000000000000110;
    assign weights1[11][699] = 16'b0000000000001000;
    assign weights1[11][700] = 16'b0000000000000110;
    assign weights1[11][701] = 16'b1111111111111111;
    assign weights1[11][702] = 16'b1111111111111110;
    assign weights1[11][703] = 16'b1111111111111011;
    assign weights1[11][704] = 16'b1111111111110111;
    assign weights1[11][705] = 16'b1111111111111010;
    assign weights1[11][706] = 16'b0000000000000100;
    assign weights1[11][707] = 16'b0000000000001000;
    assign weights1[11][708] = 16'b0000000000000111;
    assign weights1[11][709] = 16'b0000000000001100;
    assign weights1[11][710] = 16'b0000000000010011;
    assign weights1[11][711] = 16'b1111111111110111;
    assign weights1[11][712] = 16'b0000000000001100;
    assign weights1[11][713] = 16'b0000000000001010;
    assign weights1[11][714] = 16'b1111111111110111;
    assign weights1[11][715] = 16'b0000000000000000;
    assign weights1[11][716] = 16'b0000000000000101;
    assign weights1[11][717] = 16'b1111111111110110;
    assign weights1[11][718] = 16'b1111111111111101;
    assign weights1[11][719] = 16'b0000000000001010;
    assign weights1[11][720] = 16'b1111111111111100;
    assign weights1[11][721] = 16'b0000000000001001;
    assign weights1[11][722] = 16'b0000000000000110;
    assign weights1[11][723] = 16'b0000000000000110;
    assign weights1[11][724] = 16'b1111111111111010;
    assign weights1[11][725] = 16'b0000000000001011;
    assign weights1[11][726] = 16'b0000000000001010;
    assign weights1[11][727] = 16'b0000000000000110;
    assign weights1[11][728] = 16'b0000000000000001;
    assign weights1[11][729] = 16'b0000000000000010;
    assign weights1[11][730] = 16'b0000000000000000;
    assign weights1[11][731] = 16'b0000000000000011;
    assign weights1[11][732] = 16'b0000000000001011;
    assign weights1[11][733] = 16'b1111111111110011;
    assign weights1[11][734] = 16'b0000000000000100;
    assign weights1[11][735] = 16'b0000000000000001;
    assign weights1[11][736] = 16'b1111111111101111;
    assign weights1[11][737] = 16'b1111111111111011;
    assign weights1[11][738] = 16'b0000000000000010;
    assign weights1[11][739] = 16'b1111111111111100;
    assign weights1[11][740] = 16'b1111111111111101;
    assign weights1[11][741] = 16'b1111111111111111;
    assign weights1[11][742] = 16'b1111111111111111;
    assign weights1[11][743] = 16'b0000000000000010;
    assign weights1[11][744] = 16'b1111111111111110;
    assign weights1[11][745] = 16'b0000000000001001;
    assign weights1[11][746] = 16'b1111111111111001;
    assign weights1[11][747] = 16'b0000000000000011;
    assign weights1[11][748] = 16'b0000000000000100;
    assign weights1[11][749] = 16'b0000000000001100;
    assign weights1[11][750] = 16'b0000000000000011;
    assign weights1[11][751] = 16'b0000000000001000;
    assign weights1[11][752] = 16'b0000000000001000;
    assign weights1[11][753] = 16'b0000000000010001;
    assign weights1[11][754] = 16'b0000000000001001;
    assign weights1[11][755] = 16'b0000000000000011;
    assign weights1[11][756] = 16'b0000000000000110;
    assign weights1[11][757] = 16'b0000000000001000;
    assign weights1[11][758] = 16'b0000000000001101;
    assign weights1[11][759] = 16'b0000000000001100;
    assign weights1[11][760] = 16'b0000000000001010;
    assign weights1[11][761] = 16'b1111111111111110;
    assign weights1[11][762] = 16'b0000000000000100;
    assign weights1[11][763] = 16'b0000000000001100;
    assign weights1[11][764] = 16'b0000000000000101;
    assign weights1[11][765] = 16'b0000000000001001;
    assign weights1[11][766] = 16'b0000000000000010;
    assign weights1[11][767] = 16'b1111111111111011;
    assign weights1[11][768] = 16'b0000000000001010;
    assign weights1[11][769] = 16'b1111111111111100;
    assign weights1[11][770] = 16'b0000000000000001;
    assign weights1[11][771] = 16'b0000000000000011;
    assign weights1[11][772] = 16'b1111111111111100;
    assign weights1[11][773] = 16'b0000000000000010;
    assign weights1[11][774] = 16'b0000000000000101;
    assign weights1[11][775] = 16'b0000000000001001;
    assign weights1[11][776] = 16'b0000000000001110;
    assign weights1[11][777] = 16'b0000000000000101;
    assign weights1[11][778] = 16'b0000000000000111;
    assign weights1[11][779] = 16'b0000000000001101;
    assign weights1[11][780] = 16'b0000000000000111;
    assign weights1[11][781] = 16'b0000000000001000;
    assign weights1[11][782] = 16'b0000000000000110;
    assign weights1[11][783] = 16'b0000000000000100;
    assign weights1[12][0] = 16'b0000000000000000;
    assign weights1[12][1] = 16'b0000000000000010;
    assign weights1[12][2] = 16'b0000000000000011;
    assign weights1[12][3] = 16'b0000000000001000;
    assign weights1[12][4] = 16'b0000000000000011;
    assign weights1[12][5] = 16'b0000000000001100;
    assign weights1[12][6] = 16'b0000000000001111;
    assign weights1[12][7] = 16'b0000000000001001;
    assign weights1[12][8] = 16'b0000000000010101;
    assign weights1[12][9] = 16'b0000000000100001;
    assign weights1[12][10] = 16'b0000000000011111;
    assign weights1[12][11] = 16'b0000000000001110;
    assign weights1[12][12] = 16'b0000000000100001;
    assign weights1[12][13] = 16'b0000000000010111;
    assign weights1[12][14] = 16'b0000000000001101;
    assign weights1[12][15] = 16'b0000000000010100;
    assign weights1[12][16] = 16'b0000000000010101;
    assign weights1[12][17] = 16'b0000000000010000;
    assign weights1[12][18] = 16'b0000000000001011;
    assign weights1[12][19] = 16'b0000000000010001;
    assign weights1[12][20] = 16'b0000000000010011;
    assign weights1[12][21] = 16'b0000000000010000;
    assign weights1[12][22] = 16'b0000000000001000;
    assign weights1[12][23] = 16'b0000000000010100;
    assign weights1[12][24] = 16'b0000000000001001;
    assign weights1[12][25] = 16'b0000000000001011;
    assign weights1[12][26] = 16'b0000000000000110;
    assign weights1[12][27] = 16'b0000000000000101;
    assign weights1[12][28] = 16'b0000000000000001;
    assign weights1[12][29] = 16'b0000000000000101;
    assign weights1[12][30] = 16'b0000000000000111;
    assign weights1[12][31] = 16'b0000000000000110;
    assign weights1[12][32] = 16'b0000000000001000;
    assign weights1[12][33] = 16'b0000000000001110;
    assign weights1[12][34] = 16'b0000000000011101;
    assign weights1[12][35] = 16'b0000000000010001;
    assign weights1[12][36] = 16'b0000000000011000;
    assign weights1[12][37] = 16'b0000000000010110;
    assign weights1[12][38] = 16'b0000000000000111;
    assign weights1[12][39] = 16'b1111111111110010;
    assign weights1[12][40] = 16'b0000000000000111;
    assign weights1[12][41] = 16'b1111111111111110;
    assign weights1[12][42] = 16'b0000000000000011;
    assign weights1[12][43] = 16'b0000000000001010;
    assign weights1[12][44] = 16'b0000000000010001;
    assign weights1[12][45] = 16'b0000000000010011;
    assign weights1[12][46] = 16'b0000000000010110;
    assign weights1[12][47] = 16'b0000000000010010;
    assign weights1[12][48] = 16'b0000000000011010;
    assign weights1[12][49] = 16'b0000000000000100;
    assign weights1[12][50] = 16'b0000000000000101;
    assign weights1[12][51] = 16'b0000000000011011;
    assign weights1[12][52] = 16'b0000000000001011;
    assign weights1[12][53] = 16'b0000000000000111;
    assign weights1[12][54] = 16'b0000000000001011;
    assign weights1[12][55] = 16'b1111111111111010;
    assign weights1[12][56] = 16'b0000000000000111;
    assign weights1[12][57] = 16'b0000000000000111;
    assign weights1[12][58] = 16'b0000000000001010;
    assign weights1[12][59] = 16'b0000000000001001;
    assign weights1[12][60] = 16'b0000000000011011;
    assign weights1[12][61] = 16'b0000000000011111;
    assign weights1[12][62] = 16'b0000000000011111;
    assign weights1[12][63] = 16'b0000000000001011;
    assign weights1[12][64] = 16'b0000000000000111;
    assign weights1[12][65] = 16'b0000000000000011;
    assign weights1[12][66] = 16'b1111111111101101;
    assign weights1[12][67] = 16'b0000000000000011;
    assign weights1[12][68] = 16'b0000000000000110;
    assign weights1[12][69] = 16'b1111111111111110;
    assign weights1[12][70] = 16'b0000000000001000;
    assign weights1[12][71] = 16'b0000000000000111;
    assign weights1[12][72] = 16'b1111111111111001;
    assign weights1[12][73] = 16'b1111111111110010;
    assign weights1[12][74] = 16'b0000000000001110;
    assign weights1[12][75] = 16'b0000000000001100;
    assign weights1[12][76] = 16'b0000000000010001;
    assign weights1[12][77] = 16'b0000000000001111;
    assign weights1[12][78] = 16'b0000000000000010;
    assign weights1[12][79] = 16'b1111111111110100;
    assign weights1[12][80] = 16'b0000000000001010;
    assign weights1[12][81] = 16'b0000000000001010;
    assign weights1[12][82] = 16'b0000000000001001;
    assign weights1[12][83] = 16'b0000000000000110;
    assign weights1[12][84] = 16'b0000000000000010;
    assign weights1[12][85] = 16'b0000000000001101;
    assign weights1[12][86] = 16'b0000000000001011;
    assign weights1[12][87] = 16'b0000000000001111;
    assign weights1[12][88] = 16'b0000000000100000;
    assign weights1[12][89] = 16'b0000000000100000;
    assign weights1[12][90] = 16'b1111111111111111;
    assign weights1[12][91] = 16'b0000000000010011;
    assign weights1[12][92] = 16'b1111111111111100;
    assign weights1[12][93] = 16'b0000000000000011;
    assign weights1[12][94] = 16'b0000000000001010;
    assign weights1[12][95] = 16'b0000000000000110;
    assign weights1[12][96] = 16'b0000000000000001;
    assign weights1[12][97] = 16'b0000000000000111;
    assign weights1[12][98] = 16'b0000000000001010;
    assign weights1[12][99] = 16'b1111111111101011;
    assign weights1[12][100] = 16'b1111111111111101;
    assign weights1[12][101] = 16'b0000000000000110;
    assign weights1[12][102] = 16'b1111111111111100;
    assign weights1[12][103] = 16'b1111111111111111;
    assign weights1[12][104] = 16'b0000000000000011;
    assign weights1[12][105] = 16'b1111111111111100;
    assign weights1[12][106] = 16'b0000000000010000;
    assign weights1[12][107] = 16'b1111111111111001;
    assign weights1[12][108] = 16'b0000000000000110;
    assign weights1[12][109] = 16'b0000000000001011;
    assign weights1[12][110] = 16'b0000000000010101;
    assign weights1[12][111] = 16'b0000000000001110;
    assign weights1[12][112] = 16'b0000000000001000;
    assign weights1[12][113] = 16'b0000000000001101;
    assign weights1[12][114] = 16'b0000000000001110;
    assign weights1[12][115] = 16'b0000000000000111;
    assign weights1[12][116] = 16'b0000000000001101;
    assign weights1[12][117] = 16'b0000000000001100;
    assign weights1[12][118] = 16'b0000000000000011;
    assign weights1[12][119] = 16'b0000000000000000;
    assign weights1[12][120] = 16'b0000000000000110;
    assign weights1[12][121] = 16'b1111111111111110;
    assign weights1[12][122] = 16'b1111111111101011;
    assign weights1[12][123] = 16'b1111111111011110;
    assign weights1[12][124] = 16'b1111111111111101;
    assign weights1[12][125] = 16'b0000000000000101;
    assign weights1[12][126] = 16'b1111111111111110;
    assign weights1[12][127] = 16'b1111111111110010;
    assign weights1[12][128] = 16'b0000000000000000;
    assign weights1[12][129] = 16'b1111111111101101;
    assign weights1[12][130] = 16'b1111111111110110;
    assign weights1[12][131] = 16'b1111111111110111;
    assign weights1[12][132] = 16'b0000000000000011;
    assign weights1[12][133] = 16'b1111111111111010;
    assign weights1[12][134] = 16'b0000000000001010;
    assign weights1[12][135] = 16'b1111111111111010;
    assign weights1[12][136] = 16'b0000000000000001;
    assign weights1[12][137] = 16'b0000000000010110;
    assign weights1[12][138] = 16'b0000000000010001;
    assign weights1[12][139] = 16'b0000000000000101;
    assign weights1[12][140] = 16'b0000000000000010;
    assign weights1[12][141] = 16'b0000000000000010;
    assign weights1[12][142] = 16'b0000000000001000;
    assign weights1[12][143] = 16'b1111111111101100;
    assign weights1[12][144] = 16'b1111111111111011;
    assign weights1[12][145] = 16'b1111111111110100;
    assign weights1[12][146] = 16'b1111111111110100;
    assign weights1[12][147] = 16'b1111111111111011;
    assign weights1[12][148] = 16'b1111111111110111;
    assign weights1[12][149] = 16'b1111111111101101;
    assign weights1[12][150] = 16'b1111111111111000;
    assign weights1[12][151] = 16'b1111111111110100;
    assign weights1[12][152] = 16'b1111111111101100;
    assign weights1[12][153] = 16'b1111111111101100;
    assign weights1[12][154] = 16'b0000000000000001;
    assign weights1[12][155] = 16'b1111111111100000;
    assign weights1[12][156] = 16'b1111111111100111;
    assign weights1[12][157] = 16'b1111111111101101;
    assign weights1[12][158] = 16'b0000000000001001;
    assign weights1[12][159] = 16'b0000000000000010;
    assign weights1[12][160] = 16'b1111111111111000;
    assign weights1[12][161] = 16'b0000000000000111;
    assign weights1[12][162] = 16'b0000000000000000;
    assign weights1[12][163] = 16'b1111111111110000;
    assign weights1[12][164] = 16'b1111111111111101;
    assign weights1[12][165] = 16'b1111111111111110;
    assign weights1[12][166] = 16'b0000000000001100;
    assign weights1[12][167] = 16'b1111111111111101;
    assign weights1[12][168] = 16'b0000000000000100;
    assign weights1[12][169] = 16'b1111111111111100;
    assign weights1[12][170] = 16'b0000000000000001;
    assign weights1[12][171] = 16'b1111111111110000;
    assign weights1[12][172] = 16'b0000000000010010;
    assign weights1[12][173] = 16'b0000000000000101;
    assign weights1[12][174] = 16'b0000000000011111;
    assign weights1[12][175] = 16'b1111111111011111;
    assign weights1[12][176] = 16'b0000000000001011;
    assign weights1[12][177] = 16'b0000000000000110;
    assign weights1[12][178] = 16'b1111111111111111;
    assign weights1[12][179] = 16'b0000000000101000;
    assign weights1[12][180] = 16'b0000000000001011;
    assign weights1[12][181] = 16'b1111111111101100;
    assign weights1[12][182] = 16'b0000000000001001;
    assign weights1[12][183] = 16'b0000000000001000;
    assign weights1[12][184] = 16'b1111111111111010;
    assign weights1[12][185] = 16'b0000000000000110;
    assign weights1[12][186] = 16'b0000000000000010;
    assign weights1[12][187] = 16'b1111111111110010;
    assign weights1[12][188] = 16'b1111111111111111;
    assign weights1[12][189] = 16'b1111111111111110;
    assign weights1[12][190] = 16'b0000000000000010;
    assign weights1[12][191] = 16'b1111111111110111;
    assign weights1[12][192] = 16'b1111111111110101;
    assign weights1[12][193] = 16'b1111111111101011;
    assign weights1[12][194] = 16'b0000000000000010;
    assign weights1[12][195] = 16'b0000000000001001;
    assign weights1[12][196] = 16'b0000000000000010;
    assign weights1[12][197] = 16'b1111111111110101;
    assign weights1[12][198] = 16'b0000000000000001;
    assign weights1[12][199] = 16'b0000000000000100;
    assign weights1[12][200] = 16'b1111111111111010;
    assign weights1[12][201] = 16'b0000000000001010;
    assign weights1[12][202] = 16'b0000000000000111;
    assign weights1[12][203] = 16'b0000000000000010;
    assign weights1[12][204] = 16'b0000000000000110;
    assign weights1[12][205] = 16'b0000000000000111;
    assign weights1[12][206] = 16'b0000000000001000;
    assign weights1[12][207] = 16'b1111111111110000;
    assign weights1[12][208] = 16'b0000000000000101;
    assign weights1[12][209] = 16'b0000000000001110;
    assign weights1[12][210] = 16'b0000000000001001;
    assign weights1[12][211] = 16'b0000000000000010;
    assign weights1[12][212] = 16'b1111111111110100;
    assign weights1[12][213] = 16'b1111111111111001;
    assign weights1[12][214] = 16'b1111111111110111;
    assign weights1[12][215] = 16'b0000000000001111;
    assign weights1[12][216] = 16'b1111111111110111;
    assign weights1[12][217] = 16'b1111111111110111;
    assign weights1[12][218] = 16'b1111111111110001;
    assign weights1[12][219] = 16'b1111111111111111;
    assign weights1[12][220] = 16'b0000000000001001;
    assign weights1[12][221] = 16'b1111111111110111;
    assign weights1[12][222] = 16'b0000000000010000;
    assign weights1[12][223] = 16'b0000000000001111;
    assign weights1[12][224] = 16'b0000000000000010;
    assign weights1[12][225] = 16'b1111111111110110;
    assign weights1[12][226] = 16'b0000000000000010;
    assign weights1[12][227] = 16'b0000000000000100;
    assign weights1[12][228] = 16'b0000000000000001;
    assign weights1[12][229] = 16'b1111111111101111;
    assign weights1[12][230] = 16'b0000000000001001;
    assign weights1[12][231] = 16'b1111111111110111;
    assign weights1[12][232] = 16'b1111111111111011;
    assign weights1[12][233] = 16'b1111111111111011;
    assign weights1[12][234] = 16'b0000000000001101;
    assign weights1[12][235] = 16'b1111111111101111;
    assign weights1[12][236] = 16'b0000000000010000;
    assign weights1[12][237] = 16'b0000000000001000;
    assign weights1[12][238] = 16'b1111111111111100;
    assign weights1[12][239] = 16'b0000000000000101;
    assign weights1[12][240] = 16'b0000000000010100;
    assign weights1[12][241] = 16'b1111111111111100;
    assign weights1[12][242] = 16'b1111111111111100;
    assign weights1[12][243] = 16'b1111111111111110;
    assign weights1[12][244] = 16'b0000000000010110;
    assign weights1[12][245] = 16'b0000000000000000;
    assign weights1[12][246] = 16'b0000000000000100;
    assign weights1[12][247] = 16'b1111111111111111;
    assign weights1[12][248] = 16'b1111111111110111;
    assign weights1[12][249] = 16'b1111111111110100;
    assign weights1[12][250] = 16'b0000000000000001;
    assign weights1[12][251] = 16'b0000000000011000;
    assign weights1[12][252] = 16'b0000000000000100;
    assign weights1[12][253] = 16'b0000000000000000;
    assign weights1[12][254] = 16'b1111111111111010;
    assign weights1[12][255] = 16'b1111111111110101;
    assign weights1[12][256] = 16'b1111111111101000;
    assign weights1[12][257] = 16'b1111111111101010;
    assign weights1[12][258] = 16'b1111111111111110;
    assign weights1[12][259] = 16'b0000000000010000;
    assign weights1[12][260] = 16'b0000000000001001;
    assign weights1[12][261] = 16'b0000000000000010;
    assign weights1[12][262] = 16'b0000000000000000;
    assign weights1[12][263] = 16'b0000000000001011;
    assign weights1[12][264] = 16'b1111111111111111;
    assign weights1[12][265] = 16'b1111111111110011;
    assign weights1[12][266] = 16'b0000000000001111;
    assign weights1[12][267] = 16'b1111111111110100;
    assign weights1[12][268] = 16'b1111111111111101;
    assign weights1[12][269] = 16'b0000000000000000;
    assign weights1[12][270] = 16'b0000000000001000;
    assign weights1[12][271] = 16'b0000000000000101;
    assign weights1[12][272] = 16'b1111111111101110;
    assign weights1[12][273] = 16'b0000000000000001;
    assign weights1[12][274] = 16'b1111111111110111;
    assign weights1[12][275] = 16'b0000000000000010;
    assign weights1[12][276] = 16'b1111111111110001;
    assign weights1[12][277] = 16'b1111111111110100;
    assign weights1[12][278] = 16'b0000000000000001;
    assign weights1[12][279] = 16'b0000000000001000;
    assign weights1[12][280] = 16'b0000000000001000;
    assign weights1[12][281] = 16'b0000000000000111;
    assign weights1[12][282] = 16'b1111111111111100;
    assign weights1[12][283] = 16'b0000000000000111;
    assign weights1[12][284] = 16'b1111111111101001;
    assign weights1[12][285] = 16'b1111111111111000;
    assign weights1[12][286] = 16'b1111111111110110;
    assign weights1[12][287] = 16'b1111111111111001;
    assign weights1[12][288] = 16'b0000000000000010;
    assign weights1[12][289] = 16'b0000000000001101;
    assign weights1[12][290] = 16'b0000000000001101;
    assign weights1[12][291] = 16'b0000000000010001;
    assign weights1[12][292] = 16'b0000000000001100;
    assign weights1[12][293] = 16'b0000000000010110;
    assign weights1[12][294] = 16'b0000000000000000;
    assign weights1[12][295] = 16'b0000000000000111;
    assign weights1[12][296] = 16'b0000000000000011;
    assign weights1[12][297] = 16'b0000000000001100;
    assign weights1[12][298] = 16'b1111111111111111;
    assign weights1[12][299] = 16'b0000000000000011;
    assign weights1[12][300] = 16'b0000000000001110;
    assign weights1[12][301] = 16'b1111111111110110;
    assign weights1[12][302] = 16'b0000000000001010;
    assign weights1[12][303] = 16'b1111111111111000;
    assign weights1[12][304] = 16'b1111111111111101;
    assign weights1[12][305] = 16'b1111111111111100;
    assign weights1[12][306] = 16'b0000000000001001;
    assign weights1[12][307] = 16'b0000000000010100;
    assign weights1[12][308] = 16'b0000000000000000;
    assign weights1[12][309] = 16'b0000000000000001;
    assign weights1[12][310] = 16'b1111111111111100;
    assign weights1[12][311] = 16'b0000000000000110;
    assign weights1[12][312] = 16'b1111111111101010;
    assign weights1[12][313] = 16'b0000000000000100;
    assign weights1[12][314] = 16'b0000000000000001;
    assign weights1[12][315] = 16'b0000000000010110;
    assign weights1[12][316] = 16'b1111111111101110;
    assign weights1[12][317] = 16'b1111111111111001;
    assign weights1[12][318] = 16'b1111111111111010;
    assign weights1[12][319] = 16'b0000000000000000;
    assign weights1[12][320] = 16'b1111111111111111;
    assign weights1[12][321] = 16'b0000000000000011;
    assign weights1[12][322] = 16'b0000000000000110;
    assign weights1[12][323] = 16'b0000000000000001;
    assign weights1[12][324] = 16'b1111111111111001;
    assign weights1[12][325] = 16'b1111111111111000;
    assign weights1[12][326] = 16'b0000000000000000;
    assign weights1[12][327] = 16'b1111111111111010;
    assign weights1[12][328] = 16'b1111111111110101;
    assign weights1[12][329] = 16'b1111111111110100;
    assign weights1[12][330] = 16'b1111111111111001;
    assign weights1[12][331] = 16'b1111111111110101;
    assign weights1[12][332] = 16'b1111111111111101;
    assign weights1[12][333] = 16'b0000000000001000;
    assign weights1[12][334] = 16'b0000000000010101;
    assign weights1[12][335] = 16'b0000000000010100;
    assign weights1[12][336] = 16'b0000000000010010;
    assign weights1[12][337] = 16'b1111111111111001;
    assign weights1[12][338] = 16'b0000000000001101;
    assign weights1[12][339] = 16'b1111111111111000;
    assign weights1[12][340] = 16'b1111111111111101;
    assign weights1[12][341] = 16'b1111111111110010;
    assign weights1[12][342] = 16'b1111111111111011;
    assign weights1[12][343] = 16'b1111111111110100;
    assign weights1[12][344] = 16'b0000000000000010;
    assign weights1[12][345] = 16'b1111111111110100;
    assign weights1[12][346] = 16'b1111111111110010;
    assign weights1[12][347] = 16'b0000000000001010;
    assign weights1[12][348] = 16'b1111111111111010;
    assign weights1[12][349] = 16'b1111111111111110;
    assign weights1[12][350] = 16'b1111111111111011;
    assign weights1[12][351] = 16'b0000000000000001;
    assign weights1[12][352] = 16'b1111111111110101;
    assign weights1[12][353] = 16'b0000000000000101;
    assign weights1[12][354] = 16'b1111111111111101;
    assign weights1[12][355] = 16'b0000000000000111;
    assign weights1[12][356] = 16'b0000000000000100;
    assign weights1[12][357] = 16'b1111111111111011;
    assign weights1[12][358] = 16'b1111111111111100;
    assign weights1[12][359] = 16'b0000000000001100;
    assign weights1[12][360] = 16'b1111111111110010;
    assign weights1[12][361] = 16'b1111111111111110;
    assign weights1[12][362] = 16'b0000000000000011;
    assign weights1[12][363] = 16'b0000000000001000;
    assign weights1[12][364] = 16'b0000000000010111;
    assign weights1[12][365] = 16'b0000000000001001;
    assign weights1[12][366] = 16'b0000000000000101;
    assign weights1[12][367] = 16'b0000000000001110;
    assign weights1[12][368] = 16'b1111111111110110;
    assign weights1[12][369] = 16'b1111111111101011;
    assign weights1[12][370] = 16'b1111111111111011;
    assign weights1[12][371] = 16'b1111111111100000;
    assign weights1[12][372] = 16'b1111111111100110;
    assign weights1[12][373] = 16'b1111111111101100;
    assign weights1[12][374] = 16'b1111111111011001;
    assign weights1[12][375] = 16'b1111111111101000;
    assign weights1[12][376] = 16'b1111111111110100;
    assign weights1[12][377] = 16'b1111111111110010;
    assign weights1[12][378] = 16'b1111111111111100;
    assign weights1[12][379] = 16'b1111111111011111;
    assign weights1[12][380] = 16'b1111111111110110;
    assign weights1[12][381] = 16'b1111111111110001;
    assign weights1[12][382] = 16'b1111111111111111;
    assign weights1[12][383] = 16'b1111111111111100;
    assign weights1[12][384] = 16'b1111111111111110;
    assign weights1[12][385] = 16'b1111111111110111;
    assign weights1[12][386] = 16'b1111111111111000;
    assign weights1[12][387] = 16'b1111111111101000;
    assign weights1[12][388] = 16'b1111111111110101;
    assign weights1[12][389] = 16'b1111111111101010;
    assign weights1[12][390] = 16'b1111111111101010;
    assign weights1[12][391] = 16'b1111111111111100;
    assign weights1[12][392] = 16'b0000000000010000;
    assign weights1[12][393] = 16'b0000000000000011;
    assign weights1[12][394] = 16'b0000000000000010;
    assign weights1[12][395] = 16'b0000000000001000;
    assign weights1[12][396] = 16'b0000000000001100;
    assign weights1[12][397] = 16'b1111111111011000;
    assign weights1[12][398] = 16'b0000000000010011;
    assign weights1[12][399] = 16'b1111111111111011;
    assign weights1[12][400] = 16'b1111111111111010;
    assign weights1[12][401] = 16'b1111111111101111;
    assign weights1[12][402] = 16'b1111111111110101;
    assign weights1[12][403] = 16'b1111111111111101;
    assign weights1[12][404] = 16'b1111111111111010;
    assign weights1[12][405] = 16'b0000000000000100;
    assign weights1[12][406] = 16'b0000000000000110;
    assign weights1[12][407] = 16'b0000000000001111;
    assign weights1[12][408] = 16'b0000000000000010;
    assign weights1[12][409] = 16'b0000000000000101;
    assign weights1[12][410] = 16'b1111111111111101;
    assign weights1[12][411] = 16'b1111111111111011;
    assign weights1[12][412] = 16'b0000000000001101;
    assign weights1[12][413] = 16'b1111111111101101;
    assign weights1[12][414] = 16'b0000000000001001;
    assign weights1[12][415] = 16'b1111111111010101;
    assign weights1[12][416] = 16'b1111111111101100;
    assign weights1[12][417] = 16'b1111111111010001;
    assign weights1[12][418] = 16'b1111111111100101;
    assign weights1[12][419] = 16'b1111111111100110;
    assign weights1[12][420] = 16'b0000000000001011;
    assign weights1[12][421] = 16'b0000000000001010;
    assign weights1[12][422] = 16'b0000000000010100;
    assign weights1[12][423] = 16'b0000000000010001;
    assign weights1[12][424] = 16'b0000000000010011;
    assign weights1[12][425] = 16'b0000000000010011;
    assign weights1[12][426] = 16'b0000000000000111;
    assign weights1[12][427] = 16'b1111111111110110;
    assign weights1[12][428] = 16'b0000000000000111;
    assign weights1[12][429] = 16'b0000000000000000;
    assign weights1[12][430] = 16'b0000000000001100;
    assign weights1[12][431] = 16'b1111111111111111;
    assign weights1[12][432] = 16'b0000000000100000;
    assign weights1[12][433] = 16'b0000000000011001;
    assign weights1[12][434] = 16'b0000000000010011;
    assign weights1[12][435] = 16'b0000000000010000;
    assign weights1[12][436] = 16'b0000000000001111;
    assign weights1[12][437] = 16'b0000000000001110;
    assign weights1[12][438] = 16'b1111111111110101;
    assign weights1[12][439] = 16'b0000000000000010;
    assign weights1[12][440] = 16'b0000000000000101;
    assign weights1[12][441] = 16'b1111111111101101;
    assign weights1[12][442] = 16'b1111111111110010;
    assign weights1[12][443] = 16'b1111111111100111;
    assign weights1[12][444] = 16'b1111111111010001;
    assign weights1[12][445] = 16'b1111111111011111;
    assign weights1[12][446] = 16'b1111111111010111;
    assign weights1[12][447] = 16'b1111111111011011;
    assign weights1[12][448] = 16'b1111111111110111;
    assign weights1[12][449] = 16'b1111111111111011;
    assign weights1[12][450] = 16'b0000000000010110;
    assign weights1[12][451] = 16'b0000000000011101;
    assign weights1[12][452] = 16'b0000000000000001;
    assign weights1[12][453] = 16'b0000000000100111;
    assign weights1[12][454] = 16'b0000000000011111;
    assign weights1[12][455] = 16'b0000000000001000;
    assign weights1[12][456] = 16'b1111111111110111;
    assign weights1[12][457] = 16'b1111111111111001;
    assign weights1[12][458] = 16'b0000000000001100;
    assign weights1[12][459] = 16'b0000000000000101;
    assign weights1[12][460] = 16'b0000000000000110;
    assign weights1[12][461] = 16'b0000000000001101;
    assign weights1[12][462] = 16'b0000000000010100;
    assign weights1[12][463] = 16'b1111111111111111;
    assign weights1[12][464] = 16'b0000000000001011;
    assign weights1[12][465] = 16'b1111111111111100;
    assign weights1[12][466] = 16'b0000000000001111;
    assign weights1[12][467] = 16'b1111111111110001;
    assign weights1[12][468] = 16'b1111111111111010;
    assign weights1[12][469] = 16'b1111111111011000;
    assign weights1[12][470] = 16'b1111111111010110;
    assign weights1[12][471] = 16'b1111111111010111;
    assign weights1[12][472] = 16'b1111111111011111;
    assign weights1[12][473] = 16'b1111111111101001;
    assign weights1[12][474] = 16'b1111111111101111;
    assign weights1[12][475] = 16'b1111111111101101;
    assign weights1[12][476] = 16'b1111111111100011;
    assign weights1[12][477] = 16'b1111111111110001;
    assign weights1[12][478] = 16'b0000000000000011;
    assign weights1[12][479] = 16'b0000000000000110;
    assign weights1[12][480] = 16'b0000000000000100;
    assign weights1[12][481] = 16'b1111111111111111;
    assign weights1[12][482] = 16'b1111111111111011;
    assign weights1[12][483] = 16'b0000000000001000;
    assign weights1[12][484] = 16'b0000000000010011;
    assign weights1[12][485] = 16'b0000000000001111;
    assign weights1[12][486] = 16'b0000000000010011;
    assign weights1[12][487] = 16'b1111111111110110;
    assign weights1[12][488] = 16'b0000000000010111;
    assign weights1[12][489] = 16'b0000000000011100;
    assign weights1[12][490] = 16'b0000000000011110;
    assign weights1[12][491] = 16'b0000000000010001;
    assign weights1[12][492] = 16'b1111111111111110;
    assign weights1[12][493] = 16'b1111111111111111;
    assign weights1[12][494] = 16'b1111111111111100;
    assign weights1[12][495] = 16'b1111111111101110;
    assign weights1[12][496] = 16'b1111111111011111;
    assign weights1[12][497] = 16'b1111111111010101;
    assign weights1[12][498] = 16'b1111111111100101;
    assign weights1[12][499] = 16'b1111111111101010;
    assign weights1[12][500] = 16'b1111111111111111;
    assign weights1[12][501] = 16'b0000000000010011;
    assign weights1[12][502] = 16'b1111111111111001;
    assign weights1[12][503] = 16'b0000000000001100;
    assign weights1[12][504] = 16'b1111111111011011;
    assign weights1[12][505] = 16'b1111111111000111;
    assign weights1[12][506] = 16'b1111111111010101;
    assign weights1[12][507] = 16'b1111111111100011;
    assign weights1[12][508] = 16'b1111111111101010;
    assign weights1[12][509] = 16'b0000000000001100;
    assign weights1[12][510] = 16'b0000000000000110;
    assign weights1[12][511] = 16'b1111111111111011;
    assign weights1[12][512] = 16'b1111111111111100;
    assign weights1[12][513] = 16'b1111111111111101;
    assign weights1[12][514] = 16'b0000000000001100;
    assign weights1[12][515] = 16'b1111111111111100;
    assign weights1[12][516] = 16'b0000000000100011;
    assign weights1[12][517] = 16'b0000000000100000;
    assign weights1[12][518] = 16'b0000000000001000;
    assign weights1[12][519] = 16'b0000000000010111;
    assign weights1[12][520] = 16'b0000000000000111;
    assign weights1[12][521] = 16'b1111111111101011;
    assign weights1[12][522] = 16'b1111111111100010;
    assign weights1[12][523] = 16'b1111111111010011;
    assign weights1[12][524] = 16'b1111111111010111;
    assign weights1[12][525] = 16'b1111111111100101;
    assign weights1[12][526] = 16'b1111111111110000;
    assign weights1[12][527] = 16'b0000000000001010;
    assign weights1[12][528] = 16'b0000000000000010;
    assign weights1[12][529] = 16'b0000000000100000;
    assign weights1[12][530] = 16'b0000000000011001;
    assign weights1[12][531] = 16'b0000000000000100;
    assign weights1[12][532] = 16'b1111111111011000;
    assign weights1[12][533] = 16'b1111111111000011;
    assign weights1[12][534] = 16'b1111111110111110;
    assign weights1[12][535] = 16'b1111111110110010;
    assign weights1[12][536] = 16'b1111111110111010;
    assign weights1[12][537] = 16'b1111111111100000;
    assign weights1[12][538] = 16'b1111111111101111;
    assign weights1[12][539] = 16'b1111111111111000;
    assign weights1[12][540] = 16'b0000000000000101;
    assign weights1[12][541] = 16'b0000000000001001;
    assign weights1[12][542] = 16'b1111111111111001;
    assign weights1[12][543] = 16'b0000000000001010;
    assign weights1[12][544] = 16'b1111111111110010;
    assign weights1[12][545] = 16'b0000000000001010;
    assign weights1[12][546] = 16'b1111111111111100;
    assign weights1[12][547] = 16'b1111111111100001;
    assign weights1[12][548] = 16'b1111111111001110;
    assign weights1[12][549] = 16'b1111111111010010;
    assign weights1[12][550] = 16'b1111111111011011;
    assign weights1[12][551] = 16'b1111111111010111;
    assign weights1[12][552] = 16'b1111111111100010;
    assign weights1[12][553] = 16'b1111111111110100;
    assign weights1[12][554] = 16'b0000000000001011;
    assign weights1[12][555] = 16'b0000000000010101;
    assign weights1[12][556] = 16'b0000000000010001;
    assign weights1[12][557] = 16'b0000000000100001;
    assign weights1[12][558] = 16'b0000000000011000;
    assign weights1[12][559] = 16'b0000000000001010;
    assign weights1[12][560] = 16'b1111111111011000;
    assign weights1[12][561] = 16'b1111111110111011;
    assign weights1[12][562] = 16'b1111111110101110;
    assign weights1[12][563] = 16'b1111111110011101;
    assign weights1[12][564] = 16'b1111111110000111;
    assign weights1[12][565] = 16'b1111111110000100;
    assign weights1[12][566] = 16'b1111111101100001;
    assign weights1[12][567] = 16'b1111111101011101;
    assign weights1[12][568] = 16'b1111111101001111;
    assign weights1[12][569] = 16'b1111111101101101;
    assign weights1[12][570] = 16'b1111111110000100;
    assign weights1[12][571] = 16'b1111111101110010;
    assign weights1[12][572] = 16'b1111111101010100;
    assign weights1[12][573] = 16'b1111111101111011;
    assign weights1[12][574] = 16'b1111111110001000;
    assign weights1[12][575] = 16'b1111111110100000;
    assign weights1[12][576] = 16'b1111111111001000;
    assign weights1[12][577] = 16'b1111111111010101;
    assign weights1[12][578] = 16'b1111111111101011;
    assign weights1[12][579] = 16'b1111111111111101;
    assign weights1[12][580] = 16'b0000000000001111;
    assign weights1[12][581] = 16'b0000000000010010;
    assign weights1[12][582] = 16'b0000000000010100;
    assign weights1[12][583] = 16'b0000000000010111;
    assign weights1[12][584] = 16'b0000000000011001;
    assign weights1[12][585] = 16'b0000000000011001;
    assign weights1[12][586] = 16'b0000000000010010;
    assign weights1[12][587] = 16'b0000000000001100;
    assign weights1[12][588] = 16'b1111111111011111;
    assign weights1[12][589] = 16'b1111111111000101;
    assign weights1[12][590] = 16'b1111111110101011;
    assign weights1[12][591] = 16'b1111111110101010;
    assign weights1[12][592] = 16'b1111111110011110;
    assign weights1[12][593] = 16'b1111111110100010;
    assign weights1[12][594] = 16'b1111111110000100;
    assign weights1[12][595] = 16'b1111111101101101;
    assign weights1[12][596] = 16'b1111111100110010;
    assign weights1[12][597] = 16'b1111111100100111;
    assign weights1[12][598] = 16'b1111111100011100;
    assign weights1[12][599] = 16'b1111111011111001;
    assign weights1[12][600] = 16'b1111111100010001;
    assign weights1[12][601] = 16'b1111111101000010;
    assign weights1[12][602] = 16'b1111111110000001;
    assign weights1[12][603] = 16'b1111111110110100;
    assign weights1[12][604] = 16'b1111111111100001;
    assign weights1[12][605] = 16'b1111111111011101;
    assign weights1[12][606] = 16'b0000000000000011;
    assign weights1[12][607] = 16'b0000000000011100;
    assign weights1[12][608] = 16'b0000000000000100;
    assign weights1[12][609] = 16'b0000000000010110;
    assign weights1[12][610] = 16'b0000000000110000;
    assign weights1[12][611] = 16'b0000000000101000;
    assign weights1[12][612] = 16'b0000000000010101;
    assign weights1[12][613] = 16'b0000000000011000;
    assign weights1[12][614] = 16'b0000000000010010;
    assign weights1[12][615] = 16'b0000000000001011;
    assign weights1[12][616] = 16'b1111111111100111;
    assign weights1[12][617] = 16'b1111111111001101;
    assign weights1[12][618] = 16'b1111111111000011;
    assign weights1[12][619] = 16'b1111111111000100;
    assign weights1[12][620] = 16'b1111111110111101;
    assign weights1[12][621] = 16'b1111111110111000;
    assign weights1[12][622] = 16'b1111111110110101;
    assign weights1[12][623] = 16'b1111111111000001;
    assign weights1[12][624] = 16'b1111111110110011;
    assign weights1[12][625] = 16'b1111111110001001;
    assign weights1[12][626] = 16'b1111111110001001;
    assign weights1[12][627] = 16'b1111111110101011;
    assign weights1[12][628] = 16'b1111111110111110;
    assign weights1[12][629] = 16'b1111111111010100;
    assign weights1[12][630] = 16'b1111111111011111;
    assign weights1[12][631] = 16'b1111111111100000;
    assign weights1[12][632] = 16'b0000000000000000;
    assign weights1[12][633] = 16'b0000000000001100;
    assign weights1[12][634] = 16'b0000000000011101;
    assign weights1[12][635] = 16'b1111111111111101;
    assign weights1[12][636] = 16'b0000000000010010;
    assign weights1[12][637] = 16'b0000000000010000;
    assign weights1[12][638] = 16'b0000000000011010;
    assign weights1[12][639] = 16'b0000000000011001;
    assign weights1[12][640] = 16'b0000000000010011;
    assign weights1[12][641] = 16'b0000000000001101;
    assign weights1[12][642] = 16'b0000000000001010;
    assign weights1[12][643] = 16'b0000000000010010;
    assign weights1[12][644] = 16'b1111111111111010;
    assign weights1[12][645] = 16'b1111111111101000;
    assign weights1[12][646] = 16'b1111111111011101;
    assign weights1[12][647] = 16'b1111111111101000;
    assign weights1[12][648] = 16'b1111111111110010;
    assign weights1[12][649] = 16'b1111111111010111;
    assign weights1[12][650] = 16'b1111111111100010;
    assign weights1[12][651] = 16'b1111111111111101;
    assign weights1[12][652] = 16'b0000000000000001;
    assign weights1[12][653] = 16'b1111111111111101;
    assign weights1[12][654] = 16'b0000000000011000;
    assign weights1[12][655] = 16'b0000000000101000;
    assign weights1[12][656] = 16'b0000000001001010;
    assign weights1[12][657] = 16'b0000000001001001;
    assign weights1[12][658] = 16'b0000000000110100;
    assign weights1[12][659] = 16'b0000000001000001;
    assign weights1[12][660] = 16'b0000000000011010;
    assign weights1[12][661] = 16'b0000000000010010;
    assign weights1[12][662] = 16'b0000000000001111;
    assign weights1[12][663] = 16'b0000000000100110;
    assign weights1[12][664] = 16'b0000000000001101;
    assign weights1[12][665] = 16'b0000000000010010;
    assign weights1[12][666] = 16'b0000000000001100;
    assign weights1[12][667] = 16'b1111111111110001;
    assign weights1[12][668] = 16'b0000000000011101;
    assign weights1[12][669] = 16'b0000000000000111;
    assign weights1[12][670] = 16'b0000000000001011;
    assign weights1[12][671] = 16'b0000000000001100;
    assign weights1[12][672] = 16'b0000000000000001;
    assign weights1[12][673] = 16'b0000000000000111;
    assign weights1[12][674] = 16'b1111111111101101;
    assign weights1[12][675] = 16'b1111111111110101;
    assign weights1[12][676] = 16'b0000000000000011;
    assign weights1[12][677] = 16'b0000000000010010;
    assign weights1[12][678] = 16'b1111111111111101;
    assign weights1[12][679] = 16'b0000000000010010;
    assign weights1[12][680] = 16'b0000000000110100;
    assign weights1[12][681] = 16'b0000000001100011;
    assign weights1[12][682] = 16'b0000000001101110;
    assign weights1[12][683] = 16'b0000000010000100;
    assign weights1[12][684] = 16'b0000000001001000;
    assign weights1[12][685] = 16'b0000000000101000;
    assign weights1[12][686] = 16'b0000000000101111;
    assign weights1[12][687] = 16'b0000000000110111;
    assign weights1[12][688] = 16'b0000000000001010;
    assign weights1[12][689] = 16'b0000000000010011;
    assign weights1[12][690] = 16'b0000000000001111;
    assign weights1[12][691] = 16'b0000000000011101;
    assign weights1[12][692] = 16'b0000000000010011;
    assign weights1[12][693] = 16'b0000000000000000;
    assign weights1[12][694] = 16'b0000000000001011;
    assign weights1[12][695] = 16'b0000000000011000;
    assign weights1[12][696] = 16'b0000000000001100;
    assign weights1[12][697] = 16'b0000000000000010;
    assign weights1[12][698] = 16'b0000000000000010;
    assign weights1[12][699] = 16'b1111111111111111;
    assign weights1[12][700] = 16'b1111111111111111;
    assign weights1[12][701] = 16'b1111111111111111;
    assign weights1[12][702] = 16'b0000000000010010;
    assign weights1[12][703] = 16'b0000000000011011;
    assign weights1[12][704] = 16'b0000000000011011;
    assign weights1[12][705] = 16'b0000000000101101;
    assign weights1[12][706] = 16'b0000000001010010;
    assign weights1[12][707] = 16'b0000000001000100;
    assign weights1[12][708] = 16'b0000000001011111;
    assign weights1[12][709] = 16'b0000000000111111;
    assign weights1[12][710] = 16'b0000000001101100;
    assign weights1[12][711] = 16'b0000000000110000;
    assign weights1[12][712] = 16'b0000000000110100;
    assign weights1[12][713] = 16'b0000000000101001;
    assign weights1[12][714] = 16'b0000000000001110;
    assign weights1[12][715] = 16'b0000000000011001;
    assign weights1[12][716] = 16'b0000000000010001;
    assign weights1[12][717] = 16'b0000000000001110;
    assign weights1[12][718] = 16'b0000000000001111;
    assign weights1[12][719] = 16'b0000000000100011;
    assign weights1[12][720] = 16'b0000000000001010;
    assign weights1[12][721] = 16'b0000000000001011;
    assign weights1[12][722] = 16'b0000000000001111;
    assign weights1[12][723] = 16'b0000000000100000;
    assign weights1[12][724] = 16'b0000000000100001;
    assign weights1[12][725] = 16'b0000000000000001;
    assign weights1[12][726] = 16'b0000000000000111;
    assign weights1[12][727] = 16'b0000000000000010;
    assign weights1[12][728] = 16'b1111111111111101;
    assign weights1[12][729] = 16'b0000000000000111;
    assign weights1[12][730] = 16'b0000000000010011;
    assign weights1[12][731] = 16'b0000000000011011;
    assign weights1[12][732] = 16'b0000000000011101;
    assign weights1[12][733] = 16'b0000000000101100;
    assign weights1[12][734] = 16'b0000000001001111;
    assign weights1[12][735] = 16'b0000000001010110;
    assign weights1[12][736] = 16'b0000000001001000;
    assign weights1[12][737] = 16'b0000000000011001;
    assign weights1[12][738] = 16'b0000000000010101;
    assign weights1[12][739] = 16'b0000000000000111;
    assign weights1[12][740] = 16'b0000000000000100;
    assign weights1[12][741] = 16'b0000000000011001;
    assign weights1[12][742] = 16'b0000000000001001;
    assign weights1[12][743] = 16'b0000000000011000;
    assign weights1[12][744] = 16'b0000000000000110;
    assign weights1[12][745] = 16'b0000000000001001;
    assign weights1[12][746] = 16'b0000000000001111;
    assign weights1[12][747] = 16'b0000000000000010;
    assign weights1[12][748] = 16'b0000000000010000;
    assign weights1[12][749] = 16'b0000000000000010;
    assign weights1[12][750] = 16'b1111111111111110;
    assign weights1[12][751] = 16'b1111111111111011;
    assign weights1[12][752] = 16'b0000000000001001;
    assign weights1[12][753] = 16'b0000000000001011;
    assign weights1[12][754] = 16'b0000000000000100;
    assign weights1[12][755] = 16'b1111111111111111;
    assign weights1[12][756] = 16'b0000000000000011;
    assign weights1[12][757] = 16'b0000000000001101;
    assign weights1[12][758] = 16'b0000000000011000;
    assign weights1[12][759] = 16'b0000000000011111;
    assign weights1[12][760] = 16'b0000000000101010;
    assign weights1[12][761] = 16'b0000000000110111;
    assign weights1[12][762] = 16'b0000000000111110;
    assign weights1[12][763] = 16'b0000000001000001;
    assign weights1[12][764] = 16'b0000000000101010;
    assign weights1[12][765] = 16'b0000000000100100;
    assign weights1[12][766] = 16'b0000000000101011;
    assign weights1[12][767] = 16'b0000000000100110;
    assign weights1[12][768] = 16'b0000000000110010;
    assign weights1[12][769] = 16'b0000000000100000;
    assign weights1[12][770] = 16'b0000000000101000;
    assign weights1[12][771] = 16'b0000000000010011;
    assign weights1[12][772] = 16'b0000000000011000;
    assign weights1[12][773] = 16'b0000000000000111;
    assign weights1[12][774] = 16'b0000000000010111;
    assign weights1[12][775] = 16'b0000000000000111;
    assign weights1[12][776] = 16'b0000000000000001;
    assign weights1[12][777] = 16'b0000000000001010;
    assign weights1[12][778] = 16'b0000000000001110;
    assign weights1[12][779] = 16'b0000000000010011;
    assign weights1[12][780] = 16'b0000000000001000;
    assign weights1[12][781] = 16'b0000000000000110;
    assign weights1[12][782] = 16'b1111111111111100;
    assign weights1[12][783] = 16'b1111111111111100;
    assign weights1[13][0] = 16'b0000000000000001;
    assign weights1[13][1] = 16'b0000000000000000;
    assign weights1[13][2] = 16'b0000000000000010;
    assign weights1[13][3] = 16'b0000000000000100;
    assign weights1[13][4] = 16'b0000000000001010;
    assign weights1[13][5] = 16'b0000000000000101;
    assign weights1[13][6] = 16'b0000000000000111;
    assign weights1[13][7] = 16'b0000000000001011;
    assign weights1[13][8] = 16'b0000000000001101;
    assign weights1[13][9] = 16'b0000000000001010;
    assign weights1[13][10] = 16'b0000000000011101;
    assign weights1[13][11] = 16'b0000000000010011;
    assign weights1[13][12] = 16'b1111111111111110;
    assign weights1[13][13] = 16'b0000000000000001;
    assign weights1[13][14] = 16'b1111111111111110;
    assign weights1[13][15] = 16'b0000000000010000;
    assign weights1[13][16] = 16'b0000000000000101;
    assign weights1[13][17] = 16'b0000000000000011;
    assign weights1[13][18] = 16'b0000000000000010;
    assign weights1[13][19] = 16'b0000000000001100;
    assign weights1[13][20] = 16'b0000000000000001;
    assign weights1[13][21] = 16'b0000000000000110;
    assign weights1[13][22] = 16'b1111111111111100;
    assign weights1[13][23] = 16'b0000000000010101;
    assign weights1[13][24] = 16'b0000000000010000;
    assign weights1[13][25] = 16'b0000000000001011;
    assign weights1[13][26] = 16'b0000000000000100;
    assign weights1[13][27] = 16'b0000000000000010;
    assign weights1[13][28] = 16'b0000000000000001;
    assign weights1[13][29] = 16'b0000000000000001;
    assign weights1[13][30] = 16'b0000000000000100;
    assign weights1[13][31] = 16'b0000000000000100;
    assign weights1[13][32] = 16'b0000000000010010;
    assign weights1[13][33] = 16'b0000000000010010;
    assign weights1[13][34] = 16'b0000000000010011;
    assign weights1[13][35] = 16'b0000000000000011;
    assign weights1[13][36] = 16'b0000000000000010;
    assign weights1[13][37] = 16'b0000000000001101;
    assign weights1[13][38] = 16'b0000000000001001;
    assign weights1[13][39] = 16'b1111111111111110;
    assign weights1[13][40] = 16'b0000000000001100;
    assign weights1[13][41] = 16'b0000000000001100;
    assign weights1[13][42] = 16'b1111111111111101;
    assign weights1[13][43] = 16'b0000000000000000;
    assign weights1[13][44] = 16'b0000000000001010;
    assign weights1[13][45] = 16'b0000000000000100;
    assign weights1[13][46] = 16'b1111111111110111;
    assign weights1[13][47] = 16'b0000000000001001;
    assign weights1[13][48] = 16'b0000000000000110;
    assign weights1[13][49] = 16'b1111111111111111;
    assign weights1[13][50] = 16'b0000000000000110;
    assign weights1[13][51] = 16'b0000000000000010;
    assign weights1[13][52] = 16'b0000000000001010;
    assign weights1[13][53] = 16'b0000000000000010;
    assign weights1[13][54] = 16'b1111111111111111;
    assign weights1[13][55] = 16'b0000000000000001;
    assign weights1[13][56] = 16'b0000000000000010;
    assign weights1[13][57] = 16'b0000000000000101;
    assign weights1[13][58] = 16'b0000000000000100;
    assign weights1[13][59] = 16'b0000000000000100;
    assign weights1[13][60] = 16'b0000000000000101;
    assign weights1[13][61] = 16'b1111111111111011;
    assign weights1[13][62] = 16'b0000000000010000;
    assign weights1[13][63] = 16'b0000000000010111;
    assign weights1[13][64] = 16'b0000000000001010;
    assign weights1[13][65] = 16'b0000000000011000;
    assign weights1[13][66] = 16'b0000000000010011;
    assign weights1[13][67] = 16'b0000000000001010;
    assign weights1[13][68] = 16'b0000000000001010;
    assign weights1[13][69] = 16'b0000000000000101;
    assign weights1[13][70] = 16'b0000000000000001;
    assign weights1[13][71] = 16'b0000000000001000;
    assign weights1[13][72] = 16'b0000000000001000;
    assign weights1[13][73] = 16'b1111111111111111;
    assign weights1[13][74] = 16'b1111111111111000;
    assign weights1[13][75] = 16'b0000000000000111;
    assign weights1[13][76] = 16'b0000000000000011;
    assign weights1[13][77] = 16'b0000000000001010;
    assign weights1[13][78] = 16'b0000000000000001;
    assign weights1[13][79] = 16'b1111111111111011;
    assign weights1[13][80] = 16'b1111111111111100;
    assign weights1[13][81] = 16'b0000000000000001;
    assign weights1[13][82] = 16'b0000000000000101;
    assign weights1[13][83] = 16'b0000000000000111;
    assign weights1[13][84] = 16'b0000000000000011;
    assign weights1[13][85] = 16'b0000000000000111;
    assign weights1[13][86] = 16'b0000000000001101;
    assign weights1[13][87] = 16'b0000000000001011;
    assign weights1[13][88] = 16'b0000000000000101;
    assign weights1[13][89] = 16'b0000000000001111;
    assign weights1[13][90] = 16'b0000000000001010;
    assign weights1[13][91] = 16'b0000000000010001;
    assign weights1[13][92] = 16'b1111111111111001;
    assign weights1[13][93] = 16'b1111111111110111;
    assign weights1[13][94] = 16'b0000000000000000;
    assign weights1[13][95] = 16'b0000000000010100;
    assign weights1[13][96] = 16'b0000000000000100;
    assign weights1[13][97] = 16'b1111111111101111;
    assign weights1[13][98] = 16'b0000000000001010;
    assign weights1[13][99] = 16'b0000000000000100;
    assign weights1[13][100] = 16'b1111111111110110;
    assign weights1[13][101] = 16'b0000000000000001;
    assign weights1[13][102] = 16'b1111111111110100;
    assign weights1[13][103] = 16'b1111111111110111;
    assign weights1[13][104] = 16'b0000000000001001;
    assign weights1[13][105] = 16'b0000000000000010;
    assign weights1[13][106] = 16'b1111111111111101;
    assign weights1[13][107] = 16'b0000000000001101;
    assign weights1[13][108] = 16'b1111111111111011;
    assign weights1[13][109] = 16'b0000000000001101;
    assign weights1[13][110] = 16'b0000000000001111;
    assign weights1[13][111] = 16'b0000000000001101;
    assign weights1[13][112] = 16'b0000000000000111;
    assign weights1[13][113] = 16'b0000000000001000;
    assign weights1[13][114] = 16'b0000000000010010;
    assign weights1[13][115] = 16'b0000000000000001;
    assign weights1[13][116] = 16'b0000000000000001;
    assign weights1[13][117] = 16'b0000000000000010;
    assign weights1[13][118] = 16'b1111111111101110;
    assign weights1[13][119] = 16'b0000000000001101;
    assign weights1[13][120] = 16'b0000000000000111;
    assign weights1[13][121] = 16'b1111111111101111;
    assign weights1[13][122] = 16'b0000000000000001;
    assign weights1[13][123] = 16'b1111111111110111;
    assign weights1[13][124] = 16'b0000000000000011;
    assign weights1[13][125] = 16'b0000000000001000;
    assign weights1[13][126] = 16'b0000000000000101;
    assign weights1[13][127] = 16'b0000000000000010;
    assign weights1[13][128] = 16'b0000000000001001;
    assign weights1[13][129] = 16'b0000000000000101;
    assign weights1[13][130] = 16'b0000000000010011;
    assign weights1[13][131] = 16'b0000000000010001;
    assign weights1[13][132] = 16'b1111111111111110;
    assign weights1[13][133] = 16'b0000000000000001;
    assign weights1[13][134] = 16'b1111111111111001;
    assign weights1[13][135] = 16'b1111111111111011;
    assign weights1[13][136] = 16'b0000000000001100;
    assign weights1[13][137] = 16'b0000000000000100;
    assign weights1[13][138] = 16'b1111111111111111;
    assign weights1[13][139] = 16'b0000000000000100;
    assign weights1[13][140] = 16'b0000000000001001;
    assign weights1[13][141] = 16'b0000000000001010;
    assign weights1[13][142] = 16'b0000000000010001;
    assign weights1[13][143] = 16'b0000000000000010;
    assign weights1[13][144] = 16'b1111111111111110;
    assign weights1[13][145] = 16'b0000000000000010;
    assign weights1[13][146] = 16'b1111111111111100;
    assign weights1[13][147] = 16'b1111111111111010;
    assign weights1[13][148] = 16'b0000000000000100;
    assign weights1[13][149] = 16'b0000000000000001;
    assign weights1[13][150] = 16'b0000000000000011;
    assign weights1[13][151] = 16'b0000000000000011;
    assign weights1[13][152] = 16'b0000000000010011;
    assign weights1[13][153] = 16'b0000000000000011;
    assign weights1[13][154] = 16'b1111111111111011;
    assign weights1[13][155] = 16'b0000000000000010;
    assign weights1[13][156] = 16'b0000000000001100;
    assign weights1[13][157] = 16'b1111111111110110;
    assign weights1[13][158] = 16'b1111111111110001;
    assign weights1[13][159] = 16'b0000000000000100;
    assign weights1[13][160] = 16'b1111111111111101;
    assign weights1[13][161] = 16'b1111111111111111;
    assign weights1[13][162] = 16'b1111111111100001;
    assign weights1[13][163] = 16'b0000000000100110;
    assign weights1[13][164] = 16'b0000000000000001;
    assign weights1[13][165] = 16'b1111111111101001;
    assign weights1[13][166] = 16'b1111111111110010;
    assign weights1[13][167] = 16'b0000000000000110;
    assign weights1[13][168] = 16'b0000000000000111;
    assign weights1[13][169] = 16'b0000000000000011;
    assign weights1[13][170] = 16'b0000000000000010;
    assign weights1[13][171] = 16'b0000000000000101;
    assign weights1[13][172] = 16'b1111111111101100;
    assign weights1[13][173] = 16'b1111111111101101;
    assign weights1[13][174] = 16'b0000000000001010;
    assign weights1[13][175] = 16'b1111111111101100;
    assign weights1[13][176] = 16'b1111111111111111;
    assign weights1[13][177] = 16'b1111111111111110;
    assign weights1[13][178] = 16'b0000000000000010;
    assign weights1[13][179] = 16'b0000000000001100;
    assign weights1[13][180] = 16'b1111111111101100;
    assign weights1[13][181] = 16'b1111111111111001;
    assign weights1[13][182] = 16'b1111111111111110;
    assign weights1[13][183] = 16'b1111111111111011;
    assign weights1[13][184] = 16'b0000000000001011;
    assign weights1[13][185] = 16'b1111111111111110;
    assign weights1[13][186] = 16'b0000000000010000;
    assign weights1[13][187] = 16'b0000000000000100;
    assign weights1[13][188] = 16'b0000000000000011;
    assign weights1[13][189] = 16'b0000000000000110;
    assign weights1[13][190] = 16'b0000000000000101;
    assign weights1[13][191] = 16'b1111111111110100;
    assign weights1[13][192] = 16'b1111111111111001;
    assign weights1[13][193] = 16'b1111111111110011;
    assign weights1[13][194] = 16'b0000000000010101;
    assign weights1[13][195] = 16'b0000000000000111;
    assign weights1[13][196] = 16'b1111111111111110;
    assign weights1[13][197] = 16'b1111111111110111;
    assign weights1[13][198] = 16'b1111111111110000;
    assign weights1[13][199] = 16'b1111111111101101;
    assign weights1[13][200] = 16'b1111111111110101;
    assign weights1[13][201] = 16'b0000000000001101;
    assign weights1[13][202] = 16'b1111111111101111;
    assign weights1[13][203] = 16'b0000000000010110;
    assign weights1[13][204] = 16'b1111111111111100;
    assign weights1[13][205] = 16'b1111111111110010;
    assign weights1[13][206] = 16'b1111111111110110;
    assign weights1[13][207] = 16'b0000000000001111;
    assign weights1[13][208] = 16'b0000000000010000;
    assign weights1[13][209] = 16'b0000000000000110;
    assign weights1[13][210] = 16'b0000000000010101;
    assign weights1[13][211] = 16'b0000000000001000;
    assign weights1[13][212] = 16'b0000000000001000;
    assign weights1[13][213] = 16'b0000000000011010;
    assign weights1[13][214] = 16'b0000000000001010;
    assign weights1[13][215] = 16'b0000000000010001;
    assign weights1[13][216] = 16'b0000000000001110;
    assign weights1[13][217] = 16'b1111111111111101;
    assign weights1[13][218] = 16'b0000000000000100;
    assign weights1[13][219] = 16'b0000000000000010;
    assign weights1[13][220] = 16'b0000000000000111;
    assign weights1[13][221] = 16'b1111111111111100;
    assign weights1[13][222] = 16'b1111111111110111;
    assign weights1[13][223] = 16'b0000000000000101;
    assign weights1[13][224] = 16'b1111111111111110;
    assign weights1[13][225] = 16'b1111111111110001;
    assign weights1[13][226] = 16'b0000000000000001;
    assign weights1[13][227] = 16'b1111111111101001;
    assign weights1[13][228] = 16'b1111111111111001;
    assign weights1[13][229] = 16'b0000000000000011;
    assign weights1[13][230] = 16'b1111111111110111;
    assign weights1[13][231] = 16'b1111111111110111;
    assign weights1[13][232] = 16'b1111111111110100;
    assign weights1[13][233] = 16'b0000000000001000;
    assign weights1[13][234] = 16'b1111111111111111;
    assign weights1[13][235] = 16'b0000000000000110;
    assign weights1[13][236] = 16'b0000000000000101;
    assign weights1[13][237] = 16'b1111111111111000;
    assign weights1[13][238] = 16'b0000000000000101;
    assign weights1[13][239] = 16'b0000000000000101;
    assign weights1[13][240] = 16'b0000000000001010;
    assign weights1[13][241] = 16'b1111111111111100;
    assign weights1[13][242] = 16'b1111111111111011;
    assign weights1[13][243] = 16'b0000000000000010;
    assign weights1[13][244] = 16'b0000000000001111;
    assign weights1[13][245] = 16'b0000000000010011;
    assign weights1[13][246] = 16'b0000000000001011;
    assign weights1[13][247] = 16'b0000000000010000;
    assign weights1[13][248] = 16'b0000000000011000;
    assign weights1[13][249] = 16'b0000000000000101;
    assign weights1[13][250] = 16'b1111111111111000;
    assign weights1[13][251] = 16'b0000000000000011;
    assign weights1[13][252] = 16'b1111111111110110;
    assign weights1[13][253] = 16'b1111111111101011;
    assign weights1[13][254] = 16'b1111111111101011;
    assign weights1[13][255] = 16'b1111111111110001;
    assign weights1[13][256] = 16'b0000000000000000;
    assign weights1[13][257] = 16'b0000000000001100;
    assign weights1[13][258] = 16'b0000000000000000;
    assign weights1[13][259] = 16'b0000000000001101;
    assign weights1[13][260] = 16'b0000000000010101;
    assign weights1[13][261] = 16'b0000000000001110;
    assign weights1[13][262] = 16'b1111111111110110;
    assign weights1[13][263] = 16'b0000000000000101;
    assign weights1[13][264] = 16'b0000000000000100;
    assign weights1[13][265] = 16'b0000000000001101;
    assign weights1[13][266] = 16'b1111111111111111;
    assign weights1[13][267] = 16'b0000000000000100;
    assign weights1[13][268] = 16'b1111111111111101;
    assign weights1[13][269] = 16'b0000000000000011;
    assign weights1[13][270] = 16'b1111111111111101;
    assign weights1[13][271] = 16'b0000000000000000;
    assign weights1[13][272] = 16'b0000000000001000;
    assign weights1[13][273] = 16'b0000000000010101;
    assign weights1[13][274] = 16'b0000000000010011;
    assign weights1[13][275] = 16'b0000000000001100;
    assign weights1[13][276] = 16'b0000000000000001;
    assign weights1[13][277] = 16'b0000000000001010;
    assign weights1[13][278] = 16'b0000000000000010;
    assign weights1[13][279] = 16'b0000000000000111;
    assign weights1[13][280] = 16'b1111111111101111;
    assign weights1[13][281] = 16'b1111111111100111;
    assign weights1[13][282] = 16'b1111111111011111;
    assign weights1[13][283] = 16'b1111111111110000;
    assign weights1[13][284] = 16'b0000000000000110;
    assign weights1[13][285] = 16'b1111111111110100;
    assign weights1[13][286] = 16'b1111111111111010;
    assign weights1[13][287] = 16'b0000000000000111;
    assign weights1[13][288] = 16'b0000000000000100;
    assign weights1[13][289] = 16'b1111111111101000;
    assign weights1[13][290] = 16'b0000000000001100;
    assign weights1[13][291] = 16'b1111111111110011;
    assign weights1[13][292] = 16'b1111111111100111;
    assign weights1[13][293] = 16'b1111111111111110;
    assign weights1[13][294] = 16'b1111111111110010;
    assign weights1[13][295] = 16'b1111111111111010;
    assign weights1[13][296] = 16'b1111111111111000;
    assign weights1[13][297] = 16'b1111111111111110;
    assign weights1[13][298] = 16'b1111111111111101;
    assign weights1[13][299] = 16'b1111111111101000;
    assign weights1[13][300] = 16'b1111111111111101;
    assign weights1[13][301] = 16'b1111111111111001;
    assign weights1[13][302] = 16'b1111111111101011;
    assign weights1[13][303] = 16'b0000000000000110;
    assign weights1[13][304] = 16'b1111111111111000;
    assign weights1[13][305] = 16'b0000000000001101;
    assign weights1[13][306] = 16'b0000000000010101;
    assign weights1[13][307] = 16'b0000000000001111;
    assign weights1[13][308] = 16'b1111111111100110;
    assign weights1[13][309] = 16'b1111111111010101;
    assign weights1[13][310] = 16'b1111111111001010;
    assign weights1[13][311] = 16'b1111111111011011;
    assign weights1[13][312] = 16'b1111111111100101;
    assign weights1[13][313] = 16'b1111111111110111;
    assign weights1[13][314] = 16'b1111111111110100;
    assign weights1[13][315] = 16'b1111111111110011;
    assign weights1[13][316] = 16'b1111111111111100;
    assign weights1[13][317] = 16'b1111111111110000;
    assign weights1[13][318] = 16'b1111111111101111;
    assign weights1[13][319] = 16'b0000000000011011;
    assign weights1[13][320] = 16'b0000000000010010;
    assign weights1[13][321] = 16'b0000000000001100;
    assign weights1[13][322] = 16'b0000000000000011;
    assign weights1[13][323] = 16'b0000000000001001;
    assign weights1[13][324] = 16'b1111111111111100;
    assign weights1[13][325] = 16'b1111111111111111;
    assign weights1[13][326] = 16'b1111111111111001;
    assign weights1[13][327] = 16'b0000000000000110;
    assign weights1[13][328] = 16'b1111111111011001;
    assign weights1[13][329] = 16'b1111111111100110;
    assign weights1[13][330] = 16'b0000000000000000;
    assign weights1[13][331] = 16'b1111111111110101;
    assign weights1[13][332] = 16'b0000000000000100;
    assign weights1[13][333] = 16'b0000000000000110;
    assign weights1[13][334] = 16'b1111111111111110;
    assign weights1[13][335] = 16'b0000000000000111;
    assign weights1[13][336] = 16'b1111111111011110;
    assign weights1[13][337] = 16'b1111111111000111;
    assign weights1[13][338] = 16'b1111111110101001;
    assign weights1[13][339] = 16'b1111111110110101;
    assign weights1[13][340] = 16'b1111111110111001;
    assign weights1[13][341] = 16'b1111111111100111;
    assign weights1[13][342] = 16'b1111111111011111;
    assign weights1[13][343] = 16'b0000000000011110;
    assign weights1[13][344] = 16'b1111111111110010;
    assign weights1[13][345] = 16'b0000000000010000;
    assign weights1[13][346] = 16'b0000000000011001;
    assign weights1[13][347] = 16'b0000000000001101;
    assign weights1[13][348] = 16'b0000000000000001;
    assign weights1[13][349] = 16'b0000000000010101;
    assign weights1[13][350] = 16'b0000000000010101;
    assign weights1[13][351] = 16'b0000000000010101;
    assign weights1[13][352] = 16'b0000000000001111;
    assign weights1[13][353] = 16'b0000000000000101;
    assign weights1[13][354] = 16'b1111111111111001;
    assign weights1[13][355] = 16'b0000000000000001;
    assign weights1[13][356] = 16'b0000000000001000;
    assign weights1[13][357] = 16'b1111111111110101;
    assign weights1[13][358] = 16'b1111111111100111;
    assign weights1[13][359] = 16'b1111111111101010;
    assign weights1[13][360] = 16'b0000000000001001;
    assign weights1[13][361] = 16'b1111111111111101;
    assign weights1[13][362] = 16'b0000000000000111;
    assign weights1[13][363] = 16'b0000000000000110;
    assign weights1[13][364] = 16'b1111111111011111;
    assign weights1[13][365] = 16'b1111111111001001;
    assign weights1[13][366] = 16'b1111111110100010;
    assign weights1[13][367] = 16'b1111111110011101;
    assign weights1[13][368] = 16'b1111111101111101;
    assign weights1[13][369] = 16'b1111111110000111;
    assign weights1[13][370] = 16'b1111111110100110;
    assign weights1[13][371] = 16'b1111111111110001;
    assign weights1[13][372] = 16'b0000000000010101;
    assign weights1[13][373] = 16'b0000000000011011;
    assign weights1[13][374] = 16'b0000000000001010;
    assign weights1[13][375] = 16'b0000000000010100;
    assign weights1[13][376] = 16'b0000000000000011;
    assign weights1[13][377] = 16'b0000000000011101;
    assign weights1[13][378] = 16'b0000000000011001;
    assign weights1[13][379] = 16'b0000000000001011;
    assign weights1[13][380] = 16'b0000000000001101;
    assign weights1[13][381] = 16'b0000000000000010;
    assign weights1[13][382] = 16'b0000000000000111;
    assign weights1[13][383] = 16'b0000000000000000;
    assign weights1[13][384] = 16'b1111111111110101;
    assign weights1[13][385] = 16'b0000000000001000;
    assign weights1[13][386] = 16'b1111111111110100;
    assign weights1[13][387] = 16'b1111111111101111;
    assign weights1[13][388] = 16'b1111111111100110;
    assign weights1[13][389] = 16'b1111111111110111;
    assign weights1[13][390] = 16'b0000000000010001;
    assign weights1[13][391] = 16'b0000000000010111;
    assign weights1[13][392] = 16'b1111111111101110;
    assign weights1[13][393] = 16'b1111111111011010;
    assign weights1[13][394] = 16'b1111111110101100;
    assign weights1[13][395] = 16'b1111111110011011;
    assign weights1[13][396] = 16'b1111111101100011;
    assign weights1[13][397] = 16'b1111111101000110;
    assign weights1[13][398] = 16'b1111111100101010;
    assign weights1[13][399] = 16'b1111111101011011;
    assign weights1[13][400] = 16'b1111111110100010;
    assign weights1[13][401] = 16'b1111111111110100;
    assign weights1[13][402] = 16'b0000000000001001;
    assign weights1[13][403] = 16'b0000000000010110;
    assign weights1[13][404] = 16'b0000000000101111;
    assign weights1[13][405] = 16'b0000000000100001;
    assign weights1[13][406] = 16'b0000000000010111;
    assign weights1[13][407] = 16'b0000000000000011;
    assign weights1[13][408] = 16'b0000000000010110;
    assign weights1[13][409] = 16'b1111111111110111;
    assign weights1[13][410] = 16'b0000000000000011;
    assign weights1[13][411] = 16'b1111111111111111;
    assign weights1[13][412] = 16'b1111111111110001;
    assign weights1[13][413] = 16'b1111111111111100;
    assign weights1[13][414] = 16'b0000000000000010;
    assign weights1[13][415] = 16'b1111111111111011;
    assign weights1[13][416] = 16'b1111111111100110;
    assign weights1[13][417] = 16'b1111111111111011;
    assign weights1[13][418] = 16'b1111111111111101;
    assign weights1[13][419] = 16'b0000000000001010;
    assign weights1[13][420] = 16'b0000000000000101;
    assign weights1[13][421] = 16'b1111111111110111;
    assign weights1[13][422] = 16'b1111111111011101;
    assign weights1[13][423] = 16'b1111111111010100;
    assign weights1[13][424] = 16'b1111111111001010;
    assign weights1[13][425] = 16'b1111111110001010;
    assign weights1[13][426] = 16'b1111111100111110;
    assign weights1[13][427] = 16'b1111111011110000;
    assign weights1[13][428] = 16'b1111111011101000;
    assign weights1[13][429] = 16'b1111111101000100;
    assign weights1[13][430] = 16'b1111111110111010;
    assign weights1[13][431] = 16'b1111111111111100;
    assign weights1[13][432] = 16'b0000000000100010;
    assign weights1[13][433] = 16'b0000000000011100;
    assign weights1[13][434] = 16'b0000000000011010;
    assign weights1[13][435] = 16'b0000000000011011;
    assign weights1[13][436] = 16'b0000000000000111;
    assign weights1[13][437] = 16'b0000000000000100;
    assign weights1[13][438] = 16'b1111111111110111;
    assign weights1[13][439] = 16'b0000000000000111;
    assign weights1[13][440] = 16'b1111111111111111;
    assign weights1[13][441] = 16'b0000000000000101;
    assign weights1[13][442] = 16'b0000000000000000;
    assign weights1[13][443] = 16'b0000000000001010;
    assign weights1[13][444] = 16'b1111111111110000;
    assign weights1[13][445] = 16'b1111111111111010;
    assign weights1[13][446] = 16'b1111111111101001;
    assign weights1[13][447] = 16'b0000000000000001;
    assign weights1[13][448] = 16'b0000000000010110;
    assign weights1[13][449] = 16'b0000000000010100;
    assign weights1[13][450] = 16'b0000000000010010;
    assign weights1[13][451] = 16'b0000000000101110;
    assign weights1[13][452] = 16'b0000000000001011;
    assign weights1[13][453] = 16'b0000000000001100;
    assign weights1[13][454] = 16'b1111111111110000;
    assign weights1[13][455] = 16'b1111111110100000;
    assign weights1[13][456] = 16'b1111111100011011;
    assign weights1[13][457] = 16'b1111111010110000;
    assign weights1[13][458] = 16'b1111111011010000;
    assign weights1[13][459] = 16'b1111111100100010;
    assign weights1[13][460] = 16'b1111111101111110;
    assign weights1[13][461] = 16'b1111111111010111;
    assign weights1[13][462] = 16'b1111111111111000;
    assign weights1[13][463] = 16'b1111111111111011;
    assign weights1[13][464] = 16'b1111111111111110;
    assign weights1[13][465] = 16'b1111111111111001;
    assign weights1[13][466] = 16'b0000000000000100;
    assign weights1[13][467] = 16'b0000000000010000;
    assign weights1[13][468] = 16'b1111111111111001;
    assign weights1[13][469] = 16'b0000000000001010;
    assign weights1[13][470] = 16'b0000000000000010;
    assign weights1[13][471] = 16'b0000000000000010;
    assign weights1[13][472] = 16'b1111111111111000;
    assign weights1[13][473] = 16'b1111111111110100;
    assign weights1[13][474] = 16'b1111111111110101;
    assign weights1[13][475] = 16'b1111111111111001;
    assign weights1[13][476] = 16'b0000000000011100;
    assign weights1[13][477] = 16'b0000000000011001;
    assign weights1[13][478] = 16'b0000000000100110;
    assign weights1[13][479] = 16'b0000000000110001;
    assign weights1[13][480] = 16'b0000000000010111;
    assign weights1[13][481] = 16'b0000000000101110;
    assign weights1[13][482] = 16'b0000000000110000;
    assign weights1[13][483] = 16'b0000000000101101;
    assign weights1[13][484] = 16'b0000000000011111;
    assign weights1[13][485] = 16'b1111111110111011;
    assign weights1[13][486] = 16'b1111111101100011;
    assign weights1[13][487] = 16'b1111111101000111;
    assign weights1[13][488] = 16'b1111111100110100;
    assign weights1[13][489] = 16'b1111111101110001;
    assign weights1[13][490] = 16'b1111111110011111;
    assign weights1[13][491] = 16'b1111111111010010;
    assign weights1[13][492] = 16'b1111111111100000;
    assign weights1[13][493] = 16'b1111111111100101;
    assign weights1[13][494] = 16'b1111111111110010;
    assign weights1[13][495] = 16'b1111111111110001;
    assign weights1[13][496] = 16'b1111111111111011;
    assign weights1[13][497] = 16'b1111111111111001;
    assign weights1[13][498] = 16'b1111111111110101;
    assign weights1[13][499] = 16'b0000000000000011;
    assign weights1[13][500] = 16'b0000000000001000;
    assign weights1[13][501] = 16'b0000000000001000;
    assign weights1[13][502] = 16'b1111111111111101;
    assign weights1[13][503] = 16'b1111111111111011;
    assign weights1[13][504] = 16'b0000000000011010;
    assign weights1[13][505] = 16'b1111111111111011;
    assign weights1[13][506] = 16'b0000000000100010;
    assign weights1[13][507] = 16'b0000000000100010;
    assign weights1[13][508] = 16'b0000000000101001;
    assign weights1[13][509] = 16'b0000000001011011;
    assign weights1[13][510] = 16'b0000000001101010;
    assign weights1[13][511] = 16'b0000000001001111;
    assign weights1[13][512] = 16'b0000000001100100;
    assign weights1[13][513] = 16'b0000000000111000;
    assign weights1[13][514] = 16'b0000000000000100;
    assign weights1[13][515] = 16'b1111111111010011;
    assign weights1[13][516] = 16'b1111111110101001;
    assign weights1[13][517] = 16'b1111111111000110;
    assign weights1[13][518] = 16'b1111111111000110;
    assign weights1[13][519] = 16'b1111111111011010;
    assign weights1[13][520] = 16'b1111111111100010;
    assign weights1[13][521] = 16'b1111111111101100;
    assign weights1[13][522] = 16'b1111111111110011;
    assign weights1[13][523] = 16'b1111111111111101;
    assign weights1[13][524] = 16'b1111111111110011;
    assign weights1[13][525] = 16'b0000000000001100;
    assign weights1[13][526] = 16'b0000000000010001;
    assign weights1[13][527] = 16'b1111111111111110;
    assign weights1[13][528] = 16'b1111111111101101;
    assign weights1[13][529] = 16'b0000000000001111;
    assign weights1[13][530] = 16'b0000000000000101;
    assign weights1[13][531] = 16'b0000000000000000;
    assign weights1[13][532] = 16'b1111111111111010;
    assign weights1[13][533] = 16'b1111111111111101;
    assign weights1[13][534] = 16'b0000000000001111;
    assign weights1[13][535] = 16'b0000000000100000;
    assign weights1[13][536] = 16'b0000000000110100;
    assign weights1[13][537] = 16'b0000000000111011;
    assign weights1[13][538] = 16'b0000000001000010;
    assign weights1[13][539] = 16'b0000000001001010;
    assign weights1[13][540] = 16'b0000000001010110;
    assign weights1[13][541] = 16'b0000000001101011;
    assign weights1[13][542] = 16'b0000000001000111;
    assign weights1[13][543] = 16'b0000000000101011;
    assign weights1[13][544] = 16'b0000000000010000;
    assign weights1[13][545] = 16'b1111111111110001;
    assign weights1[13][546] = 16'b1111111111100011;
    assign weights1[13][547] = 16'b1111111111110000;
    assign weights1[13][548] = 16'b1111111111100110;
    assign weights1[13][549] = 16'b1111111111011111;
    assign weights1[13][550] = 16'b0000000000000100;
    assign weights1[13][551] = 16'b1111111111100011;
    assign weights1[13][552] = 16'b1111111111111110;
    assign weights1[13][553] = 16'b0000000000000000;
    assign weights1[13][554] = 16'b0000000000000111;
    assign weights1[13][555] = 16'b1111111111111000;
    assign weights1[13][556] = 16'b0000000000000010;
    assign weights1[13][557] = 16'b1111111111111100;
    assign weights1[13][558] = 16'b0000000000000000;
    assign weights1[13][559] = 16'b1111111111110111;
    assign weights1[13][560] = 16'b1111111111110011;
    assign weights1[13][561] = 16'b1111111111011110;
    assign weights1[13][562] = 16'b1111111111111111;
    assign weights1[13][563] = 16'b1111111111111001;
    assign weights1[13][564] = 16'b0000000000100111;
    assign weights1[13][565] = 16'b0000000000001100;
    assign weights1[13][566] = 16'b0000000000010010;
    assign weights1[13][567] = 16'b0000000000001101;
    assign weights1[13][568] = 16'b0000000000001110;
    assign weights1[13][569] = 16'b0000000000010000;
    assign weights1[13][570] = 16'b0000000000100010;
    assign weights1[13][571] = 16'b0000000000011100;
    assign weights1[13][572] = 16'b0000000000101011;
    assign weights1[13][573] = 16'b1111111111111011;
    assign weights1[13][574] = 16'b1111111111110111;
    assign weights1[13][575] = 16'b1111111111111100;
    assign weights1[13][576] = 16'b1111111111111101;
    assign weights1[13][577] = 16'b0000000000000100;
    assign weights1[13][578] = 16'b1111111111101100;
    assign weights1[13][579] = 16'b0000000000001001;
    assign weights1[13][580] = 16'b1111111111110010;
    assign weights1[13][581] = 16'b0000000000000111;
    assign weights1[13][582] = 16'b1111111111101110;
    assign weights1[13][583] = 16'b0000000000000000;
    assign weights1[13][584] = 16'b0000000000000100;
    assign weights1[13][585] = 16'b1111111111111100;
    assign weights1[13][586] = 16'b1111111111111100;
    assign weights1[13][587] = 16'b1111111111111110;
    assign weights1[13][588] = 16'b1111111111101101;
    assign weights1[13][589] = 16'b1111111111010111;
    assign weights1[13][590] = 16'b1111111111000111;
    assign weights1[13][591] = 16'b1111111111010110;
    assign weights1[13][592] = 16'b1111111111111101;
    assign weights1[13][593] = 16'b0000000000001110;
    assign weights1[13][594] = 16'b0000000000001010;
    assign weights1[13][595] = 16'b0000000000001011;
    assign weights1[13][596] = 16'b0000000000010100;
    assign weights1[13][597] = 16'b1111111111111000;
    assign weights1[13][598] = 16'b0000000000010010;
    assign weights1[13][599] = 16'b0000000000011010;
    assign weights1[13][600] = 16'b0000000000010110;
    assign weights1[13][601] = 16'b0000000000011100;
    assign weights1[13][602] = 16'b0000000000100010;
    assign weights1[13][603] = 16'b0000000000001110;
    assign weights1[13][604] = 16'b1111111111111011;
    assign weights1[13][605] = 16'b0000000000000011;
    assign weights1[13][606] = 16'b1111111111111000;
    assign weights1[13][607] = 16'b0000000000000011;
    assign weights1[13][608] = 16'b0000000000000000;
    assign weights1[13][609] = 16'b1111111111110100;
    assign weights1[13][610] = 16'b0000000000001011;
    assign weights1[13][611] = 16'b1111111111110111;
    assign weights1[13][612] = 16'b1111111111110100;
    assign weights1[13][613] = 16'b1111111111111001;
    assign weights1[13][614] = 16'b1111111111101110;
    assign weights1[13][615] = 16'b1111111111110010;
    assign weights1[13][616] = 16'b1111111111101100;
    assign weights1[13][617] = 16'b1111111111011000;
    assign weights1[13][618] = 16'b1111111111000011;
    assign weights1[13][619] = 16'b1111111110111011;
    assign weights1[13][620] = 16'b1111111111000111;
    assign weights1[13][621] = 16'b1111111111000110;
    assign weights1[13][622] = 16'b1111111111110100;
    assign weights1[13][623] = 16'b1111111111101110;
    assign weights1[13][624] = 16'b0000000000000000;
    assign weights1[13][625] = 16'b0000000000011010;
    assign weights1[13][626] = 16'b0000000000000111;
    assign weights1[13][627] = 16'b0000000000000110;
    assign weights1[13][628] = 16'b0000000000000100;
    assign weights1[13][629] = 16'b0000000000001010;
    assign weights1[13][630] = 16'b0000000000000000;
    assign weights1[13][631] = 16'b0000000000001001;
    assign weights1[13][632] = 16'b0000000000001010;
    assign weights1[13][633] = 16'b1111111111111001;
    assign weights1[13][634] = 16'b0000000000001110;
    assign weights1[13][635] = 16'b1111111111111000;
    assign weights1[13][636] = 16'b1111111111110111;
    assign weights1[13][637] = 16'b1111111111110111;
    assign weights1[13][638] = 16'b1111111111101110;
    assign weights1[13][639] = 16'b0000000000001101;
    assign weights1[13][640] = 16'b1111111111110110;
    assign weights1[13][641] = 16'b1111111111111111;
    assign weights1[13][642] = 16'b1111111111101111;
    assign weights1[13][643] = 16'b1111111111111000;
    assign weights1[13][644] = 16'b1111111111110110;
    assign weights1[13][645] = 16'b1111111111100110;
    assign weights1[13][646] = 16'b1111111111011001;
    assign weights1[13][647] = 16'b1111111111001111;
    assign weights1[13][648] = 16'b1111111111001011;
    assign weights1[13][649] = 16'b1111111111100101;
    assign weights1[13][650] = 16'b1111111111101110;
    assign weights1[13][651] = 16'b1111111111111011;
    assign weights1[13][652] = 16'b1111111111111001;
    assign weights1[13][653] = 16'b1111111111111100;
    assign weights1[13][654] = 16'b0000000000110110;
    assign weights1[13][655] = 16'b0000000000011000;
    assign weights1[13][656] = 16'b0000000000001100;
    assign weights1[13][657] = 16'b0000000000001111;
    assign weights1[13][658] = 16'b0000000000001111;
    assign weights1[13][659] = 16'b0000000000000111;
    assign weights1[13][660] = 16'b1111111111110111;
    assign weights1[13][661] = 16'b0000000000000011;
    assign weights1[13][662] = 16'b0000000000001111;
    assign weights1[13][663] = 16'b0000000000000111;
    assign weights1[13][664] = 16'b0000000000010000;
    assign weights1[13][665] = 16'b0000000000000110;
    assign weights1[13][666] = 16'b1111111111111001;
    assign weights1[13][667] = 16'b1111111111101101;
    assign weights1[13][668] = 16'b1111111111110110;
    assign weights1[13][669] = 16'b1111111111110110;
    assign weights1[13][670] = 16'b1111111111110100;
    assign weights1[13][671] = 16'b1111111111110110;
    assign weights1[13][672] = 16'b1111111111111010;
    assign weights1[13][673] = 16'b1111111111110011;
    assign weights1[13][674] = 16'b1111111111101101;
    assign weights1[13][675] = 16'b1111111111011011;
    assign weights1[13][676] = 16'b1111111111011110;
    assign weights1[13][677] = 16'b1111111111010110;
    assign weights1[13][678] = 16'b1111111111011010;
    assign weights1[13][679] = 16'b1111111111111100;
    assign weights1[13][680] = 16'b0000000000000000;
    assign weights1[13][681] = 16'b1111111111111110;
    assign weights1[13][682] = 16'b0000000000000001;
    assign weights1[13][683] = 16'b1111111111111110;
    assign weights1[13][684] = 16'b0000000000010000;
    assign weights1[13][685] = 16'b1111111111111000;
    assign weights1[13][686] = 16'b0000000000000101;
    assign weights1[13][687] = 16'b0000000000000101;
    assign weights1[13][688] = 16'b1111111111110101;
    assign weights1[13][689] = 16'b0000000000000010;
    assign weights1[13][690] = 16'b0000000000000011;
    assign weights1[13][691] = 16'b1111111111101100;
    assign weights1[13][692] = 16'b1111111111110011;
    assign weights1[13][693] = 16'b0000000000000110;
    assign weights1[13][694] = 16'b1111111111011111;
    assign weights1[13][695] = 16'b1111111111101001;
    assign weights1[13][696] = 16'b1111111111110001;
    assign weights1[13][697] = 16'b1111111111110011;
    assign weights1[13][698] = 16'b1111111111111001;
    assign weights1[13][699] = 16'b1111111111111101;
    assign weights1[13][700] = 16'b1111111111111111;
    assign weights1[13][701] = 16'b1111111111111101;
    assign weights1[13][702] = 16'b1111111111111000;
    assign weights1[13][703] = 16'b1111111111111011;
    assign weights1[13][704] = 16'b1111111111101101;
    assign weights1[13][705] = 16'b1111111111011111;
    assign weights1[13][706] = 16'b1111111111100110;
    assign weights1[13][707] = 16'b1111111111110111;
    assign weights1[13][708] = 16'b1111111111111011;
    assign weights1[13][709] = 16'b1111111111100000;
    assign weights1[13][710] = 16'b1111111111111111;
    assign weights1[13][711] = 16'b1111111111101010;
    assign weights1[13][712] = 16'b1111111111110011;
    assign weights1[13][713] = 16'b0000000000001101;
    assign weights1[13][714] = 16'b0000000000010100;
    assign weights1[13][715] = 16'b0000000000000110;
    assign weights1[13][716] = 16'b0000000000000110;
    assign weights1[13][717] = 16'b0000000000001110;
    assign weights1[13][718] = 16'b0000000000000010;
    assign weights1[13][719] = 16'b1111111111111001;
    assign weights1[13][720] = 16'b1111111111110110;
    assign weights1[13][721] = 16'b1111111111101000;
    assign weights1[13][722] = 16'b1111111111011011;
    assign weights1[13][723] = 16'b1111111111101011;
    assign weights1[13][724] = 16'b1111111111110101;
    assign weights1[13][725] = 16'b1111111111110101;
    assign weights1[13][726] = 16'b1111111111111010;
    assign weights1[13][727] = 16'b0000000000000000;
    assign weights1[13][728] = 16'b1111111111111110;
    assign weights1[13][729] = 16'b1111111111111100;
    assign weights1[13][730] = 16'b0000000000000001;
    assign weights1[13][731] = 16'b0000000000000000;
    assign weights1[13][732] = 16'b1111111111111010;
    assign weights1[13][733] = 16'b1111111111110111;
    assign weights1[13][734] = 16'b1111111111101011;
    assign weights1[13][735] = 16'b1111111111011001;
    assign weights1[13][736] = 16'b1111111111100011;
    assign weights1[13][737] = 16'b1111111111100110;
    assign weights1[13][738] = 16'b1111111111110100;
    assign weights1[13][739] = 16'b1111111111100110;
    assign weights1[13][740] = 16'b1111111111111000;
    assign weights1[13][741] = 16'b1111111111111000;
    assign weights1[13][742] = 16'b1111111111100111;
    assign weights1[13][743] = 16'b1111111111110110;
    assign weights1[13][744] = 16'b0000000000000010;
    assign weights1[13][745] = 16'b1111111111111110;
    assign weights1[13][746] = 16'b1111111111101111;
    assign weights1[13][747] = 16'b1111111111101100;
    assign weights1[13][748] = 16'b1111111111101111;
    assign weights1[13][749] = 16'b1111111111100000;
    assign weights1[13][750] = 16'b1111111111101001;
    assign weights1[13][751] = 16'b1111111111111000;
    assign weights1[13][752] = 16'b1111111111111000;
    assign weights1[13][753] = 16'b1111111111111001;
    assign weights1[13][754] = 16'b1111111111111110;
    assign weights1[13][755] = 16'b0000000000000000;
    assign weights1[13][756] = 16'b0000000000000001;
    assign weights1[13][757] = 16'b0000000000000000;
    assign weights1[13][758] = 16'b0000000000000010;
    assign weights1[13][759] = 16'b0000000000001001;
    assign weights1[13][760] = 16'b0000000000000110;
    assign weights1[13][761] = 16'b0000000000000100;
    assign weights1[13][762] = 16'b0000000000000110;
    assign weights1[13][763] = 16'b1111111111111010;
    assign weights1[13][764] = 16'b1111111111100111;
    assign weights1[13][765] = 16'b1111111111101001;
    assign weights1[13][766] = 16'b1111111111011011;
    assign weights1[13][767] = 16'b1111111111011000;
    assign weights1[13][768] = 16'b1111111111100111;
    assign weights1[13][769] = 16'b1111111111100000;
    assign weights1[13][770] = 16'b1111111111101001;
    assign weights1[13][771] = 16'b1111111111101110;
    assign weights1[13][772] = 16'b1111111111100111;
    assign weights1[13][773] = 16'b1111111111100001;
    assign weights1[13][774] = 16'b1111111111110010;
    assign weights1[13][775] = 16'b1111111111110110;
    assign weights1[13][776] = 16'b1111111111110011;
    assign weights1[13][777] = 16'b1111111111101110;
    assign weights1[13][778] = 16'b1111111111110010;
    assign weights1[13][779] = 16'b1111111111110110;
    assign weights1[13][780] = 16'b1111111111111011;
    assign weights1[13][781] = 16'b1111111111111100;
    assign weights1[13][782] = 16'b0000000000000000;
    assign weights1[13][783] = 16'b0000000000000000;
    assign weights1[14][0] = 16'b0000000000000000;
    assign weights1[14][1] = 16'b0000000000000000;
    assign weights1[14][2] = 16'b0000000000000000;
    assign weights1[14][3] = 16'b0000000000000000;
    assign weights1[14][4] = 16'b1111111111111011;
    assign weights1[14][5] = 16'b1111111111111001;
    assign weights1[14][6] = 16'b1111111111111010;
    assign weights1[14][7] = 16'b1111111111111010;
    assign weights1[14][8] = 16'b1111111111110011;
    assign weights1[14][9] = 16'b1111111111101010;
    assign weights1[14][10] = 16'b1111111111110001;
    assign weights1[14][11] = 16'b1111111111110100;
    assign weights1[14][12] = 16'b1111111111110110;
    assign weights1[14][13] = 16'b1111111111111101;
    assign weights1[14][14] = 16'b1111111111110010;
    assign weights1[14][15] = 16'b1111111111111011;
    assign weights1[14][16] = 16'b0000000000001111;
    assign weights1[14][17] = 16'b0000000000000011;
    assign weights1[14][18] = 16'b1111111111111111;
    assign weights1[14][19] = 16'b1111111111111001;
    assign weights1[14][20] = 16'b1111111111110010;
    assign weights1[14][21] = 16'b1111111111111110;
    assign weights1[14][22] = 16'b0000000000000011;
    assign weights1[14][23] = 16'b0000000000000001;
    assign weights1[14][24] = 16'b1111111111111101;
    assign weights1[14][25] = 16'b1111111111111101;
    assign weights1[14][26] = 16'b1111111111111100;
    assign weights1[14][27] = 16'b1111111111111101;
    assign weights1[14][28] = 16'b0000000000000000;
    assign weights1[14][29] = 16'b0000000000000000;
    assign weights1[14][30] = 16'b1111111111111011;
    assign weights1[14][31] = 16'b1111111111111000;
    assign weights1[14][32] = 16'b1111111111111111;
    assign weights1[14][33] = 16'b1111111111110110;
    assign weights1[14][34] = 16'b1111111111110110;
    assign weights1[14][35] = 16'b1111111111110110;
    assign weights1[14][36] = 16'b1111111111111111;
    assign weights1[14][37] = 16'b1111111111101110;
    assign weights1[14][38] = 16'b1111111111110101;
    assign weights1[14][39] = 16'b1111111111110001;
    assign weights1[14][40] = 16'b1111111111110101;
    assign weights1[14][41] = 16'b1111111111111000;
    assign weights1[14][42] = 16'b0000000000000000;
    assign weights1[14][43] = 16'b1111111111111110;
    assign weights1[14][44] = 16'b1111111111111111;
    assign weights1[14][45] = 16'b1111111111110011;
    assign weights1[14][46] = 16'b0000000000000101;
    assign weights1[14][47] = 16'b1111111111111010;
    assign weights1[14][48] = 16'b1111111111111101;
    assign weights1[14][49] = 16'b1111111111111010;
    assign weights1[14][50] = 16'b0000000000000101;
    assign weights1[14][51] = 16'b1111111111110111;
    assign weights1[14][52] = 16'b1111111111110110;
    assign weights1[14][53] = 16'b1111111111111110;
    assign weights1[14][54] = 16'b1111111111111110;
    assign weights1[14][55] = 16'b1111111111111111;
    assign weights1[14][56] = 16'b1111111111111110;
    assign weights1[14][57] = 16'b1111111111111101;
    assign weights1[14][58] = 16'b1111111111110111;
    assign weights1[14][59] = 16'b1111111111111010;
    assign weights1[14][60] = 16'b1111111111110011;
    assign weights1[14][61] = 16'b1111111111111010;
    assign weights1[14][62] = 16'b1111111111111010;
    assign weights1[14][63] = 16'b1111111111111001;
    assign weights1[14][64] = 16'b1111111111111111;
    assign weights1[14][65] = 16'b0000000000000001;
    assign weights1[14][66] = 16'b1111111111110111;
    assign weights1[14][67] = 16'b1111111111111101;
    assign weights1[14][68] = 16'b1111111111111010;
    assign weights1[14][69] = 16'b0000000000000011;
    assign weights1[14][70] = 16'b1111111111111101;
    assign weights1[14][71] = 16'b0000000000001001;
    assign weights1[14][72] = 16'b1111111111111001;
    assign weights1[14][73] = 16'b1111111111111010;
    assign weights1[14][74] = 16'b1111111111110010;
    assign weights1[14][75] = 16'b1111111111111101;
    assign weights1[14][76] = 16'b0000000000000111;
    assign weights1[14][77] = 16'b1111111111111100;
    assign weights1[14][78] = 16'b1111111111110110;
    assign weights1[14][79] = 16'b0000000000000011;
    assign weights1[14][80] = 16'b1111111111111001;
    assign weights1[14][81] = 16'b0000000000001000;
    assign weights1[14][82] = 16'b1111111111111111;
    assign weights1[14][83] = 16'b1111111111111100;
    assign weights1[14][84] = 16'b1111111111111111;
    assign weights1[14][85] = 16'b1111111111111101;
    assign weights1[14][86] = 16'b0000000000000001;
    assign weights1[14][87] = 16'b0000000000000101;
    assign weights1[14][88] = 16'b1111111111111001;
    assign weights1[14][89] = 16'b1111111111111111;
    assign weights1[14][90] = 16'b0000000000001111;
    assign weights1[14][91] = 16'b1111111111111111;
    assign weights1[14][92] = 16'b1111111111111111;
    assign weights1[14][93] = 16'b0000000000000001;
    assign weights1[14][94] = 16'b1111111111111011;
    assign weights1[14][95] = 16'b1111111111111110;
    assign weights1[14][96] = 16'b1111111111110010;
    assign weights1[14][97] = 16'b1111111111110110;
    assign weights1[14][98] = 16'b1111111111110100;
    assign weights1[14][99] = 16'b0000000000000000;
    assign weights1[14][100] = 16'b1111111111101011;
    assign weights1[14][101] = 16'b0000000000010010;
    assign weights1[14][102] = 16'b0000000000010100;
    assign weights1[14][103] = 16'b0000000000000100;
    assign weights1[14][104] = 16'b1111111111111001;
    assign weights1[14][105] = 16'b1111111111101100;
    assign weights1[14][106] = 16'b1111111111111000;
    assign weights1[14][107] = 16'b1111111111101111;
    assign weights1[14][108] = 16'b1111111111111101;
    assign weights1[14][109] = 16'b1111111111110101;
    assign weights1[14][110] = 16'b0000000000000000;
    assign weights1[14][111] = 16'b0000000000000100;
    assign weights1[14][112] = 16'b1111111111111110;
    assign weights1[14][113] = 16'b1111111111111100;
    assign weights1[14][114] = 16'b1111111111111100;
    assign weights1[14][115] = 16'b0000000000000011;
    assign weights1[14][116] = 16'b1111111111111001;
    assign weights1[14][117] = 16'b0000000000001011;
    assign weights1[14][118] = 16'b0000000000000000;
    assign weights1[14][119] = 16'b1111111111110100;
    assign weights1[14][120] = 16'b1111111111111110;
    assign weights1[14][121] = 16'b1111111111111011;
    assign weights1[14][122] = 16'b1111111111111001;
    assign weights1[14][123] = 16'b1111111111111110;
    assign weights1[14][124] = 16'b0000000000000011;
    assign weights1[14][125] = 16'b0000000000001100;
    assign weights1[14][126] = 16'b1111111111110101;
    assign weights1[14][127] = 16'b0000000000001110;
    assign weights1[14][128] = 16'b0000000000010010;
    assign weights1[14][129] = 16'b1111111111101011;
    assign weights1[14][130] = 16'b1111111111110110;
    assign weights1[14][131] = 16'b0000000000000010;
    assign weights1[14][132] = 16'b0000000000000101;
    assign weights1[14][133] = 16'b0000000000001011;
    assign weights1[14][134] = 16'b0000000000000000;
    assign weights1[14][135] = 16'b1111111111111011;
    assign weights1[14][136] = 16'b0000000000001011;
    assign weights1[14][137] = 16'b1111111111111100;
    assign weights1[14][138] = 16'b1111111111111101;
    assign weights1[14][139] = 16'b0000000000000110;
    assign weights1[14][140] = 16'b0000000000000100;
    assign weights1[14][141] = 16'b1111111111111011;
    assign weights1[14][142] = 16'b0000000000000010;
    assign weights1[14][143] = 16'b1111111111111010;
    assign weights1[14][144] = 16'b1111111111111100;
    assign weights1[14][145] = 16'b0000000000001000;
    assign weights1[14][146] = 16'b0000000000000010;
    assign weights1[14][147] = 16'b1111111111111110;
    assign weights1[14][148] = 16'b0000000000001010;
    assign weights1[14][149] = 16'b0000000000000001;
    assign weights1[14][150] = 16'b1111111111111001;
    assign weights1[14][151] = 16'b1111111111111001;
    assign weights1[14][152] = 16'b0000000000001001;
    assign weights1[14][153] = 16'b0000000000000110;
    assign weights1[14][154] = 16'b1111111111110111;
    assign weights1[14][155] = 16'b1111111111110101;
    assign weights1[14][156] = 16'b0000000000000100;
    assign weights1[14][157] = 16'b1111111111111001;
    assign weights1[14][158] = 16'b0000000000001011;
    assign weights1[14][159] = 16'b1111111111111011;
    assign weights1[14][160] = 16'b1111111111111110;
    assign weights1[14][161] = 16'b1111111111111101;
    assign weights1[14][162] = 16'b1111111111110101;
    assign weights1[14][163] = 16'b1111111111111010;
    assign weights1[14][164] = 16'b0000000000000111;
    assign weights1[14][165] = 16'b0000000000000101;
    assign weights1[14][166] = 16'b0000000000000010;
    assign weights1[14][167] = 16'b0000000000000010;
    assign weights1[14][168] = 16'b0000000000000101;
    assign weights1[14][169] = 16'b1111111111111101;
    assign weights1[14][170] = 16'b1111111111110110;
    assign weights1[14][171] = 16'b0000000000001001;
    assign weights1[14][172] = 16'b1111111111111111;
    assign weights1[14][173] = 16'b1111111111101110;
    assign weights1[14][174] = 16'b0000000000000011;
    assign weights1[14][175] = 16'b0000000000000001;
    assign weights1[14][176] = 16'b1111111111111001;
    assign weights1[14][177] = 16'b0000000000001111;
    assign weights1[14][178] = 16'b1111111111110110;
    assign weights1[14][179] = 16'b1111111111111110;
    assign weights1[14][180] = 16'b1111111111110010;
    assign weights1[14][181] = 16'b1111111111101101;
    assign weights1[14][182] = 16'b0000000000000000;
    assign weights1[14][183] = 16'b0000000000000101;
    assign weights1[14][184] = 16'b1111111111111011;
    assign weights1[14][185] = 16'b0000000000000001;
    assign weights1[14][186] = 16'b0000000000010000;
    assign weights1[14][187] = 16'b1111111111110011;
    assign weights1[14][188] = 16'b0000000000000100;
    assign weights1[14][189] = 16'b1111111111110100;
    assign weights1[14][190] = 16'b1111111111111100;
    assign weights1[14][191] = 16'b0000000000001101;
    assign weights1[14][192] = 16'b0000000000000001;
    assign weights1[14][193] = 16'b1111111111111111;
    assign weights1[14][194] = 16'b0000000000000100;
    assign weights1[14][195] = 16'b0000000000001000;
    assign weights1[14][196] = 16'b0000000000000000;
    assign weights1[14][197] = 16'b1111111111111100;
    assign weights1[14][198] = 16'b0000000000000001;
    assign weights1[14][199] = 16'b1111111111110111;
    assign weights1[14][200] = 16'b0000000000000100;
    assign weights1[14][201] = 16'b1111111111111011;
    assign weights1[14][202] = 16'b0000000000001011;
    assign weights1[14][203] = 16'b0000000000001001;
    assign weights1[14][204] = 16'b1111111111111000;
    assign weights1[14][205] = 16'b1111111111110111;
    assign weights1[14][206] = 16'b0000000000000011;
    assign weights1[14][207] = 16'b1111111111110111;
    assign weights1[14][208] = 16'b1111111111111001;
    assign weights1[14][209] = 16'b1111111111111010;
    assign weights1[14][210] = 16'b0000000000000011;
    assign weights1[14][211] = 16'b1111111111110010;
    assign weights1[14][212] = 16'b1111111111111100;
    assign weights1[14][213] = 16'b1111111111111111;
    assign weights1[14][214] = 16'b0000000000000001;
    assign weights1[14][215] = 16'b1111111111101100;
    assign weights1[14][216] = 16'b0000000000001111;
    assign weights1[14][217] = 16'b1111111111101111;
    assign weights1[14][218] = 16'b0000000000001110;
    assign weights1[14][219] = 16'b0000000000001011;
    assign weights1[14][220] = 16'b1111111111110111;
    assign weights1[14][221] = 16'b0000000000001010;
    assign weights1[14][222] = 16'b0000000000000111;
    assign weights1[14][223] = 16'b1111111111111110;
    assign weights1[14][224] = 16'b0000000000001000;
    assign weights1[14][225] = 16'b0000000000000110;
    assign weights1[14][226] = 16'b0000000000001011;
    assign weights1[14][227] = 16'b0000000000001000;
    assign weights1[14][228] = 16'b1111111111110110;
    assign weights1[14][229] = 16'b0000000000010000;
    assign weights1[14][230] = 16'b0000000000000110;
    assign weights1[14][231] = 16'b0000000000000111;
    assign weights1[14][232] = 16'b1111111111110101;
    assign weights1[14][233] = 16'b1111111111111010;
    assign weights1[14][234] = 16'b1111111111110111;
    assign weights1[14][235] = 16'b0000000000000001;
    assign weights1[14][236] = 16'b0000000000001001;
    assign weights1[14][237] = 16'b0000000000001010;
    assign weights1[14][238] = 16'b0000000000000010;
    assign weights1[14][239] = 16'b0000000000001010;
    assign weights1[14][240] = 16'b1111111111101110;
    assign weights1[14][241] = 16'b0000000000001011;
    assign weights1[14][242] = 16'b0000000000000110;
    assign weights1[14][243] = 16'b1111111111111010;
    assign weights1[14][244] = 16'b0000000000001101;
    assign weights1[14][245] = 16'b0000000000000010;
    assign weights1[14][246] = 16'b0000000000000010;
    assign weights1[14][247] = 16'b0000000000000000;
    assign weights1[14][248] = 16'b0000000000001000;
    assign weights1[14][249] = 16'b1111111111111001;
    assign weights1[14][250] = 16'b1111111111111111;
    assign weights1[14][251] = 16'b1111111111101111;
    assign weights1[14][252] = 16'b0000000000001010;
    assign weights1[14][253] = 16'b0000000000000101;
    assign weights1[14][254] = 16'b0000000000000100;
    assign weights1[14][255] = 16'b1111111111111101;
    assign weights1[14][256] = 16'b1111111111110111;
    assign weights1[14][257] = 16'b0000000000000000;
    assign weights1[14][258] = 16'b1111111111111011;
    assign weights1[14][259] = 16'b0000000000001011;
    assign weights1[14][260] = 16'b0000000000001100;
    assign weights1[14][261] = 16'b0000000000011001;
    assign weights1[14][262] = 16'b0000000000000010;
    assign weights1[14][263] = 16'b1111111111101110;
    assign weights1[14][264] = 16'b1111111111111111;
    assign weights1[14][265] = 16'b0000000000000110;
    assign weights1[14][266] = 16'b1111111111111110;
    assign weights1[14][267] = 16'b0000000000000010;
    assign weights1[14][268] = 16'b1111111111110111;
    assign weights1[14][269] = 16'b1111111111111010;
    assign weights1[14][270] = 16'b1111111111111100;
    assign weights1[14][271] = 16'b1111111111110110;
    assign weights1[14][272] = 16'b1111111111110111;
    assign weights1[14][273] = 16'b1111111111101010;
    assign weights1[14][274] = 16'b0000000000000110;
    assign weights1[14][275] = 16'b1111111111111111;
    assign weights1[14][276] = 16'b1111111111111101;
    assign weights1[14][277] = 16'b0000000000001100;
    assign weights1[14][278] = 16'b0000000000000110;
    assign weights1[14][279] = 16'b1111111111111110;
    assign weights1[14][280] = 16'b0000000000010000;
    assign weights1[14][281] = 16'b0000000000000100;
    assign weights1[14][282] = 16'b0000000000001001;
    assign weights1[14][283] = 16'b0000000000000001;
    assign weights1[14][284] = 16'b1111111111111100;
    assign weights1[14][285] = 16'b0000000000000001;
    assign weights1[14][286] = 16'b1111111111110100;
    assign weights1[14][287] = 16'b1111111111111010;
    assign weights1[14][288] = 16'b0000000000000011;
    assign weights1[14][289] = 16'b0000000000000010;
    assign weights1[14][290] = 16'b1111111111101001;
    assign weights1[14][291] = 16'b0000000000000100;
    assign weights1[14][292] = 16'b0000000000001100;
    assign weights1[14][293] = 16'b1111111111111010;
    assign weights1[14][294] = 16'b0000000000001110;
    assign weights1[14][295] = 16'b0000000000000011;
    assign weights1[14][296] = 16'b1111111111101011;
    assign weights1[14][297] = 16'b0000000000001110;
    assign weights1[14][298] = 16'b1111111111110110;
    assign weights1[14][299] = 16'b1111111111111001;
    assign weights1[14][300] = 16'b0000000000001010;
    assign weights1[14][301] = 16'b0000000000001010;
    assign weights1[14][302] = 16'b1111111111111000;
    assign weights1[14][303] = 16'b0000000000000101;
    assign weights1[14][304] = 16'b1111111111111100;
    assign weights1[14][305] = 16'b1111111111111011;
    assign weights1[14][306] = 16'b0000000000000001;
    assign weights1[14][307] = 16'b0000000000000111;
    assign weights1[14][308] = 16'b0000000000001101;
    assign weights1[14][309] = 16'b0000000000001000;
    assign weights1[14][310] = 16'b0000000000010001;
    assign weights1[14][311] = 16'b0000000000001001;
    assign weights1[14][312] = 16'b0000000000000111;
    assign weights1[14][313] = 16'b0000000000001100;
    assign weights1[14][314] = 16'b0000000000010110;
    assign weights1[14][315] = 16'b1111111111110101;
    assign weights1[14][316] = 16'b0000000000001000;
    assign weights1[14][317] = 16'b0000000000001011;
    assign weights1[14][318] = 16'b0000000000000011;
    assign weights1[14][319] = 16'b0000000000000010;
    assign weights1[14][320] = 16'b0000000000000110;
    assign weights1[14][321] = 16'b1111111111101100;
    assign weights1[14][322] = 16'b0000000000000000;
    assign weights1[14][323] = 16'b0000000000001011;
    assign weights1[14][324] = 16'b0000000000000011;
    assign weights1[14][325] = 16'b0000000000000111;
    assign weights1[14][326] = 16'b1111111111111100;
    assign weights1[14][327] = 16'b1111111111111101;
    assign weights1[14][328] = 16'b1111111111111001;
    assign weights1[14][329] = 16'b0000000000000010;
    assign weights1[14][330] = 16'b0000000000001100;
    assign weights1[14][331] = 16'b0000000000000110;
    assign weights1[14][332] = 16'b0000000000000011;
    assign weights1[14][333] = 16'b1111111111111010;
    assign weights1[14][334] = 16'b1111111111110010;
    assign weights1[14][335] = 16'b0000000000000101;
    assign weights1[14][336] = 16'b0000000000000010;
    assign weights1[14][337] = 16'b0000000000000010;
    assign weights1[14][338] = 16'b1111111111111111;
    assign weights1[14][339] = 16'b0000000000001011;
    assign weights1[14][340] = 16'b0000000000010011;
    assign weights1[14][341] = 16'b1111111111111100;
    assign weights1[14][342] = 16'b1111111111111001;
    assign weights1[14][343] = 16'b0000000000001100;
    assign weights1[14][344] = 16'b0000000000000100;
    assign weights1[14][345] = 16'b0000000000000001;
    assign weights1[14][346] = 16'b1111111111110101;
    assign weights1[14][347] = 16'b0000000000000011;
    assign weights1[14][348] = 16'b0000000000000111;
    assign weights1[14][349] = 16'b1111111111111101;
    assign weights1[14][350] = 16'b1111111111111010;
    assign weights1[14][351] = 16'b1111111111111111;
    assign weights1[14][352] = 16'b0000000000000111;
    assign weights1[14][353] = 16'b1111111111101101;
    assign weights1[14][354] = 16'b1111111111111100;
    assign weights1[14][355] = 16'b0000000000000111;
    assign weights1[14][356] = 16'b0000000000000000;
    assign weights1[14][357] = 16'b0000000000000010;
    assign weights1[14][358] = 16'b1111111111101110;
    assign weights1[14][359] = 16'b1111111111110011;
    assign weights1[14][360] = 16'b1111111111111011;
    assign weights1[14][361] = 16'b1111111111111011;
    assign weights1[14][362] = 16'b1111111111111010;
    assign weights1[14][363] = 16'b1111111111111011;
    assign weights1[14][364] = 16'b0000000000000100;
    assign weights1[14][365] = 16'b1111111111110101;
    assign weights1[14][366] = 16'b0000000000000011;
    assign weights1[14][367] = 16'b0000000000000111;
    assign weights1[14][368] = 16'b0000000000000000;
    assign weights1[14][369] = 16'b1111111111111101;
    assign weights1[14][370] = 16'b1111111111111111;
    assign weights1[14][371] = 16'b0000000000001001;
    assign weights1[14][372] = 16'b0000000000000100;
    assign weights1[14][373] = 16'b0000000000001000;
    assign weights1[14][374] = 16'b1111111111111001;
    assign weights1[14][375] = 16'b0000000000010011;
    assign weights1[14][376] = 16'b1111111111110011;
    assign weights1[14][377] = 16'b1111111111111100;
    assign weights1[14][378] = 16'b1111111111111111;
    assign weights1[14][379] = 16'b0000000000000111;
    assign weights1[14][380] = 16'b1111111111111101;
    assign weights1[14][381] = 16'b0000000000000110;
    assign weights1[14][382] = 16'b0000000000000000;
    assign weights1[14][383] = 16'b1111111111110101;
    assign weights1[14][384] = 16'b1111111111111011;
    assign weights1[14][385] = 16'b0000000000010000;
    assign weights1[14][386] = 16'b0000000000001110;
    assign weights1[14][387] = 16'b1111111111110010;
    assign weights1[14][388] = 16'b0000000000000100;
    assign weights1[14][389] = 16'b0000000000000001;
    assign weights1[14][390] = 16'b0000000000001001;
    assign weights1[14][391] = 16'b1111111111110110;
    assign weights1[14][392] = 16'b0000000000000001;
    assign weights1[14][393] = 16'b0000000000000011;
    assign weights1[14][394] = 16'b0000000000001110;
    assign weights1[14][395] = 16'b1111111111110101;
    assign weights1[14][396] = 16'b0000000000001001;
    assign weights1[14][397] = 16'b0000000000000000;
    assign weights1[14][398] = 16'b0000000000000010;
    assign weights1[14][399] = 16'b1111111111111100;
    assign weights1[14][400] = 16'b1111111111111000;
    assign weights1[14][401] = 16'b1111111111111111;
    assign weights1[14][402] = 16'b0000000000001000;
    assign weights1[14][403] = 16'b1111111111111000;
    assign weights1[14][404] = 16'b1111111111111000;
    assign weights1[14][405] = 16'b1111111111110101;
    assign weights1[14][406] = 16'b1111111111111101;
    assign weights1[14][407] = 16'b1111111111110110;
    assign weights1[14][408] = 16'b1111111111110110;
    assign weights1[14][409] = 16'b0000000000001001;
    assign weights1[14][410] = 16'b1111111111111100;
    assign weights1[14][411] = 16'b0000000000000110;
    assign weights1[14][412] = 16'b1111111111111111;
    assign weights1[14][413] = 16'b1111111111111111;
    assign weights1[14][414] = 16'b0000000000000101;
    assign weights1[14][415] = 16'b0000000000000101;
    assign weights1[14][416] = 16'b1111111111101100;
    assign weights1[14][417] = 16'b0000000000010111;
    assign weights1[14][418] = 16'b1111111111101101;
    assign weights1[14][419] = 16'b1111111111110111;
    assign weights1[14][420] = 16'b1111111111111110;
    assign weights1[14][421] = 16'b0000000000000100;
    assign weights1[14][422] = 16'b1111111111111010;
    assign weights1[14][423] = 16'b1111111111111100;
    assign weights1[14][424] = 16'b0000000000000111;
    assign weights1[14][425] = 16'b1111111111111101;
    assign weights1[14][426] = 16'b1111111111111110;
    assign weights1[14][427] = 16'b1111111111111100;
    assign weights1[14][428] = 16'b0000000000001110;
    assign weights1[14][429] = 16'b0000000000001100;
    assign weights1[14][430] = 16'b0000000000001010;
    assign weights1[14][431] = 16'b1111111111111000;
    assign weights1[14][432] = 16'b1111111111111110;
    assign weights1[14][433] = 16'b0000000000000000;
    assign weights1[14][434] = 16'b0000000000001000;
    assign weights1[14][435] = 16'b0000000000000110;
    assign weights1[14][436] = 16'b0000000000000001;
    assign weights1[14][437] = 16'b0000000000000101;
    assign weights1[14][438] = 16'b1111111111111111;
    assign weights1[14][439] = 16'b0000000000000011;
    assign weights1[14][440] = 16'b0000000000001000;
    assign weights1[14][441] = 16'b0000000000000111;
    assign weights1[14][442] = 16'b1111111111111111;
    assign weights1[14][443] = 16'b0000000000000010;
    assign weights1[14][444] = 16'b1111111111111011;
    assign weights1[14][445] = 16'b0000000000000001;
    assign weights1[14][446] = 16'b0000000000000000;
    assign weights1[14][447] = 16'b1111111111111011;
    assign weights1[14][448] = 16'b1111111111110010;
    assign weights1[14][449] = 16'b1111111111110011;
    assign weights1[14][450] = 16'b1111111111110001;
    assign weights1[14][451] = 16'b1111111111101000;
    assign weights1[14][452] = 16'b1111111111110111;
    assign weights1[14][453] = 16'b1111111111101011;
    assign weights1[14][454] = 16'b1111111111101110;
    assign weights1[14][455] = 16'b0000000000001100;
    assign weights1[14][456] = 16'b0000000000010010;
    assign weights1[14][457] = 16'b0000000000000101;
    assign weights1[14][458] = 16'b0000000000000110;
    assign weights1[14][459] = 16'b1111111111110011;
    assign weights1[14][460] = 16'b1111111111110000;
    assign weights1[14][461] = 16'b1111111111111000;
    assign weights1[14][462] = 16'b1111111111111101;
    assign weights1[14][463] = 16'b0000000000000001;
    assign weights1[14][464] = 16'b0000000000000010;
    assign weights1[14][465] = 16'b1111111111111100;
    assign weights1[14][466] = 16'b1111111111110000;
    assign weights1[14][467] = 16'b0000000000000011;
    assign weights1[14][468] = 16'b0000000000001010;
    assign weights1[14][469] = 16'b0000000000001110;
    assign weights1[14][470] = 16'b0000000000011010;
    assign weights1[14][471] = 16'b0000000000010111;
    assign weights1[14][472] = 16'b0000000000000100;
    assign weights1[14][473] = 16'b1111111111110010;
    assign weights1[14][474] = 16'b1111111111111011;
    assign weights1[14][475] = 16'b1111111111111011;
    assign weights1[14][476] = 16'b1111111111101100;
    assign weights1[14][477] = 16'b1111111111101110;
    assign weights1[14][478] = 16'b1111111111100111;
    assign weights1[14][479] = 16'b1111111111101110;
    assign weights1[14][480] = 16'b1111111111110101;
    assign weights1[14][481] = 16'b1111111111101110;
    assign weights1[14][482] = 16'b0000000000010000;
    assign weights1[14][483] = 16'b0000000000010000;
    assign weights1[14][484] = 16'b0000000000011111;
    assign weights1[14][485] = 16'b0000000000000011;
    assign weights1[14][486] = 16'b1111111111110110;
    assign weights1[14][487] = 16'b1111111111100101;
    assign weights1[14][488] = 16'b1111111111101000;
    assign weights1[14][489] = 16'b1111111111111001;
    assign weights1[14][490] = 16'b0000000000001110;
    assign weights1[14][491] = 16'b0000000000000110;
    assign weights1[14][492] = 16'b0000000000001101;
    assign weights1[14][493] = 16'b1111111111110000;
    assign weights1[14][494] = 16'b1111111111111000;
    assign weights1[14][495] = 16'b1111111111111000;
    assign weights1[14][496] = 16'b1111111111111101;
    assign weights1[14][497] = 16'b1111111111111111;
    assign weights1[14][498] = 16'b0000000000100110;
    assign weights1[14][499] = 16'b0000000000010111;
    assign weights1[14][500] = 16'b0000000000010010;
    assign weights1[14][501] = 16'b0000000000000011;
    assign weights1[14][502] = 16'b1111111111111010;
    assign weights1[14][503] = 16'b1111111111111011;
    assign weights1[14][504] = 16'b1111111111101000;
    assign weights1[14][505] = 16'b1111111111011101;
    assign weights1[14][506] = 16'b1111111111010100;
    assign weights1[14][507] = 16'b1111111111110010;
    assign weights1[14][508] = 16'b1111111111111000;
    assign weights1[14][509] = 16'b0000000000000101;
    assign weights1[14][510] = 16'b0000000000100011;
    assign weights1[14][511] = 16'b0000000000110011;
    assign weights1[14][512] = 16'b0000000000101000;
    assign weights1[14][513] = 16'b1111111111111111;
    assign weights1[14][514] = 16'b1111111111101001;
    assign weights1[14][515] = 16'b1111111111101001;
    assign weights1[14][516] = 16'b1111111111001111;
    assign weights1[14][517] = 16'b0000000000000010;
    assign weights1[14][518] = 16'b0000000000011010;
    assign weights1[14][519] = 16'b0000000000101110;
    assign weights1[14][520] = 16'b1111111111110110;
    assign weights1[14][521] = 16'b1111111111110100;
    assign weights1[14][522] = 16'b1111111111101111;
    assign weights1[14][523] = 16'b1111111111100101;
    assign weights1[14][524] = 16'b0000000000001101;
    assign weights1[14][525] = 16'b0000000000001000;
    assign weights1[14][526] = 16'b0000000000011110;
    assign weights1[14][527] = 16'b0000000000010001;
    assign weights1[14][528] = 16'b0000000000010010;
    assign weights1[14][529] = 16'b0000000000010110;
    assign weights1[14][530] = 16'b0000000000001100;
    assign weights1[14][531] = 16'b0000000000000000;
    assign weights1[14][532] = 16'b1111111111100010;
    assign weights1[14][533] = 16'b1111111111011110;
    assign weights1[14][534] = 16'b1111111111110010;
    assign weights1[14][535] = 16'b1111111111101111;
    assign weights1[14][536] = 16'b0000000000000101;
    assign weights1[14][537] = 16'b0000000000011111;
    assign weights1[14][538] = 16'b0000000000101101;
    assign weights1[14][539] = 16'b0000000000100011;
    assign weights1[14][540] = 16'b0000000000010101;
    assign weights1[14][541] = 16'b1111111111101101;
    assign weights1[14][542] = 16'b1111111111011111;
    assign weights1[14][543] = 16'b1111111110111010;
    assign weights1[14][544] = 16'b1111111111010110;
    assign weights1[14][545] = 16'b0000000000010011;
    assign weights1[14][546] = 16'b0000000000100100;
    assign weights1[14][547] = 16'b0000000000100101;
    assign weights1[14][548] = 16'b1111111111110010;
    assign weights1[14][549] = 16'b1111111111010100;
    assign weights1[14][550] = 16'b1111111111100001;
    assign weights1[14][551] = 16'b1111111111100000;
    assign weights1[14][552] = 16'b1111111111111000;
    assign weights1[14][553] = 16'b1111111111110001;
    assign weights1[14][554] = 16'b0000000000011111;
    assign weights1[14][555] = 16'b0000000000100101;
    assign weights1[14][556] = 16'b0000000000010111;
    assign weights1[14][557] = 16'b0000000000011000;
    assign weights1[14][558] = 16'b0000000000001100;
    assign weights1[14][559] = 16'b0000000000000011;
    assign weights1[14][560] = 16'b1111111111101001;
    assign weights1[14][561] = 16'b1111111111110111;
    assign weights1[14][562] = 16'b0000000000000011;
    assign weights1[14][563] = 16'b0000000000010001;
    assign weights1[14][564] = 16'b0000000000111010;
    assign weights1[14][565] = 16'b0000000000101111;
    assign weights1[14][566] = 16'b0000000000101010;
    assign weights1[14][567] = 16'b0000000000000010;
    assign weights1[14][568] = 16'b1111111111111011;
    assign weights1[14][569] = 16'b1111111111010111;
    assign weights1[14][570] = 16'b1111111111000001;
    assign weights1[14][571] = 16'b1111111110110001;
    assign weights1[14][572] = 16'b1111111111101100;
    assign weights1[14][573] = 16'b0000000000010011;
    assign weights1[14][574] = 16'b0000000000110110;
    assign weights1[14][575] = 16'b0000000000101101;
    assign weights1[14][576] = 16'b0000000000000010;
    assign weights1[14][577] = 16'b1111111111010100;
    assign weights1[14][578] = 16'b1111111111001100;
    assign weights1[14][579] = 16'b1111111111011010;
    assign weights1[14][580] = 16'b1111111111011101;
    assign weights1[14][581] = 16'b1111111111110011;
    assign weights1[14][582] = 16'b0000000000100111;
    assign weights1[14][583] = 16'b0000000000100011;
    assign weights1[14][584] = 16'b0000000000110100;
    assign weights1[14][585] = 16'b0000000000010101;
    assign weights1[14][586] = 16'b0000000000000110;
    assign weights1[14][587] = 16'b0000000000000000;
    assign weights1[14][588] = 16'b0000000000001010;
    assign weights1[14][589] = 16'b0000000000010010;
    assign weights1[14][590] = 16'b0000000000011111;
    assign weights1[14][591] = 16'b0000000000100101;
    assign weights1[14][592] = 16'b0000000000101101;
    assign weights1[14][593] = 16'b0000000000110100;
    assign weights1[14][594] = 16'b0000000000101010;
    assign weights1[14][595] = 16'b1111111111110101;
    assign weights1[14][596] = 16'b1111111111011001;
    assign weights1[14][597] = 16'b1111111110011000;
    assign weights1[14][598] = 16'b1111111110001111;
    assign weights1[14][599] = 16'b1111111111000011;
    assign weights1[14][600] = 16'b0000000000000100;
    assign weights1[14][601] = 16'b0000000000101011;
    assign weights1[14][602] = 16'b0000000000111110;
    assign weights1[14][603] = 16'b0000000000100111;
    assign weights1[14][604] = 16'b0000000000000000;
    assign weights1[14][605] = 16'b1111111111010101;
    assign weights1[14][606] = 16'b1111111110011010;
    assign weights1[14][607] = 16'b1111111110111101;
    assign weights1[14][608] = 16'b1111111110111111;
    assign weights1[14][609] = 16'b1111111111111010;
    assign weights1[14][610] = 16'b0000000000001110;
    assign weights1[14][611] = 16'b0000000000101101;
    assign weights1[14][612] = 16'b0000000000101110;
    assign weights1[14][613] = 16'b0000000000011001;
    assign weights1[14][614] = 16'b0000000000001111;
    assign weights1[14][615] = 16'b0000000000001001;
    assign weights1[14][616] = 16'b0000000000010111;
    assign weights1[14][617] = 16'b0000000000011010;
    assign weights1[14][618] = 16'b0000000000101101;
    assign weights1[14][619] = 16'b0000000000101101;
    assign weights1[14][620] = 16'b0000000000101011;
    assign weights1[14][621] = 16'b0000000000011011;
    assign weights1[14][622] = 16'b1111111111111010;
    assign weights1[14][623] = 16'b1111111110110001;
    assign weights1[14][624] = 16'b1111111110000111;
    assign weights1[14][625] = 16'b1111111101110001;
    assign weights1[14][626] = 16'b1111111110000011;
    assign weights1[14][627] = 16'b1111111111010100;
    assign weights1[14][628] = 16'b0000000000100010;
    assign weights1[14][629] = 16'b0000000000101100;
    assign weights1[14][630] = 16'b0000000000100100;
    assign weights1[14][631] = 16'b0000000001000001;
    assign weights1[14][632] = 16'b1111111111110101;
    assign weights1[14][633] = 16'b1111111110111100;
    assign weights1[14][634] = 16'b1111111110100000;
    assign weights1[14][635] = 16'b1111111111000100;
    assign weights1[14][636] = 16'b1111111110111111;
    assign weights1[14][637] = 16'b1111111111001010;
    assign weights1[14][638] = 16'b1111111111110110;
    assign weights1[14][639] = 16'b0000000000010100;
    assign weights1[14][640] = 16'b0000000000100001;
    assign weights1[14][641] = 16'b0000000000011110;
    assign weights1[14][642] = 16'b0000000000010010;
    assign weights1[14][643] = 16'b0000000000001111;
    assign weights1[14][644] = 16'b0000000000001110;
    assign weights1[14][645] = 16'b0000000000011001;
    assign weights1[14][646] = 16'b0000000000011101;
    assign weights1[14][647] = 16'b0000000000001011;
    assign weights1[14][648] = 16'b0000000000000010;
    assign weights1[14][649] = 16'b1111111111000001;
    assign weights1[14][650] = 16'b1111111110101101;
    assign weights1[14][651] = 16'b1111111110000100;
    assign weights1[14][652] = 16'b1111111101101100;
    assign weights1[14][653] = 16'b1111111100111110;
    assign weights1[14][654] = 16'b1111111110110000;
    assign weights1[14][655] = 16'b0000000000010000;
    assign weights1[14][656] = 16'b0000000000110101;
    assign weights1[14][657] = 16'b0000000000111011;
    assign weights1[14][658] = 16'b0000000000111000;
    assign weights1[14][659] = 16'b0000000000101111;
    assign weights1[14][660] = 16'b0000000000010011;
    assign weights1[14][661] = 16'b1111111111001100;
    assign weights1[14][662] = 16'b1111111110100100;
    assign weights1[14][663] = 16'b1111111110111001;
    assign weights1[14][664] = 16'b1111111110111101;
    assign weights1[14][665] = 16'b1111111111000000;
    assign weights1[14][666] = 16'b1111111111101011;
    assign weights1[14][667] = 16'b0000000000000000;
    assign weights1[14][668] = 16'b0000000000010110;
    assign weights1[14][669] = 16'b0000000000001110;
    assign weights1[14][670] = 16'b0000000000011010;
    assign weights1[14][671] = 16'b0000000000010100;
    assign weights1[14][672] = 16'b0000000000001010;
    assign weights1[14][673] = 16'b0000000000000101;
    assign weights1[14][674] = 16'b0000000000000010;
    assign weights1[14][675] = 16'b1111111111110111;
    assign weights1[14][676] = 16'b1111111111011110;
    assign weights1[14][677] = 16'b1111111110110011;
    assign weights1[14][678] = 16'b1111111110100010;
    assign weights1[14][679] = 16'b1111111101111110;
    assign weights1[14][680] = 16'b1111111101001111;
    assign weights1[14][681] = 16'b1111111110000101;
    assign weights1[14][682] = 16'b0000000000010010;
    assign weights1[14][683] = 16'b0000000000110111;
    assign weights1[14][684] = 16'b0000000000110011;
    assign weights1[14][685] = 16'b0000000000010110;
    assign weights1[14][686] = 16'b0000000000001101;
    assign weights1[14][687] = 16'b0000000001000011;
    assign weights1[14][688] = 16'b1111111111100000;
    assign weights1[14][689] = 16'b1111111110101101;
    assign weights1[14][690] = 16'b1111111101101111;
    assign weights1[14][691] = 16'b1111111110101001;
    assign weights1[14][692] = 16'b1111111110111110;
    assign weights1[14][693] = 16'b1111111111000000;
    assign weights1[14][694] = 16'b1111111111011000;
    assign weights1[14][695] = 16'b1111111111101001;
    assign weights1[14][696] = 16'b1111111111111001;
    assign weights1[14][697] = 16'b0000000000000001;
    assign weights1[14][698] = 16'b0000000000001010;
    assign weights1[14][699] = 16'b0000000000001100;
    assign weights1[14][700] = 16'b1111111111111100;
    assign weights1[14][701] = 16'b1111111111110011;
    assign weights1[14][702] = 16'b1111111111101100;
    assign weights1[14][703] = 16'b1111111111010010;
    assign weights1[14][704] = 16'b1111111111001000;
    assign weights1[14][705] = 16'b1111111110110001;
    assign weights1[14][706] = 16'b1111111110000110;
    assign weights1[14][707] = 16'b1111111101111110;
    assign weights1[14][708] = 16'b1111111101110101;
    assign weights1[14][709] = 16'b1111111111001010;
    assign weights1[14][710] = 16'b0000000000000000;
    assign weights1[14][711] = 16'b0000000000100100;
    assign weights1[14][712] = 16'b0000000000101000;
    assign weights1[14][713] = 16'b0000000000011010;
    assign weights1[14][714] = 16'b0000000000110110;
    assign weights1[14][715] = 16'b0000000000111001;
    assign weights1[14][716] = 16'b0000000000001100;
    assign weights1[14][717] = 16'b1111111111000100;
    assign weights1[14][718] = 16'b1111111110100000;
    assign weights1[14][719] = 16'b1111111110101101;
    assign weights1[14][720] = 16'b1111111110111100;
    assign weights1[14][721] = 16'b1111111110110111;
    assign weights1[14][722] = 16'b1111111111001100;
    assign weights1[14][723] = 16'b1111111111011100;
    assign weights1[14][724] = 16'b1111111111101011;
    assign weights1[14][725] = 16'b0000000000000000;
    assign weights1[14][726] = 16'b0000000000001001;
    assign weights1[14][727] = 16'b0000000000001000;
    assign weights1[14][728] = 16'b1111111111110111;
    assign weights1[14][729] = 16'b1111111111101011;
    assign weights1[14][730] = 16'b1111111111100000;
    assign weights1[14][731] = 16'b1111111111001110;
    assign weights1[14][732] = 16'b1111111110111001;
    assign weights1[14][733] = 16'b1111111110110100;
    assign weights1[14][734] = 16'b1111111110100011;
    assign weights1[14][735] = 16'b1111111110010101;
    assign weights1[14][736] = 16'b1111111110111110;
    assign weights1[14][737] = 16'b1111111111111101;
    assign weights1[14][738] = 16'b0000000000011110;
    assign weights1[14][739] = 16'b0000000000101001;
    assign weights1[14][740] = 16'b0000000000101100;
    assign weights1[14][741] = 16'b0000000000100101;
    assign weights1[14][742] = 16'b0000000000101000;
    assign weights1[14][743] = 16'b0000000000010001;
    assign weights1[14][744] = 16'b1111111111101011;
    assign weights1[14][745] = 16'b1111111111001100;
    assign weights1[14][746] = 16'b1111111110101111;
    assign weights1[14][747] = 16'b1111111110111010;
    assign weights1[14][748] = 16'b1111111111000011;
    assign weights1[14][749] = 16'b1111111111000001;
    assign weights1[14][750] = 16'b1111111111011001;
    assign weights1[14][751] = 16'b1111111111011110;
    assign weights1[14][752] = 16'b1111111111101111;
    assign weights1[14][753] = 16'b1111111111111110;
    assign weights1[14][754] = 16'b0000000000000111;
    assign weights1[14][755] = 16'b0000000000000010;
    assign weights1[14][756] = 16'b1111111111111010;
    assign weights1[14][757] = 16'b1111111111110010;
    assign weights1[14][758] = 16'b1111111111100010;
    assign weights1[14][759] = 16'b1111111111001100;
    assign weights1[14][760] = 16'b1111111110110010;
    assign weights1[14][761] = 16'b1111111110100011;
    assign weights1[14][762] = 16'b1111111110010111;
    assign weights1[14][763] = 16'b1111111110100101;
    assign weights1[14][764] = 16'b1111111111100000;
    assign weights1[14][765] = 16'b0000000000000000;
    assign weights1[14][766] = 16'b0000000000101000;
    assign weights1[14][767] = 16'b0000000000100100;
    assign weights1[14][768] = 16'b0000000000110010;
    assign weights1[14][769] = 16'b0000000000101111;
    assign weights1[14][770] = 16'b0000000000011110;
    assign weights1[14][771] = 16'b0000000000010000;
    assign weights1[14][772] = 16'b0000000000000110;
    assign weights1[14][773] = 16'b1111111111010011;
    assign weights1[14][774] = 16'b1111111111000101;
    assign weights1[14][775] = 16'b1111111110110110;
    assign weights1[14][776] = 16'b1111111111000000;
    assign weights1[14][777] = 16'b1111111111001001;
    assign weights1[14][778] = 16'b1111111111011010;
    assign weights1[14][779] = 16'b1111111111100011;
    assign weights1[14][780] = 16'b1111111111110001;
    assign weights1[14][781] = 16'b0000000000000001;
    assign weights1[14][782] = 16'b0000000000001000;
    assign weights1[14][783] = 16'b0000000000001000;
    assign weights1[15][0] = 16'b0000000000000000;
    assign weights1[15][1] = 16'b0000000000000000;
    assign weights1[15][2] = 16'b0000000000000000;
    assign weights1[15][3] = 16'b0000000000000000;
    assign weights1[15][4] = 16'b0000000000000000;
    assign weights1[15][5] = 16'b1111111111111110;
    assign weights1[15][6] = 16'b0000000000000000;
    assign weights1[15][7] = 16'b0000000000000000;
    assign weights1[15][8] = 16'b0000000000000000;
    assign weights1[15][9] = 16'b0000000000000000;
    assign weights1[15][10] = 16'b0000000000000010;
    assign weights1[15][11] = 16'b0000000000000010;
    assign weights1[15][12] = 16'b0000000000000100;
    assign weights1[15][13] = 16'b0000000000000110;
    assign weights1[15][14] = 16'b0000000000001001;
    assign weights1[15][15] = 16'b0000000000001010;
    assign weights1[15][16] = 16'b0000000000000110;
    assign weights1[15][17] = 16'b0000000000001000;
    assign weights1[15][18] = 16'b0000000000000010;
    assign weights1[15][19] = 16'b1111111111111111;
    assign weights1[15][20] = 16'b0000000000000011;
    assign weights1[15][21] = 16'b0000000000000100;
    assign weights1[15][22] = 16'b0000000000000011;
    assign weights1[15][23] = 16'b0000000000000001;
    assign weights1[15][24] = 16'b0000000000000000;
    assign weights1[15][25] = 16'b1111111111111111;
    assign weights1[15][26] = 16'b0000000000000000;
    assign weights1[15][27] = 16'b0000000000000000;
    assign weights1[15][28] = 16'b0000000000000000;
    assign weights1[15][29] = 16'b0000000000000000;
    assign weights1[15][30] = 16'b0000000000000000;
    assign weights1[15][31] = 16'b1111111111111111;
    assign weights1[15][32] = 16'b1111111111111110;
    assign weights1[15][33] = 16'b1111111111111110;
    assign weights1[15][34] = 16'b1111111111111100;
    assign weights1[15][35] = 16'b1111111111111111;
    assign weights1[15][36] = 16'b1111111111111111;
    assign weights1[15][37] = 16'b0000000000000010;
    assign weights1[15][38] = 16'b0000000000000001;
    assign weights1[15][39] = 16'b0000000000000100;
    assign weights1[15][40] = 16'b0000000000001001;
    assign weights1[15][41] = 16'b0000000000001110;
    assign weights1[15][42] = 16'b0000000000001100;
    assign weights1[15][43] = 16'b0000000000001101;
    assign weights1[15][44] = 16'b0000000000001010;
    assign weights1[15][45] = 16'b0000000000001000;
    assign weights1[15][46] = 16'b0000000000001101;
    assign weights1[15][47] = 16'b0000000000000101;
    assign weights1[15][48] = 16'b0000000000000110;
    assign weights1[15][49] = 16'b0000000000001010;
    assign weights1[15][50] = 16'b0000000000000111;
    assign weights1[15][51] = 16'b0000000000000100;
    assign weights1[15][52] = 16'b1111111111111111;
    assign weights1[15][53] = 16'b1111111111111110;
    assign weights1[15][54] = 16'b1111111111111110;
    assign weights1[15][55] = 16'b0000000000000001;
    assign weights1[15][56] = 16'b0000000000000000;
    assign weights1[15][57] = 16'b0000000000000000;
    assign weights1[15][58] = 16'b0000000000000000;
    assign weights1[15][59] = 16'b1111111111111111;
    assign weights1[15][60] = 16'b1111111111111110;
    assign weights1[15][61] = 16'b1111111111111100;
    assign weights1[15][62] = 16'b1111111111111101;
    assign weights1[15][63] = 16'b0000000000000000;
    assign weights1[15][64] = 16'b1111111111111110;
    assign weights1[15][65] = 16'b1111111111111111;
    assign weights1[15][66] = 16'b0000000000000001;
    assign weights1[15][67] = 16'b0000000000000101;
    assign weights1[15][68] = 16'b0000000000001111;
    assign weights1[15][69] = 16'b0000000000010001;
    assign weights1[15][70] = 16'b0000000000001000;
    assign weights1[15][71] = 16'b0000000000001000;
    assign weights1[15][72] = 16'b0000000000000100;
    assign weights1[15][73] = 16'b0000000000001001;
    assign weights1[15][74] = 16'b0000000000001110;
    assign weights1[15][75] = 16'b0000000000001111;
    assign weights1[15][76] = 16'b0000000000000000;
    assign weights1[15][77] = 16'b0000000000000101;
    assign weights1[15][78] = 16'b0000000000001000;
    assign weights1[15][79] = 16'b0000000000001010;
    assign weights1[15][80] = 16'b0000000000000101;
    assign weights1[15][81] = 16'b0000000000000001;
    assign weights1[15][82] = 16'b0000000000000001;
    assign weights1[15][83] = 16'b0000000000000001;
    assign weights1[15][84] = 16'b1111111111111111;
    assign weights1[15][85] = 16'b1111111111111111;
    assign weights1[15][86] = 16'b1111111111111110;
    assign weights1[15][87] = 16'b1111111111111101;
    assign weights1[15][88] = 16'b1111111111111011;
    assign weights1[15][89] = 16'b1111111111110010;
    assign weights1[15][90] = 16'b1111111111110100;
    assign weights1[15][91] = 16'b1111111111111101;
    assign weights1[15][92] = 16'b1111111111111111;
    assign weights1[15][93] = 16'b1111111111111011;
    assign weights1[15][94] = 16'b1111111111111011;
    assign weights1[15][95] = 16'b1111111111110101;
    assign weights1[15][96] = 16'b1111111111110100;
    assign weights1[15][97] = 16'b1111111111110111;
    assign weights1[15][98] = 16'b1111111111110000;
    assign weights1[15][99] = 16'b1111111111111001;
    assign weights1[15][100] = 16'b1111111111111100;
    assign weights1[15][101] = 16'b1111111111110001;
    assign weights1[15][102] = 16'b1111111111110111;
    assign weights1[15][103] = 16'b1111111111111011;
    assign weights1[15][104] = 16'b1111111111110100;
    assign weights1[15][105] = 16'b1111111111111000;
    assign weights1[15][106] = 16'b0000000000000101;
    assign weights1[15][107] = 16'b0000000000000111;
    assign weights1[15][108] = 16'b0000000000000011;
    assign weights1[15][109] = 16'b0000000000000100;
    assign weights1[15][110] = 16'b1111111111111101;
    assign weights1[15][111] = 16'b1111111111111110;
    assign weights1[15][112] = 16'b1111111111111111;
    assign weights1[15][113] = 16'b1111111111111110;
    assign weights1[15][114] = 16'b1111111111111101;
    assign weights1[15][115] = 16'b1111111111111101;
    assign weights1[15][116] = 16'b1111111111111100;
    assign weights1[15][117] = 16'b1111111111111010;
    assign weights1[15][118] = 16'b1111111111110101;
    assign weights1[15][119] = 16'b1111111111110111;
    assign weights1[15][120] = 16'b1111111111111010;
    assign weights1[15][121] = 16'b0000000000000110;
    assign weights1[15][122] = 16'b0000000000001000;
    assign weights1[15][123] = 16'b1111111111111100;
    assign weights1[15][124] = 16'b1111111111111110;
    assign weights1[15][125] = 16'b0000000000000111;
    assign weights1[15][126] = 16'b0000000000000111;
    assign weights1[15][127] = 16'b1111111111111000;
    assign weights1[15][128] = 16'b1111111111111000;
    assign weights1[15][129] = 16'b1111111111111001;
    assign weights1[15][130] = 16'b1111111111110000;
    assign weights1[15][131] = 16'b1111111111111110;
    assign weights1[15][132] = 16'b1111111111101011;
    assign weights1[15][133] = 16'b1111111111110100;
    assign weights1[15][134] = 16'b0000000000000000;
    assign weights1[15][135] = 16'b1111111111111001;
    assign weights1[15][136] = 16'b1111111111111011;
    assign weights1[15][137] = 16'b1111111111111001;
    assign weights1[15][138] = 16'b1111111111111101;
    assign weights1[15][139] = 16'b1111111111111100;
    assign weights1[15][140] = 16'b1111111111111110;
    assign weights1[15][141] = 16'b1111111111111010;
    assign weights1[15][142] = 16'b1111111111111011;
    assign weights1[15][143] = 16'b1111111111110100;
    assign weights1[15][144] = 16'b1111111111111001;
    assign weights1[15][145] = 16'b1111111111110101;
    assign weights1[15][146] = 16'b0000000000000000;
    assign weights1[15][147] = 16'b1111111111111001;
    assign weights1[15][148] = 16'b1111111111100011;
    assign weights1[15][149] = 16'b0000000000000100;
    assign weights1[15][150] = 16'b1111111111111110;
    assign weights1[15][151] = 16'b0000000000010011;
    assign weights1[15][152] = 16'b0000000000000111;
    assign weights1[15][153] = 16'b1111111111011100;
    assign weights1[15][154] = 16'b1111111111111000;
    assign weights1[15][155] = 16'b1111111111111100;
    assign weights1[15][156] = 16'b0000000000001100;
    assign weights1[15][157] = 16'b0000000000001100;
    assign weights1[15][158] = 16'b0000000000001101;
    assign weights1[15][159] = 16'b0000000000000000;
    assign weights1[15][160] = 16'b0000000000001111;
    assign weights1[15][161] = 16'b0000000000000101;
    assign weights1[15][162] = 16'b1111111111110111;
    assign weights1[15][163] = 16'b1111111111110010;
    assign weights1[15][164] = 16'b1111111111101011;
    assign weights1[15][165] = 16'b1111111111110000;
    assign weights1[15][166] = 16'b1111111111111000;
    assign weights1[15][167] = 16'b1111111111111010;
    assign weights1[15][168] = 16'b1111111111111100;
    assign weights1[15][169] = 16'b1111111111111000;
    assign weights1[15][170] = 16'b1111111111110111;
    assign weights1[15][171] = 16'b1111111111111001;
    assign weights1[15][172] = 16'b1111111111101101;
    assign weights1[15][173] = 16'b1111111111011011;
    assign weights1[15][174] = 16'b0000000000001101;
    assign weights1[15][175] = 16'b1111111111101110;
    assign weights1[15][176] = 16'b1111111111110010;
    assign weights1[15][177] = 16'b0000000000001001;
    assign weights1[15][178] = 16'b0000000000100000;
    assign weights1[15][179] = 16'b1111111111110000;
    assign weights1[15][180] = 16'b1111111111101101;
    assign weights1[15][181] = 16'b1111111111111110;
    assign weights1[15][182] = 16'b1111111111101001;
    assign weights1[15][183] = 16'b1111111111111110;
    assign weights1[15][184] = 16'b1111111111110110;
    assign weights1[15][185] = 16'b1111111111101111;
    assign weights1[15][186] = 16'b0000000000011011;
    assign weights1[15][187] = 16'b1111111111110111;
    assign weights1[15][188] = 16'b0000000000001110;
    assign weights1[15][189] = 16'b0000000000010100;
    assign weights1[15][190] = 16'b0000000000001100;
    assign weights1[15][191] = 16'b1111111111111011;
    assign weights1[15][192] = 16'b0000000000001101;
    assign weights1[15][193] = 16'b1111111111110100;
    assign weights1[15][194] = 16'b0000000000000001;
    assign weights1[15][195] = 16'b1111111111111111;
    assign weights1[15][196] = 16'b1111111111111000;
    assign weights1[15][197] = 16'b1111111111110101;
    assign weights1[15][198] = 16'b1111111111110001;
    assign weights1[15][199] = 16'b1111111111101110;
    assign weights1[15][200] = 16'b1111111111110010;
    assign weights1[15][201] = 16'b1111111111111010;
    assign weights1[15][202] = 16'b0000000000001000;
    assign weights1[15][203] = 16'b0000000000000111;
    assign weights1[15][204] = 16'b0000000000001111;
    assign weights1[15][205] = 16'b1111111111110101;
    assign weights1[15][206] = 16'b1111111111110111;
    assign weights1[15][207] = 16'b0000000000000101;
    assign weights1[15][208] = 16'b1111111111111011;
    assign weights1[15][209] = 16'b1111111111110011;
    assign weights1[15][210] = 16'b1111111111111111;
    assign weights1[15][211] = 16'b0000000000010010;
    assign weights1[15][212] = 16'b1111111111111100;
    assign weights1[15][213] = 16'b1111111111111011;
    assign weights1[15][214] = 16'b0000000000001100;
    assign weights1[15][215] = 16'b1111111111110000;
    assign weights1[15][216] = 16'b1111111111111101;
    assign weights1[15][217] = 16'b0000000000011001;
    assign weights1[15][218] = 16'b1111111111110010;
    assign weights1[15][219] = 16'b1111111111101100;
    assign weights1[15][220] = 16'b1111111111110110;
    assign weights1[15][221] = 16'b1111111111111011;
    assign weights1[15][222] = 16'b0000000000000010;
    assign weights1[15][223] = 16'b1111111111111111;
    assign weights1[15][224] = 16'b1111111111111001;
    assign weights1[15][225] = 16'b1111111111111011;
    assign weights1[15][226] = 16'b1111111111110011;
    assign weights1[15][227] = 16'b1111111111101110;
    assign weights1[15][228] = 16'b1111111111111000;
    assign weights1[15][229] = 16'b1111111111101000;
    assign weights1[15][230] = 16'b0000000000010001;
    assign weights1[15][231] = 16'b0000000000001011;
    assign weights1[15][232] = 16'b1111111111010001;
    assign weights1[15][233] = 16'b1111111111100100;
    assign weights1[15][234] = 16'b1111111111110111;
    assign weights1[15][235] = 16'b1111111111111000;
    assign weights1[15][236] = 16'b0000000000000100;
    assign weights1[15][237] = 16'b0000000000010001;
    assign weights1[15][238] = 16'b1111111111110101;
    assign weights1[15][239] = 16'b1111111111100011;
    assign weights1[15][240] = 16'b0000000000001001;
    assign weights1[15][241] = 16'b0000000000000100;
    assign weights1[15][242] = 16'b1111111111110101;
    assign weights1[15][243] = 16'b0000000000001000;
    assign weights1[15][244] = 16'b0000000000000100;
    assign weights1[15][245] = 16'b1111111111101000;
    assign weights1[15][246] = 16'b0000000000000010;
    assign weights1[15][247] = 16'b1111111111101011;
    assign weights1[15][248] = 16'b1111111111110011;
    assign weights1[15][249] = 16'b1111111111111011;
    assign weights1[15][250] = 16'b0000000000000000;
    assign weights1[15][251] = 16'b1111111111111111;
    assign weights1[15][252] = 16'b1111111111111111;
    assign weights1[15][253] = 16'b1111111111110111;
    assign weights1[15][254] = 16'b1111111111101110;
    assign weights1[15][255] = 16'b1111111111110000;
    assign weights1[15][256] = 16'b1111111111110010;
    assign weights1[15][257] = 16'b1111111111100010;
    assign weights1[15][258] = 16'b1111111111101011;
    assign weights1[15][259] = 16'b1111111111111000;
    assign weights1[15][260] = 16'b1111111111111100;
    assign weights1[15][261] = 16'b0000000000000011;
    assign weights1[15][262] = 16'b1111111111110001;
    assign weights1[15][263] = 16'b1111111111111010;
    assign weights1[15][264] = 16'b1111111111111100;
    assign weights1[15][265] = 16'b1111111111111001;
    assign weights1[15][266] = 16'b1111111111110000;
    assign weights1[15][267] = 16'b1111111111111111;
    assign weights1[15][268] = 16'b0000000000000001;
    assign weights1[15][269] = 16'b1111111111101001;
    assign weights1[15][270] = 16'b0000000000000001;
    assign weights1[15][271] = 16'b1111111111110010;
    assign weights1[15][272] = 16'b0000000000000000;
    assign weights1[15][273] = 16'b0000000000000100;
    assign weights1[15][274] = 16'b0000000000001001;
    assign weights1[15][275] = 16'b0000000000000100;
    assign weights1[15][276] = 16'b1111111111101110;
    assign weights1[15][277] = 16'b0000000000000101;
    assign weights1[15][278] = 16'b0000000000010000;
    assign weights1[15][279] = 16'b0000000000000100;
    assign weights1[15][280] = 16'b1111111111111000;
    assign weights1[15][281] = 16'b1111111111101110;
    assign weights1[15][282] = 16'b1111111111111000;
    assign weights1[15][283] = 16'b0000000000000001;
    assign weights1[15][284] = 16'b1111111111111110;
    assign weights1[15][285] = 16'b1111111111110001;
    assign weights1[15][286] = 16'b1111111111111101;
    assign weights1[15][287] = 16'b1111111111111010;
    assign weights1[15][288] = 16'b1111111111101001;
    assign weights1[15][289] = 16'b0000000000001010;
    assign weights1[15][290] = 16'b1111111111101110;
    assign weights1[15][291] = 16'b1111111111110110;
    assign weights1[15][292] = 16'b1111111111111010;
    assign weights1[15][293] = 16'b1111111111111101;
    assign weights1[15][294] = 16'b1111111111111000;
    assign weights1[15][295] = 16'b1111111111110110;
    assign weights1[15][296] = 16'b0000000000001010;
    assign weights1[15][297] = 16'b1111111111111100;
    assign weights1[15][298] = 16'b0000000000000000;
    assign weights1[15][299] = 16'b1111111111111101;
    assign weights1[15][300] = 16'b1111111111111111;
    assign weights1[15][301] = 16'b1111111111111100;
    assign weights1[15][302] = 16'b1111111111111000;
    assign weights1[15][303] = 16'b0000000000000000;
    assign weights1[15][304] = 16'b1111111111100111;
    assign weights1[15][305] = 16'b1111111111111010;
    assign weights1[15][306] = 16'b1111111111110111;
    assign weights1[15][307] = 16'b1111111111110110;
    assign weights1[15][308] = 16'b1111111111110100;
    assign weights1[15][309] = 16'b1111111111110010;
    assign weights1[15][310] = 16'b1111111111110001;
    assign weights1[15][311] = 16'b1111111111110100;
    assign weights1[15][312] = 16'b0000000000000100;
    assign weights1[15][313] = 16'b1111111111101111;
    assign weights1[15][314] = 16'b0000000000001110;
    assign weights1[15][315] = 16'b1111111111100101;
    assign weights1[15][316] = 16'b1111111111101110;
    assign weights1[15][317] = 16'b1111111111110100;
    assign weights1[15][318] = 16'b1111111111110111;
    assign weights1[15][319] = 16'b1111111111110110;
    assign weights1[15][320] = 16'b1111111111101110;
    assign weights1[15][321] = 16'b1111111111111011;
    assign weights1[15][322] = 16'b1111111111100001;
    assign weights1[15][323] = 16'b1111111111111000;
    assign weights1[15][324] = 16'b1111111111100001;
    assign weights1[15][325] = 16'b1111111111110101;
    assign weights1[15][326] = 16'b1111111111101101;
    assign weights1[15][327] = 16'b0000000000000001;
    assign weights1[15][328] = 16'b1111111111110001;
    assign weights1[15][329] = 16'b0000000000000000;
    assign weights1[15][330] = 16'b1111111111110101;
    assign weights1[15][331] = 16'b1111111111101100;
    assign weights1[15][332] = 16'b1111111111100111;
    assign weights1[15][333] = 16'b1111111111101100;
    assign weights1[15][334] = 16'b1111111111110100;
    assign weights1[15][335] = 16'b1111111111111001;
    assign weights1[15][336] = 16'b1111111111110111;
    assign weights1[15][337] = 16'b1111111111110101;
    assign weights1[15][338] = 16'b1111111111111101;
    assign weights1[15][339] = 16'b1111111111110011;
    assign weights1[15][340] = 16'b1111111111111111;
    assign weights1[15][341] = 16'b1111111111111001;
    assign weights1[15][342] = 16'b1111111111110000;
    assign weights1[15][343] = 16'b1111111111101001;
    assign weights1[15][344] = 16'b0000000000000110;
    assign weights1[15][345] = 16'b0000000000000100;
    assign weights1[15][346] = 16'b1111111111110001;
    assign weights1[15][347] = 16'b1111111111101011;
    assign weights1[15][348] = 16'b0000000000000011;
    assign weights1[15][349] = 16'b1111111111101101;
    assign weights1[15][350] = 16'b1111111111101110;
    assign weights1[15][351] = 16'b1111111111110010;
    assign weights1[15][352] = 16'b1111111111110100;
    assign weights1[15][353] = 16'b1111111111100000;
    assign weights1[15][354] = 16'b1111111111011011;
    assign weights1[15][355] = 16'b1111111111111000;
    assign weights1[15][356] = 16'b1111111111100101;
    assign weights1[15][357] = 16'b1111111111110100;
    assign weights1[15][358] = 16'b1111111111100001;
    assign weights1[15][359] = 16'b1111111111011100;
    assign weights1[15][360] = 16'b1111111111011000;
    assign weights1[15][361] = 16'b1111111111101100;
    assign weights1[15][362] = 16'b1111111111101011;
    assign weights1[15][363] = 16'b1111111111110010;
    assign weights1[15][364] = 16'b1111111111101110;
    assign weights1[15][365] = 16'b0000000000000000;
    assign weights1[15][366] = 16'b1111111111111000;
    assign weights1[15][367] = 16'b1111111111110010;
    assign weights1[15][368] = 16'b1111111111110110;
    assign weights1[15][369] = 16'b1111111111100000;
    assign weights1[15][370] = 16'b0000000000000011;
    assign weights1[15][371] = 16'b1111111111110111;
    assign weights1[15][372] = 16'b1111111111100000;
    assign weights1[15][373] = 16'b1111111111100010;
    assign weights1[15][374] = 16'b1111111111110000;
    assign weights1[15][375] = 16'b1111111111100110;
    assign weights1[15][376] = 16'b1111111111101111;
    assign weights1[15][377] = 16'b0000000000001010;
    assign weights1[15][378] = 16'b0000000000000011;
    assign weights1[15][379] = 16'b1111111111101000;
    assign weights1[15][380] = 16'b1111111111110000;
    assign weights1[15][381] = 16'b1111111111111001;
    assign weights1[15][382] = 16'b0000000000000000;
    assign weights1[15][383] = 16'b1111111111101111;
    assign weights1[15][384] = 16'b1111111111100111;
    assign weights1[15][385] = 16'b1111111111010110;
    assign weights1[15][386] = 16'b1111111111011011;
    assign weights1[15][387] = 16'b1111111111011011;
    assign weights1[15][388] = 16'b1111111111011010;
    assign weights1[15][389] = 16'b1111111111110001;
    assign weights1[15][390] = 16'b1111111111101100;
    assign weights1[15][391] = 16'b1111111111111000;
    assign weights1[15][392] = 16'b1111111111110111;
    assign weights1[15][393] = 16'b1111111111111111;
    assign weights1[15][394] = 16'b1111111111110000;
    assign weights1[15][395] = 16'b1111111111101010;
    assign weights1[15][396] = 16'b0000000000010010;
    assign weights1[15][397] = 16'b1111111111100010;
    assign weights1[15][398] = 16'b1111111111101010;
    assign weights1[15][399] = 16'b1111111111101001;
    assign weights1[15][400] = 16'b1111111111100110;
    assign weights1[15][401] = 16'b1111111111110101;
    assign weights1[15][402] = 16'b1111111111111110;
    assign weights1[15][403] = 16'b1111111111110000;
    assign weights1[15][404] = 16'b1111111111101100;
    assign weights1[15][405] = 16'b1111111111110001;
    assign weights1[15][406] = 16'b1111111111111100;
    assign weights1[15][407] = 16'b0000000000001011;
    assign weights1[15][408] = 16'b1111111111110011;
    assign weights1[15][409] = 16'b1111111111101001;
    assign weights1[15][410] = 16'b1111111111100100;
    assign weights1[15][411] = 16'b1111111111110110;
    assign weights1[15][412] = 16'b1111111111101110;
    assign weights1[15][413] = 16'b1111111111101000;
    assign weights1[15][414] = 16'b1111111111001000;
    assign weights1[15][415] = 16'b1111111111011010;
    assign weights1[15][416] = 16'b1111111111100100;
    assign weights1[15][417] = 16'b1111111111100010;
    assign weights1[15][418] = 16'b1111111111100111;
    assign weights1[15][419] = 16'b0000000000000101;
    assign weights1[15][420] = 16'b1111111111111001;
    assign weights1[15][421] = 16'b0000000000000101;
    assign weights1[15][422] = 16'b1111111111101110;
    assign weights1[15][423] = 16'b1111111111110001;
    assign weights1[15][424] = 16'b1111111111111101;
    assign weights1[15][425] = 16'b1111111111110010;
    assign weights1[15][426] = 16'b1111111111110000;
    assign weights1[15][427] = 16'b1111111111101010;
    assign weights1[15][428] = 16'b0000000000001010;
    assign weights1[15][429] = 16'b1111111111101100;
    assign weights1[15][430] = 16'b1111111111110111;
    assign weights1[15][431] = 16'b0000000000001000;
    assign weights1[15][432] = 16'b0000000000001010;
    assign weights1[15][433] = 16'b1111111111110111;
    assign weights1[15][434] = 16'b1111111111110011;
    assign weights1[15][435] = 16'b0000000000001111;
    assign weights1[15][436] = 16'b0000000000000010;
    assign weights1[15][437] = 16'b1111111111111100;
    assign weights1[15][438] = 16'b1111111111010100;
    assign weights1[15][439] = 16'b1111111111101001;
    assign weights1[15][440] = 16'b1111111111100000;
    assign weights1[15][441] = 16'b1111111111101110;
    assign weights1[15][442] = 16'b1111111111100000;
    assign weights1[15][443] = 16'b1111111111101010;
    assign weights1[15][444] = 16'b1111111111011100;
    assign weights1[15][445] = 16'b1111111111010111;
    assign weights1[15][446] = 16'b1111111111111110;
    assign weights1[15][447] = 16'b0000000000011011;
    assign weights1[15][448] = 16'b1111111111110000;
    assign weights1[15][449] = 16'b1111111111101111;
    assign weights1[15][450] = 16'b1111111111101001;
    assign weights1[15][451] = 16'b1111111111100110;
    assign weights1[15][452] = 16'b1111111111101101;
    assign weights1[15][453] = 16'b1111111111100010;
    assign weights1[15][454] = 16'b1111111111111100;
    assign weights1[15][455] = 16'b1111111111111111;
    assign weights1[15][456] = 16'b0000000000001000;
    assign weights1[15][457] = 16'b0000000000010100;
    assign weights1[15][458] = 16'b0000000000001010;
    assign weights1[15][459] = 16'b1111111111111100;
    assign weights1[15][460] = 16'b1111111111110100;
    assign weights1[15][461] = 16'b1111111111110010;
    assign weights1[15][462] = 16'b1111111111110011;
    assign weights1[15][463] = 16'b1111111111110011;
    assign weights1[15][464] = 16'b1111111111101110;
    assign weights1[15][465] = 16'b1111111111111000;
    assign weights1[15][466] = 16'b1111111111111100;
    assign weights1[15][467] = 16'b1111111111111101;
    assign weights1[15][468] = 16'b1111111111100000;
    assign weights1[15][469] = 16'b1111111111110011;
    assign weights1[15][470] = 16'b1111111111101000;
    assign weights1[15][471] = 16'b1111111111110001;
    assign weights1[15][472] = 16'b1111111111101111;
    assign weights1[15][473] = 16'b1111111111110010;
    assign weights1[15][474] = 16'b0000000000100000;
    assign weights1[15][475] = 16'b0000000000101001;
    assign weights1[15][476] = 16'b1111111111110001;
    assign weights1[15][477] = 16'b1111111111101011;
    assign weights1[15][478] = 16'b1111111111110001;
    assign weights1[15][479] = 16'b1111111111010100;
    assign weights1[15][480] = 16'b1111111111011100;
    assign weights1[15][481] = 16'b1111111111101011;
    assign weights1[15][482] = 16'b0000000000001001;
    assign weights1[15][483] = 16'b0000000000000000;
    assign weights1[15][484] = 16'b1111111111110101;
    assign weights1[15][485] = 16'b1111111111111111;
    assign weights1[15][486] = 16'b1111111111111111;
    assign weights1[15][487] = 16'b1111111111110000;
    assign weights1[15][488] = 16'b1111111111111110;
    assign weights1[15][489] = 16'b1111111111111010;
    assign weights1[15][490] = 16'b1111111111111010;
    assign weights1[15][491] = 16'b1111111111101011;
    assign weights1[15][492] = 16'b1111111111111100;
    assign weights1[15][493] = 16'b0000000000000000;
    assign weights1[15][494] = 16'b0000000000000000;
    assign weights1[15][495] = 16'b1111111111111101;
    assign weights1[15][496] = 16'b1111111111100110;
    assign weights1[15][497] = 16'b1111111111111010;
    assign weights1[15][498] = 16'b1111111111101011;
    assign weights1[15][499] = 16'b1111111111101100;
    assign weights1[15][500] = 16'b0000000000000100;
    assign weights1[15][501] = 16'b0000000000011000;
    assign weights1[15][502] = 16'b0000000000100100;
    assign weights1[15][503] = 16'b0000000000111101;
    assign weights1[15][504] = 16'b1111111111111010;
    assign weights1[15][505] = 16'b1111111111101011;
    assign weights1[15][506] = 16'b1111111111111100;
    assign weights1[15][507] = 16'b1111111111110101;
    assign weights1[15][508] = 16'b1111111111111001;
    assign weights1[15][509] = 16'b0000000000000001;
    assign weights1[15][510] = 16'b1111111111111000;
    assign weights1[15][511] = 16'b1111111111111110;
    assign weights1[15][512] = 16'b1111111111111110;
    assign weights1[15][513] = 16'b1111111111111110;
    assign weights1[15][514] = 16'b1111111111111010;
    assign weights1[15][515] = 16'b1111111111110100;
    assign weights1[15][516] = 16'b1111111111111001;
    assign weights1[15][517] = 16'b1111111111111010;
    assign weights1[15][518] = 16'b1111111111100000;
    assign weights1[15][519] = 16'b1111111111111001;
    assign weights1[15][520] = 16'b1111111111111000;
    assign weights1[15][521] = 16'b0000000000001101;
    assign weights1[15][522] = 16'b0000000000010000;
    assign weights1[15][523] = 16'b1111111111111110;
    assign weights1[15][524] = 16'b1111111111011010;
    assign weights1[15][525] = 16'b1111111111011100;
    assign weights1[15][526] = 16'b1111111111110101;
    assign weights1[15][527] = 16'b1111111111110000;
    assign weights1[15][528] = 16'b0000000000000010;
    assign weights1[15][529] = 16'b0000000000110011;
    assign weights1[15][530] = 16'b0000000000111000;
    assign weights1[15][531] = 16'b0000000000101110;
    assign weights1[15][532] = 16'b0000000000001000;
    assign weights1[15][533] = 16'b1111111111111100;
    assign weights1[15][534] = 16'b1111111111101111;
    assign weights1[15][535] = 16'b1111111111111100;
    assign weights1[15][536] = 16'b0000000000001000;
    assign weights1[15][537] = 16'b1111111111110111;
    assign weights1[15][538] = 16'b0000000000000001;
    assign weights1[15][539] = 16'b1111111111110101;
    assign weights1[15][540] = 16'b1111111111111101;
    assign weights1[15][541] = 16'b1111111111011110;
    assign weights1[15][542] = 16'b1111111111110100;
    assign weights1[15][543] = 16'b1111111111111110;
    assign weights1[15][544] = 16'b0000000000000111;
    assign weights1[15][545] = 16'b1111111111111011;
    assign weights1[15][546] = 16'b1111111111100011;
    assign weights1[15][547] = 16'b1111111111100110;
    assign weights1[15][548] = 16'b1111111111110001;
    assign weights1[15][549] = 16'b1111111111110001;
    assign weights1[15][550] = 16'b1111111111111010;
    assign weights1[15][551] = 16'b1111111111110010;
    assign weights1[15][552] = 16'b1111111111101000;
    assign weights1[15][553] = 16'b1111111111110110;
    assign weights1[15][554] = 16'b0000000000001101;
    assign weights1[15][555] = 16'b0000000000010101;
    assign weights1[15][556] = 16'b0000000000011110;
    assign weights1[15][557] = 16'b0000000001001000;
    assign weights1[15][558] = 16'b0000000000110110;
    assign weights1[15][559] = 16'b0000000000100100;
    assign weights1[15][560] = 16'b0000000000010111;
    assign weights1[15][561] = 16'b0000000000001110;
    assign weights1[15][562] = 16'b0000000000001110;
    assign weights1[15][563] = 16'b0000000000010010;
    assign weights1[15][564] = 16'b0000000000001111;
    assign weights1[15][565] = 16'b1111111111101111;
    assign weights1[15][566] = 16'b1111111111111110;
    assign weights1[15][567] = 16'b0000000000011011;
    assign weights1[15][568] = 16'b1111111111101001;
    assign weights1[15][569] = 16'b0000000000001001;
    assign weights1[15][570] = 16'b1111111111100110;
    assign weights1[15][571] = 16'b1111111111100101;
    assign weights1[15][572] = 16'b1111111111101000;
    assign weights1[15][573] = 16'b1111111111010001;
    assign weights1[15][574] = 16'b1111111111101101;
    assign weights1[15][575] = 16'b1111111111101000;
    assign weights1[15][576] = 16'b1111111111011101;
    assign weights1[15][577] = 16'b1111111111010010;
    assign weights1[15][578] = 16'b1111111111101010;
    assign weights1[15][579] = 16'b0000000000001010;
    assign weights1[15][580] = 16'b1111111111101011;
    assign weights1[15][581] = 16'b0000000000001110;
    assign weights1[15][582] = 16'b0000000000100001;
    assign weights1[15][583] = 16'b0000000000110110;
    assign weights1[15][584] = 16'b0000000000111110;
    assign weights1[15][585] = 16'b0000000001010011;
    assign weights1[15][586] = 16'b0000000000111000;
    assign weights1[15][587] = 16'b0000000000100111;
    assign weights1[15][588] = 16'b0000000000101000;
    assign weights1[15][589] = 16'b0000000000101101;
    assign weights1[15][590] = 16'b0000000000100001;
    assign weights1[15][591] = 16'b0000000000100100;
    assign weights1[15][592] = 16'b0000000000010100;
    assign weights1[15][593] = 16'b1111111111111000;
    assign weights1[15][594] = 16'b1111111111111100;
    assign weights1[15][595] = 16'b0000000000001001;
    assign weights1[15][596] = 16'b0000000000000000;
    assign weights1[15][597] = 16'b1111111111100110;
    assign weights1[15][598] = 16'b1111111111010000;
    assign weights1[15][599] = 16'b1111111111011100;
    assign weights1[15][600] = 16'b1111111111010100;
    assign weights1[15][601] = 16'b0000000000001001;
    assign weights1[15][602] = 16'b0000000000000000;
    assign weights1[15][603] = 16'b0000000000000011;
    assign weights1[15][604] = 16'b1111111111100111;
    assign weights1[15][605] = 16'b1111111111100010;
    assign weights1[15][606] = 16'b1111111111111001;
    assign weights1[15][607] = 16'b0000000000010011;
    assign weights1[15][608] = 16'b0000000000101011;
    assign weights1[15][609] = 16'b0000000000111001;
    assign weights1[15][610] = 16'b0000000001100001;
    assign weights1[15][611] = 16'b0000000001010001;
    assign weights1[15][612] = 16'b0000000001100010;
    assign weights1[15][613] = 16'b0000000001010110;
    assign weights1[15][614] = 16'b0000000000110011;
    assign weights1[15][615] = 16'b0000000000110000;
    assign weights1[15][616] = 16'b0000000000110011;
    assign weights1[15][617] = 16'b0000000001000010;
    assign weights1[15][618] = 16'b0000000001000011;
    assign weights1[15][619] = 16'b0000000000110000;
    assign weights1[15][620] = 16'b0000000000100001;
    assign weights1[15][621] = 16'b0000000000110101;
    assign weights1[15][622] = 16'b0000000000101100;
    assign weights1[15][623] = 16'b0000000000001100;
    assign weights1[15][624] = 16'b0000000000001001;
    assign weights1[15][625] = 16'b0000000000101111;
    assign weights1[15][626] = 16'b0000000000001000;
    assign weights1[15][627] = 16'b0000000000011011;
    assign weights1[15][628] = 16'b0000000000100010;
    assign weights1[15][629] = 16'b0000000000000000;
    assign weights1[15][630] = 16'b0000000000101001;
    assign weights1[15][631] = 16'b0000000000110110;
    assign weights1[15][632] = 16'b0000000001001010;
    assign weights1[15][633] = 16'b0000000000101111;
    assign weights1[15][634] = 16'b0000000000111010;
    assign weights1[15][635] = 16'b0000000001011011;
    assign weights1[15][636] = 16'b0000000001011101;
    assign weights1[15][637] = 16'b0000000001101011;
    assign weights1[15][638] = 16'b0000000001100000;
    assign weights1[15][639] = 16'b0000000001100010;
    assign weights1[15][640] = 16'b0000000001010000;
    assign weights1[15][641] = 16'b0000000001010001;
    assign weights1[15][642] = 16'b0000000000110100;
    assign weights1[15][643] = 16'b0000000000101010;
    assign weights1[15][644] = 16'b0000000000110010;
    assign weights1[15][645] = 16'b0000000000111111;
    assign weights1[15][646] = 16'b0000000001001011;
    assign weights1[15][647] = 16'b0000000001011011;
    assign weights1[15][648] = 16'b0000000001001100;
    assign weights1[15][649] = 16'b0000000001011011;
    assign weights1[15][650] = 16'b0000000001011100;
    assign weights1[15][651] = 16'b0000000001001100;
    assign weights1[15][652] = 16'b0000000001101010;
    assign weights1[15][653] = 16'b0000000001101010;
    assign weights1[15][654] = 16'b0000000001010100;
    assign weights1[15][655] = 16'b0000000001101100;
    assign weights1[15][656] = 16'b0000000001100101;
    assign weights1[15][657] = 16'b0000000001000001;
    assign weights1[15][658] = 16'b0000000001001110;
    assign weights1[15][659] = 16'b0000000001011110;
    assign weights1[15][660] = 16'b0000000001100010;
    assign weights1[15][661] = 16'b0000000001101010;
    assign weights1[15][662] = 16'b0000000001101000;
    assign weights1[15][663] = 16'b0000000001100011;
    assign weights1[15][664] = 16'b0000000001010100;
    assign weights1[15][665] = 16'b0000000001000001;
    assign weights1[15][666] = 16'b0000000001010011;
    assign weights1[15][667] = 16'b0000000000101111;
    assign weights1[15][668] = 16'b0000000000110011;
    assign weights1[15][669] = 16'b0000000000111101;
    assign weights1[15][670] = 16'b0000000000100101;
    assign weights1[15][671] = 16'b0000000000011010;
    assign weights1[15][672] = 16'b0000000000101010;
    assign weights1[15][673] = 16'b0000000000111010;
    assign weights1[15][674] = 16'b0000000000111010;
    assign weights1[15][675] = 16'b0000000001001111;
    assign weights1[15][676] = 16'b0000000001000110;
    assign weights1[15][677] = 16'b0000000001010000;
    assign weights1[15][678] = 16'b0000000001000100;
    assign weights1[15][679] = 16'b0000000001010011;
    assign weights1[15][680] = 16'b0000000001100010;
    assign weights1[15][681] = 16'b0000000001001111;
    assign weights1[15][682] = 16'b0000000001110000;
    assign weights1[15][683] = 16'b0000000001101101;
    assign weights1[15][684] = 16'b0000000001011110;
    assign weights1[15][685] = 16'b0000000001010000;
    assign weights1[15][686] = 16'b0000000001001000;
    assign weights1[15][687] = 16'b0000000001001100;
    assign weights1[15][688] = 16'b0000000001011011;
    assign weights1[15][689] = 16'b0000000001001001;
    assign weights1[15][690] = 16'b0000000001000111;
    assign weights1[15][691] = 16'b0000000001000100;
    assign weights1[15][692] = 16'b0000000000110111;
    assign weights1[15][693] = 16'b0000000000101100;
    assign weights1[15][694] = 16'b0000000000111010;
    assign weights1[15][695] = 16'b0000000000010110;
    assign weights1[15][696] = 16'b0000000000101100;
    assign weights1[15][697] = 16'b0000000000110010;
    assign weights1[15][698] = 16'b0000000000011111;
    assign weights1[15][699] = 16'b0000000000001001;
    assign weights1[15][700] = 16'b0000000000011000;
    assign weights1[15][701] = 16'b0000000000101011;
    assign weights1[15][702] = 16'b0000000000100101;
    assign weights1[15][703] = 16'b0000000000101110;
    assign weights1[15][704] = 16'b0000000000110001;
    assign weights1[15][705] = 16'b0000000000100011;
    assign weights1[15][706] = 16'b0000000000101101;
    assign weights1[15][707] = 16'b0000000000011110;
    assign weights1[15][708] = 16'b0000000000110100;
    assign weights1[15][709] = 16'b0000000000101001;
    assign weights1[15][710] = 16'b0000000000111111;
    assign weights1[15][711] = 16'b0000000000110111;
    assign weights1[15][712] = 16'b0000000001001010;
    assign weights1[15][713] = 16'b0000000000110100;
    assign weights1[15][714] = 16'b0000000001000101;
    assign weights1[15][715] = 16'b0000000000110111;
    assign weights1[15][716] = 16'b0000000000110011;
    assign weights1[15][717] = 16'b0000000000011111;
    assign weights1[15][718] = 16'b0000000000010110;
    assign weights1[15][719] = 16'b0000000000100001;
    assign weights1[15][720] = 16'b0000000000110011;
    assign weights1[15][721] = 16'b0000000000010100;
    assign weights1[15][722] = 16'b0000000000011001;
    assign weights1[15][723] = 16'b0000000000010110;
    assign weights1[15][724] = 16'b0000000000011110;
    assign weights1[15][725] = 16'b0000000000011110;
    assign weights1[15][726] = 16'b0000000000010000;
    assign weights1[15][727] = 16'b0000000000000010;
    assign weights1[15][728] = 16'b0000000000000100;
    assign weights1[15][729] = 16'b0000000000000111;
    assign weights1[15][730] = 16'b0000000000010000;
    assign weights1[15][731] = 16'b0000000000010110;
    assign weights1[15][732] = 16'b0000000000010100;
    assign weights1[15][733] = 16'b0000000000011101;
    assign weights1[15][734] = 16'b0000000000010101;
    assign weights1[15][735] = 16'b0000000000011010;
    assign weights1[15][736] = 16'b0000000000010010;
    assign weights1[15][737] = 16'b0000000000010010;
    assign weights1[15][738] = 16'b0000000000100000;
    assign weights1[15][739] = 16'b0000000000001110;
    assign weights1[15][740] = 16'b0000000000100011;
    assign weights1[15][741] = 16'b0000000000011011;
    assign weights1[15][742] = 16'b0000000000010111;
    assign weights1[15][743] = 16'b0000000000010001;
    assign weights1[15][744] = 16'b0000000000001110;
    assign weights1[15][745] = 16'b0000000000001111;
    assign weights1[15][746] = 16'b0000000000100011;
    assign weights1[15][747] = 16'b0000000000011001;
    assign weights1[15][748] = 16'b0000000000010101;
    assign weights1[15][749] = 16'b0000000000011111;
    assign weights1[15][750] = 16'b0000000000010111;
    assign weights1[15][751] = 16'b0000000000010100;
    assign weights1[15][752] = 16'b0000000000010100;
    assign weights1[15][753] = 16'b0000000000000010;
    assign weights1[15][754] = 16'b0000000000000110;
    assign weights1[15][755] = 16'b1111111111111100;
    assign weights1[15][756] = 16'b1111111111111011;
    assign weights1[15][757] = 16'b0000000000000001;
    assign weights1[15][758] = 16'b0000000000000001;
    assign weights1[15][759] = 16'b1111111111111111;
    assign weights1[15][760] = 16'b0000000000001010;
    assign weights1[15][761] = 16'b0000000000010111;
    assign weights1[15][762] = 16'b0000000000001100;
    assign weights1[15][763] = 16'b0000000000001110;
    assign weights1[15][764] = 16'b0000000000001101;
    assign weights1[15][765] = 16'b0000000000001100;
    assign weights1[15][766] = 16'b0000000000011010;
    assign weights1[15][767] = 16'b0000000000011100;
    assign weights1[15][768] = 16'b0000000000010010;
    assign weights1[15][769] = 16'b0000000000010010;
    assign weights1[15][770] = 16'b0000000000010101;
    assign weights1[15][771] = 16'b0000000000100011;
    assign weights1[15][772] = 16'b0000000000001111;
    assign weights1[15][773] = 16'b0000000000001000;
    assign weights1[15][774] = 16'b0000000000101010;
    assign weights1[15][775] = 16'b0000000000101001;
    assign weights1[15][776] = 16'b0000000000001100;
    assign weights1[15][777] = 16'b0000000000001001;
    assign weights1[15][778] = 16'b0000000000010010;
    assign weights1[15][779] = 16'b0000000000000111;
    assign weights1[15][780] = 16'b0000000000000101;
    assign weights1[15][781] = 16'b0000000000001001;
    assign weights1[15][782] = 16'b1111111111111110;
    assign weights1[15][783] = 16'b1111111111111001;
    assign weights1[16][0] = 16'b0000000000000000;
    assign weights1[16][1] = 16'b1111111111111111;
    assign weights1[16][2] = 16'b1111111111111101;
    assign weights1[16][3] = 16'b1111111111111010;
    assign weights1[16][4] = 16'b1111111111110001;
    assign weights1[16][5] = 16'b1111111111110001;
    assign weights1[16][6] = 16'b1111111111101010;
    assign weights1[16][7] = 16'b1111111111101000;
    assign weights1[16][8] = 16'b1111111111101011;
    assign weights1[16][9] = 16'b1111111111100000;
    assign weights1[16][10] = 16'b1111111111011011;
    assign weights1[16][11] = 16'b1111111111011001;
    assign weights1[16][12] = 16'b1111111111011100;
    assign weights1[16][13] = 16'b1111111111011010;
    assign weights1[16][14] = 16'b1111111111100001;
    assign weights1[16][15] = 16'b1111111111100000;
    assign weights1[16][16] = 16'b1111111111011100;
    assign weights1[16][17] = 16'b1111111111101001;
    assign weights1[16][18] = 16'b1111111111100111;
    assign weights1[16][19] = 16'b1111111111100110;
    assign weights1[16][20] = 16'b1111111111101111;
    assign weights1[16][21] = 16'b1111111111101101;
    assign weights1[16][22] = 16'b1111111111110110;
    assign weights1[16][23] = 16'b1111111111111000;
    assign weights1[16][24] = 16'b1111111111110101;
    assign weights1[16][25] = 16'b1111111111111001;
    assign weights1[16][26] = 16'b1111111111111101;
    assign weights1[16][27] = 16'b1111111111111111;
    assign weights1[16][28] = 16'b0000000000000000;
    assign weights1[16][29] = 16'b1111111111111101;
    assign weights1[16][30] = 16'b1111111111110111;
    assign weights1[16][31] = 16'b1111111111110001;
    assign weights1[16][32] = 16'b1111111111101010;
    assign weights1[16][33] = 16'b1111111111100101;
    assign weights1[16][34] = 16'b1111111111100000;
    assign weights1[16][35] = 16'b1111111111011000;
    assign weights1[16][36] = 16'b1111111111011110;
    assign weights1[16][37] = 16'b1111111111001111;
    assign weights1[16][38] = 16'b1111111111001010;
    assign weights1[16][39] = 16'b1111111111001001;
    assign weights1[16][40] = 16'b1111111111000110;
    assign weights1[16][41] = 16'b1111111111000111;
    assign weights1[16][42] = 16'b1111111111001001;
    assign weights1[16][43] = 16'b1111111111000100;
    assign weights1[16][44] = 16'b1111111111000101;
    assign weights1[16][45] = 16'b1111111111010001;
    assign weights1[16][46] = 16'b1111111111010111;
    assign weights1[16][47] = 16'b1111111111010111;
    assign weights1[16][48] = 16'b1111111111011000;
    assign weights1[16][49] = 16'b1111111111011110;
    assign weights1[16][50] = 16'b1111111111100001;
    assign weights1[16][51] = 16'b1111111111101011;
    assign weights1[16][52] = 16'b1111111111101100;
    assign weights1[16][53] = 16'b1111111111110011;
    assign weights1[16][54] = 16'b1111111111111100;
    assign weights1[16][55] = 16'b1111111111111110;
    assign weights1[16][56] = 16'b0000000000000000;
    assign weights1[16][57] = 16'b1111111111111011;
    assign weights1[16][58] = 16'b1111111111101110;
    assign weights1[16][59] = 16'b1111111111101011;
    assign weights1[16][60] = 16'b1111111111100101;
    assign weights1[16][61] = 16'b1111111111011101;
    assign weights1[16][62] = 16'b1111111111010000;
    assign weights1[16][63] = 16'b1111111111001000;
    assign weights1[16][64] = 16'b1111111111001010;
    assign weights1[16][65] = 16'b1111111110111101;
    assign weights1[16][66] = 16'b1111111110111000;
    assign weights1[16][67] = 16'b1111111110101010;
    assign weights1[16][68] = 16'b1111111110100011;
    assign weights1[16][69] = 16'b1111111110101100;
    assign weights1[16][70] = 16'b1111111110101001;
    assign weights1[16][71] = 16'b1111111110001111;
    assign weights1[16][72] = 16'b1111111110100111;
    assign weights1[16][73] = 16'b1111111110101001;
    assign weights1[16][74] = 16'b1111111110101101;
    assign weights1[16][75] = 16'b1111111110101100;
    assign weights1[16][76] = 16'b1111111111000101;
    assign weights1[16][77] = 16'b1111111111010010;
    assign weights1[16][78] = 16'b1111111111010100;
    assign weights1[16][79] = 16'b1111111111011000;
    assign weights1[16][80] = 16'b1111111111100011;
    assign weights1[16][81] = 16'b1111111111110000;
    assign weights1[16][82] = 16'b1111111111111100;
    assign weights1[16][83] = 16'b1111111111110111;
    assign weights1[16][84] = 16'b0000000000000001;
    assign weights1[16][85] = 16'b1111111111111001;
    assign weights1[16][86] = 16'b1111111111110010;
    assign weights1[16][87] = 16'b1111111111100100;
    assign weights1[16][88] = 16'b1111111111100010;
    assign weights1[16][89] = 16'b1111111111010101;
    assign weights1[16][90] = 16'b1111111111000110;
    assign weights1[16][91] = 16'b1111111110110110;
    assign weights1[16][92] = 16'b1111111111000110;
    assign weights1[16][93] = 16'b1111111110101101;
    assign weights1[16][94] = 16'b1111111110011110;
    assign weights1[16][95] = 16'b1111111110100000;
    assign weights1[16][96] = 16'b1111111110001010;
    assign weights1[16][97] = 16'b1111111101110001;
    assign weights1[16][98] = 16'b1111111110011111;
    assign weights1[16][99] = 16'b1111111110011010;
    assign weights1[16][100] = 16'b1111111110111110;
    assign weights1[16][101] = 16'b1111111111000001;
    assign weights1[16][102] = 16'b1111111110101001;
    assign weights1[16][103] = 16'b1111111111000111;
    assign weights1[16][104] = 16'b1111111111000011;
    assign weights1[16][105] = 16'b1111111111010101;
    assign weights1[16][106] = 16'b1111111111011010;
    assign weights1[16][107] = 16'b1111111111001011;
    assign weights1[16][108] = 16'b1111111111100001;
    assign weights1[16][109] = 16'b1111111111100111;
    assign weights1[16][110] = 16'b1111111111110010;
    assign weights1[16][111] = 16'b1111111111110101;
    assign weights1[16][112] = 16'b0000000000000001;
    assign weights1[16][113] = 16'b1111111111111001;
    assign weights1[16][114] = 16'b1111111111110010;
    assign weights1[16][115] = 16'b1111111111100011;
    assign weights1[16][116] = 16'b1111111111011111;
    assign weights1[16][117] = 16'b1111111111001011;
    assign weights1[16][118] = 16'b1111111111010111;
    assign weights1[16][119] = 16'b1111111111001101;
    assign weights1[16][120] = 16'b1111111111001010;
    assign weights1[16][121] = 16'b1111111111100100;
    assign weights1[16][122] = 16'b1111111111010110;
    assign weights1[16][123] = 16'b1111111111100001;
    assign weights1[16][124] = 16'b1111111111100101;
    assign weights1[16][125] = 16'b1111111111011010;
    assign weights1[16][126] = 16'b1111111111011101;
    assign weights1[16][127] = 16'b1111111111111001;
    assign weights1[16][128] = 16'b1111111111110000;
    assign weights1[16][129] = 16'b1111111111101100;
    assign weights1[16][130] = 16'b1111111111101100;
    assign weights1[16][131] = 16'b1111111111100011;
    assign weights1[16][132] = 16'b0000000000000001;
    assign weights1[16][133] = 16'b1111111111011110;
    assign weights1[16][134] = 16'b1111111111101100;
    assign weights1[16][135] = 16'b1111111111101011;
    assign weights1[16][136] = 16'b1111111111010110;
    assign weights1[16][137] = 16'b1111111111001011;
    assign weights1[16][138] = 16'b1111111111101001;
    assign weights1[16][139] = 16'b1111111111110001;
    assign weights1[16][140] = 16'b0000000000000101;
    assign weights1[16][141] = 16'b1111111111111111;
    assign weights1[16][142] = 16'b1111111111110001;
    assign weights1[16][143] = 16'b1111111111110001;
    assign weights1[16][144] = 16'b1111111111111000;
    assign weights1[16][145] = 16'b1111111111111000;
    assign weights1[16][146] = 16'b0000000000000101;
    assign weights1[16][147] = 16'b0000000000001001;
    assign weights1[16][148] = 16'b0000000000010101;
    assign weights1[16][149] = 16'b0000000000001110;
    assign weights1[16][150] = 16'b0000000000000101;
    assign weights1[16][151] = 16'b0000000000110110;
    assign weights1[16][152] = 16'b0000000000111010;
    assign weights1[16][153] = 16'b0000000000011100;
    assign weights1[16][154] = 16'b0000000000011100;
    assign weights1[16][155] = 16'b0000000000100100;
    assign weights1[16][156] = 16'b0000000000001111;
    assign weights1[16][157] = 16'b0000000000000101;
    assign weights1[16][158] = 16'b0000000000000010;
    assign weights1[16][159] = 16'b0000000000000110;
    assign weights1[16][160] = 16'b1111111111110010;
    assign weights1[16][161] = 16'b1111111111110110;
    assign weights1[16][162] = 16'b1111111111110100;
    assign weights1[16][163] = 16'b1111111111110110;
    assign weights1[16][164] = 16'b1111111111101001;
    assign weights1[16][165] = 16'b1111111111000101;
    assign weights1[16][166] = 16'b1111111111010110;
    assign weights1[16][167] = 16'b1111111111100010;
    assign weights1[16][168] = 16'b0000000000000100;
    assign weights1[16][169] = 16'b0000000000000100;
    assign weights1[16][170] = 16'b0000000000000010;
    assign weights1[16][171] = 16'b0000000000010000;
    assign weights1[16][172] = 16'b0000000000011101;
    assign weights1[16][173] = 16'b0000000000110010;
    assign weights1[16][174] = 16'b0000000001000010;
    assign weights1[16][175] = 16'b0000000001010010;
    assign weights1[16][176] = 16'b0000000001010100;
    assign weights1[16][177] = 16'b0000000001001001;
    assign weights1[16][178] = 16'b0000000000110100;
    assign weights1[16][179] = 16'b0000000000101000;
    assign weights1[16][180] = 16'b0000000000011101;
    assign weights1[16][181] = 16'b0000000000111101;
    assign weights1[16][182] = 16'b0000000000101100;
    assign weights1[16][183] = 16'b0000000000101100;
    assign weights1[16][184] = 16'b0000000000001111;
    assign weights1[16][185] = 16'b0000000000010000;
    assign weights1[16][186] = 16'b0000000000101000;
    assign weights1[16][187] = 16'b0000000000011011;
    assign weights1[16][188] = 16'b0000000000000000;
    assign weights1[16][189] = 16'b0000000000010001;
    assign weights1[16][190] = 16'b0000000000010101;
    assign weights1[16][191] = 16'b1111111111110011;
    assign weights1[16][192] = 16'b1111111111101111;
    assign weights1[16][193] = 16'b1111111111101101;
    assign weights1[16][194] = 16'b1111111111101001;
    assign weights1[16][195] = 16'b1111111111100100;
    assign weights1[16][196] = 16'b0000000000000111;
    assign weights1[16][197] = 16'b0000000000010101;
    assign weights1[16][198] = 16'b0000000000100100;
    assign weights1[16][199] = 16'b0000000000101010;
    assign weights1[16][200] = 16'b0000000001000101;
    assign weights1[16][201] = 16'b0000000000111100;
    assign weights1[16][202] = 16'b0000000001000010;
    assign weights1[16][203] = 16'b0000000001001100;
    assign weights1[16][204] = 16'b0000000000100110;
    assign weights1[16][205] = 16'b0000000000100100;
    assign weights1[16][206] = 16'b0000000001001000;
    assign weights1[16][207] = 16'b0000000000111100;
    assign weights1[16][208] = 16'b0000000000111000;
    assign weights1[16][209] = 16'b0000000000101011;
    assign weights1[16][210] = 16'b0000000000100010;
    assign weights1[16][211] = 16'b0000000000001110;
    assign weights1[16][212] = 16'b0000000000011110;
    assign weights1[16][213] = 16'b0000000000100001;
    assign weights1[16][214] = 16'b0000000000011001;
    assign weights1[16][215] = 16'b1111111111111101;
    assign weights1[16][216] = 16'b0000000000011101;
    assign weights1[16][217] = 16'b0000000000001110;
    assign weights1[16][218] = 16'b0000000000100100;
    assign weights1[16][219] = 16'b0000000000001110;
    assign weights1[16][220] = 16'b0000000000000101;
    assign weights1[16][221] = 16'b0000000000000010;
    assign weights1[16][222] = 16'b1111111111100001;
    assign weights1[16][223] = 16'b1111111111100101;
    assign weights1[16][224] = 16'b0000000000010011;
    assign weights1[16][225] = 16'b0000000000011110;
    assign weights1[16][226] = 16'b0000000000101000;
    assign weights1[16][227] = 16'b0000000000101111;
    assign weights1[16][228] = 16'b0000000000110111;
    assign weights1[16][229] = 16'b0000000000101111;
    assign weights1[16][230] = 16'b0000000000110101;
    assign weights1[16][231] = 16'b0000000000001101;
    assign weights1[16][232] = 16'b0000000000100110;
    assign weights1[16][233] = 16'b0000000000110110;
    assign weights1[16][234] = 16'b0000000000111001;
    assign weights1[16][235] = 16'b0000000000101110;
    assign weights1[16][236] = 16'b0000000001001001;
    assign weights1[16][237] = 16'b0000000000110011;
    assign weights1[16][238] = 16'b0000000001001101;
    assign weights1[16][239] = 16'b0000000000111000;
    assign weights1[16][240] = 16'b0000000001010110;
    assign weights1[16][241] = 16'b0000000000100110;
    assign weights1[16][242] = 16'b0000000000110110;
    assign weights1[16][243] = 16'b0000000000011011;
    assign weights1[16][244] = 16'b0000000000010111;
    assign weights1[16][245] = 16'b1111111111111111;
    assign weights1[16][246] = 16'b0000000000000111;
    assign weights1[16][247] = 16'b1111111111111110;
    assign weights1[16][248] = 16'b0000000000001111;
    assign weights1[16][249] = 16'b1111111111110100;
    assign weights1[16][250] = 16'b1111111111101010;
    assign weights1[16][251] = 16'b1111111111101001;
    assign weights1[16][252] = 16'b0000000000010001;
    assign weights1[16][253] = 16'b0000000000011010;
    assign weights1[16][254] = 16'b0000000000010001;
    assign weights1[16][255] = 16'b0000000000100100;
    assign weights1[16][256] = 16'b0000000000001011;
    assign weights1[16][257] = 16'b0000000000010100;
    assign weights1[16][258] = 16'b0000000000010101;
    assign weights1[16][259] = 16'b1111111111110000;
    assign weights1[16][260] = 16'b1111111111100101;
    assign weights1[16][261] = 16'b1111111111100100;
    assign weights1[16][262] = 16'b1111111111111100;
    assign weights1[16][263] = 16'b1111111111101001;
    assign weights1[16][264] = 16'b0000000000000001;
    assign weights1[16][265] = 16'b0000000000010100;
    assign weights1[16][266] = 16'b0000000000001101;
    assign weights1[16][267] = 16'b0000000000011110;
    assign weights1[16][268] = 16'b0000000000011111;
    assign weights1[16][269] = 16'b0000000000100010;
    assign weights1[16][270] = 16'b0000000000101000;
    assign weights1[16][271] = 16'b0000000000000111;
    assign weights1[16][272] = 16'b0000000000101001;
    assign weights1[16][273] = 16'b0000000000010000;
    assign weights1[16][274] = 16'b0000000000001010;
    assign weights1[16][275] = 16'b0000000000011100;
    assign weights1[16][276] = 16'b1111111111111110;
    assign weights1[16][277] = 16'b0000000000010010;
    assign weights1[16][278] = 16'b0000000000000111;
    assign weights1[16][279] = 16'b1111111111101100;
    assign weights1[16][280] = 16'b0000000000001101;
    assign weights1[16][281] = 16'b0000000000000000;
    assign weights1[16][282] = 16'b1111111111111011;
    assign weights1[16][283] = 16'b1111111111111011;
    assign weights1[16][284] = 16'b1111111111100001;
    assign weights1[16][285] = 16'b1111111111111011;
    assign weights1[16][286] = 16'b1111111111110001;
    assign weights1[16][287] = 16'b1111111111110000;
    assign weights1[16][288] = 16'b1111111111011000;
    assign weights1[16][289] = 16'b1111111111011101;
    assign weights1[16][290] = 16'b1111111111010100;
    assign weights1[16][291] = 16'b1111111111000101;
    assign weights1[16][292] = 16'b1111111111011111;
    assign weights1[16][293] = 16'b1111111111000011;
    assign weights1[16][294] = 16'b1111111111011010;
    assign weights1[16][295] = 16'b1111111111100100;
    assign weights1[16][296] = 16'b0000000000011000;
    assign weights1[16][297] = 16'b1111111111110101;
    assign weights1[16][298] = 16'b0000000000101011;
    assign weights1[16][299] = 16'b0000000000100011;
    assign weights1[16][300] = 16'b0000000000100100;
    assign weights1[16][301] = 16'b0000000000100101;
    assign weights1[16][302] = 16'b0000000000100100;
    assign weights1[16][303] = 16'b0000000000011101;
    assign weights1[16][304] = 16'b0000000000010011;
    assign weights1[16][305] = 16'b0000000000100000;
    assign weights1[16][306] = 16'b0000000000000100;
    assign weights1[16][307] = 16'b0000000000000100;
    assign weights1[16][308] = 16'b0000000000000000;
    assign weights1[16][309] = 16'b1111111111111000;
    assign weights1[16][310] = 16'b1111111111110000;
    assign weights1[16][311] = 16'b1111111111010010;
    assign weights1[16][312] = 16'b1111111111001101;
    assign weights1[16][313] = 16'b1111111111100101;
    assign weights1[16][314] = 16'b1111111111000000;
    assign weights1[16][315] = 16'b1111111111000111;
    assign weights1[16][316] = 16'b1111111111100110;
    assign weights1[16][317] = 16'b1111111111010001;
    assign weights1[16][318] = 16'b1111111111011001;
    assign weights1[16][319] = 16'b1111111111011010;
    assign weights1[16][320] = 16'b1111111111010101;
    assign weights1[16][321] = 16'b1111111111100000;
    assign weights1[16][322] = 16'b1111111111011000;
    assign weights1[16][323] = 16'b1111111111000011;
    assign weights1[16][324] = 16'b1111111111100100;
    assign weights1[16][325] = 16'b0000000000000001;
    assign weights1[16][326] = 16'b0000000000001000;
    assign weights1[16][327] = 16'b0000000000000111;
    assign weights1[16][328] = 16'b0000000000010111;
    assign weights1[16][329] = 16'b0000000000010001;
    assign weights1[16][330] = 16'b0000000000101011;
    assign weights1[16][331] = 16'b0000000000101001;
    assign weights1[16][332] = 16'b0000000000010100;
    assign weights1[16][333] = 16'b0000000000010101;
    assign weights1[16][334] = 16'b0000000000010011;
    assign weights1[16][335] = 16'b0000000000000100;
    assign weights1[16][336] = 16'b1111111111110110;
    assign weights1[16][337] = 16'b1111111111100111;
    assign weights1[16][338] = 16'b1111111111101001;
    assign weights1[16][339] = 16'b1111111111011100;
    assign weights1[16][340] = 16'b1111111111011000;
    assign weights1[16][341] = 16'b1111111111000111;
    assign weights1[16][342] = 16'b1111111110110110;
    assign weights1[16][343] = 16'b1111111111101100;
    assign weights1[16][344] = 16'b1111111111101111;
    assign weights1[16][345] = 16'b0000000000000011;
    assign weights1[16][346] = 16'b1111111111101100;
    assign weights1[16][347] = 16'b1111111111110010;
    assign weights1[16][348] = 16'b1111111111101000;
    assign weights1[16][349] = 16'b1111111111011001;
    assign weights1[16][350] = 16'b1111111111010111;
    assign weights1[16][351] = 16'b1111111111101010;
    assign weights1[16][352] = 16'b1111111111100000;
    assign weights1[16][353] = 16'b1111111111110010;
    assign weights1[16][354] = 16'b0000000000001111;
    assign weights1[16][355] = 16'b0000000000001011;
    assign weights1[16][356] = 16'b0000000000000010;
    assign weights1[16][357] = 16'b0000000000001101;
    assign weights1[16][358] = 16'b0000000000001011;
    assign weights1[16][359] = 16'b0000000000000001;
    assign weights1[16][360] = 16'b1111111111110010;
    assign weights1[16][361] = 16'b0000000000011101;
    assign weights1[16][362] = 16'b0000000000001000;
    assign weights1[16][363] = 16'b0000000000000110;
    assign weights1[16][364] = 16'b1111111111101000;
    assign weights1[16][365] = 16'b1111111111011111;
    assign weights1[16][366] = 16'b1111111111011111;
    assign weights1[16][367] = 16'b1111111111011101;
    assign weights1[16][368] = 16'b1111111111011101;
    assign weights1[16][369] = 16'b1111111111011000;
    assign weights1[16][370] = 16'b1111111111000010;
    assign weights1[16][371] = 16'b1111111111101110;
    assign weights1[16][372] = 16'b0000000000001001;
    assign weights1[16][373] = 16'b1111111111111101;
    assign weights1[16][374] = 16'b1111111111111110;
    assign weights1[16][375] = 16'b0000000000000101;
    assign weights1[16][376] = 16'b0000000000001000;
    assign weights1[16][377] = 16'b1111111111111001;
    assign weights1[16][378] = 16'b1111111111100011;
    assign weights1[16][379] = 16'b0000000000000001;
    assign weights1[16][380] = 16'b0000000000001010;
    assign weights1[16][381] = 16'b1111111111101100;
    assign weights1[16][382] = 16'b0000000000000100;
    assign weights1[16][383] = 16'b0000000000000001;
    assign weights1[16][384] = 16'b0000000000010001;
    assign weights1[16][385] = 16'b0000000000011001;
    assign weights1[16][386] = 16'b0000000000000001;
    assign weights1[16][387] = 16'b0000000000001111;
    assign weights1[16][388] = 16'b0000000000000101;
    assign weights1[16][389] = 16'b0000000000001011;
    assign weights1[16][390] = 16'b0000000000001001;
    assign weights1[16][391] = 16'b0000000000001100;
    assign weights1[16][392] = 16'b1111111111100110;
    assign weights1[16][393] = 16'b1111111111011100;
    assign weights1[16][394] = 16'b1111111111101000;
    assign weights1[16][395] = 16'b1111111111100010;
    assign weights1[16][396] = 16'b0000000000000111;
    assign weights1[16][397] = 16'b1111111111011011;
    assign weights1[16][398] = 16'b1111111111011010;
    assign weights1[16][399] = 16'b1111111111111110;
    assign weights1[16][400] = 16'b1111111111110010;
    assign weights1[16][401] = 16'b1111111111100101;
    assign weights1[16][402] = 16'b1111111111111001;
    assign weights1[16][403] = 16'b0000000000000010;
    assign weights1[16][404] = 16'b1111111111111101;
    assign weights1[16][405] = 16'b0000000000001010;
    assign weights1[16][406] = 16'b0000000000000100;
    assign weights1[16][407] = 16'b1111111111110100;
    assign weights1[16][408] = 16'b1111111111100100;
    assign weights1[16][409] = 16'b1111111111101110;
    assign weights1[16][410] = 16'b1111111111100111;
    assign weights1[16][411] = 16'b1111111111111001;
    assign weights1[16][412] = 16'b1111111111110111;
    assign weights1[16][413] = 16'b0000000000001000;
    assign weights1[16][414] = 16'b0000000000011001;
    assign weights1[16][415] = 16'b1111111111111101;
    assign weights1[16][416] = 16'b0000000000011110;
    assign weights1[16][417] = 16'b0000000000000110;
    assign weights1[16][418] = 16'b0000000000001000;
    assign weights1[16][419] = 16'b0000000000001011;
    assign weights1[16][420] = 16'b1111111111110100;
    assign weights1[16][421] = 16'b1111111111101001;
    assign weights1[16][422] = 16'b1111111111100010;
    assign weights1[16][423] = 16'b1111111111101001;
    assign weights1[16][424] = 16'b0000000000001000;
    assign weights1[16][425] = 16'b0000000000000010;
    assign weights1[16][426] = 16'b0000000000001100;
    assign weights1[16][427] = 16'b1111111111101010;
    assign weights1[16][428] = 16'b1111111111110000;
    assign weights1[16][429] = 16'b1111111111111000;
    assign weights1[16][430] = 16'b0000000000001000;
    assign weights1[16][431] = 16'b1111111111110001;
    assign weights1[16][432] = 16'b0000000000000110;
    assign weights1[16][433] = 16'b1111111111111110;
    assign weights1[16][434] = 16'b0000000000001000;
    assign weights1[16][435] = 16'b1111111111110100;
    assign weights1[16][436] = 16'b1111111111110010;
    assign weights1[16][437] = 16'b0000000000000101;
    assign weights1[16][438] = 16'b1111111111111001;
    assign weights1[16][439] = 16'b1111111111011111;
    assign weights1[16][440] = 16'b1111111111111000;
    assign weights1[16][441] = 16'b1111111111111010;
    assign weights1[16][442] = 16'b0000000000011010;
    assign weights1[16][443] = 16'b0000000000000100;
    assign weights1[16][444] = 16'b0000000000000110;
    assign weights1[16][445] = 16'b1111111111110111;
    assign weights1[16][446] = 16'b1111111111110100;
    assign weights1[16][447] = 16'b0000000000000110;
    assign weights1[16][448] = 16'b1111111111111010;
    assign weights1[16][449] = 16'b1111111111111101;
    assign weights1[16][450] = 16'b1111111111111000;
    assign weights1[16][451] = 16'b1111111111111010;
    assign weights1[16][452] = 16'b1111111111111010;
    assign weights1[16][453] = 16'b0000000000010010;
    assign weights1[16][454] = 16'b1111111111110110;
    assign weights1[16][455] = 16'b1111111111111001;
    assign weights1[16][456] = 16'b0000000000000011;
    assign weights1[16][457] = 16'b1111111111111100;
    assign weights1[16][458] = 16'b0000000000010010;
    assign weights1[16][459] = 16'b0000000000010111;
    assign weights1[16][460] = 16'b1111111111111001;
    assign weights1[16][461] = 16'b0000000000000001;
    assign weights1[16][462] = 16'b1111111111110110;
    assign weights1[16][463] = 16'b0000000000000100;
    assign weights1[16][464] = 16'b0000000000001000;
    assign weights1[16][465] = 16'b1111111111101100;
    assign weights1[16][466] = 16'b1111111111101000;
    assign weights1[16][467] = 16'b1111111111011000;
    assign weights1[16][468] = 16'b0000000000000101;
    assign weights1[16][469] = 16'b1111111111111110;
    assign weights1[16][470] = 16'b0000000000000011;
    assign weights1[16][471] = 16'b0000000000001111;
    assign weights1[16][472] = 16'b0000000000001011;
    assign weights1[16][473] = 16'b0000000000000011;
    assign weights1[16][474] = 16'b0000000000000000;
    assign weights1[16][475] = 16'b0000000000000001;
    assign weights1[16][476] = 16'b1111111111110110;
    assign weights1[16][477] = 16'b0000000000000010;
    assign weights1[16][478] = 16'b1111111111111100;
    assign weights1[16][479] = 16'b1111111111111101;
    assign weights1[16][480] = 16'b0000000000011101;
    assign weights1[16][481] = 16'b0000000000010010;
    assign weights1[16][482] = 16'b0000000000000111;
    assign weights1[16][483] = 16'b1111111111111100;
    assign weights1[16][484] = 16'b0000000000001000;
    assign weights1[16][485] = 16'b0000000000000011;
    assign weights1[16][486] = 16'b1111111111100100;
    assign weights1[16][487] = 16'b0000000000000001;
    assign weights1[16][488] = 16'b0000000000000010;
    assign weights1[16][489] = 16'b1111111111100110;
    assign weights1[16][490] = 16'b1111111111101110;
    assign weights1[16][491] = 16'b1111111111111101;
    assign weights1[16][492] = 16'b0000000000000000;
    assign weights1[16][493] = 16'b1111111111111100;
    assign weights1[16][494] = 16'b1111111111110111;
    assign weights1[16][495] = 16'b1111111111110010;
    assign weights1[16][496] = 16'b1111111111101110;
    assign weights1[16][497] = 16'b1111111111110001;
    assign weights1[16][498] = 16'b1111111111110000;
    assign weights1[16][499] = 16'b0000000000001001;
    assign weights1[16][500] = 16'b0000000000000000;
    assign weights1[16][501] = 16'b1111111111111011;
    assign weights1[16][502] = 16'b1111111111111101;
    assign weights1[16][503] = 16'b0000000000000111;
    assign weights1[16][504] = 16'b1111111111110111;
    assign weights1[16][505] = 16'b0000000000000001;
    assign weights1[16][506] = 16'b0000000000001000;
    assign weights1[16][507] = 16'b1111111111111001;
    assign weights1[16][508] = 16'b0000000000001110;
    assign weights1[16][509] = 16'b0000000000010011;
    assign weights1[16][510] = 16'b0000000000010000;
    assign weights1[16][511] = 16'b1111111111110110;
    assign weights1[16][512] = 16'b0000000000001111;
    assign weights1[16][513] = 16'b0000000000000110;
    assign weights1[16][514] = 16'b0000000000000100;
    assign weights1[16][515] = 16'b1111111111111010;
    assign weights1[16][516] = 16'b0000000000000101;
    assign weights1[16][517] = 16'b0000000000001001;
    assign weights1[16][518] = 16'b1111111111100101;
    assign weights1[16][519] = 16'b1111111111110000;
    assign weights1[16][520] = 16'b0000000000001001;
    assign weights1[16][521] = 16'b0000000000010000;
    assign weights1[16][522] = 16'b0000000000010111;
    assign weights1[16][523] = 16'b0000000000001000;
    assign weights1[16][524] = 16'b1111111111110110;
    assign weights1[16][525] = 16'b1111111111101011;
    assign weights1[16][526] = 16'b0000000000001100;
    assign weights1[16][527] = 16'b0000000000000011;
    assign weights1[16][528] = 16'b0000000000000111;
    assign weights1[16][529] = 16'b1111111111111000;
    assign weights1[16][530] = 16'b1111111111111011;
    assign weights1[16][531] = 16'b0000000000001111;
    assign weights1[16][532] = 16'b1111111111111011;
    assign weights1[16][533] = 16'b1111111111110101;
    assign weights1[16][534] = 16'b0000000000000111;
    assign weights1[16][535] = 16'b1111111111111101;
    assign weights1[16][536] = 16'b1111111111111100;
    assign weights1[16][537] = 16'b0000000000000110;
    assign weights1[16][538] = 16'b1111111111111001;
    assign weights1[16][539] = 16'b1111111111111110;
    assign weights1[16][540] = 16'b0000000000010010;
    assign weights1[16][541] = 16'b0000000000000100;
    assign weights1[16][542] = 16'b0000000000000100;
    assign weights1[16][543] = 16'b1111111111110010;
    assign weights1[16][544] = 16'b0000000000011010;
    assign weights1[16][545] = 16'b1111111111101011;
    assign weights1[16][546] = 16'b1111111111111110;
    assign weights1[16][547] = 16'b0000000000000100;
    assign weights1[16][548] = 16'b1111111111101110;
    assign weights1[16][549] = 16'b1111111111111101;
    assign weights1[16][550] = 16'b1111111111110000;
    assign weights1[16][551] = 16'b0000000000001111;
    assign weights1[16][552] = 16'b0000000000001100;
    assign weights1[16][553] = 16'b0000000000000111;
    assign weights1[16][554] = 16'b0000000000000010;
    assign weights1[16][555] = 16'b0000000000011111;
    assign weights1[16][556] = 16'b0000000000001010;
    assign weights1[16][557] = 16'b0000000000000010;
    assign weights1[16][558] = 16'b0000000000000001;
    assign weights1[16][559] = 16'b1111111111110110;
    assign weights1[16][560] = 16'b0000000000000110;
    assign weights1[16][561] = 16'b0000000000001100;
    assign weights1[16][562] = 16'b1111111111111001;
    assign weights1[16][563] = 16'b1111111111111111;
    assign weights1[16][564] = 16'b0000000000010000;
    assign weights1[16][565] = 16'b1111111111111110;
    assign weights1[16][566] = 16'b1111111111111111;
    assign weights1[16][567] = 16'b0000000000011101;
    assign weights1[16][568] = 16'b0000000000001001;
    assign weights1[16][569] = 16'b1111111111110111;
    assign weights1[16][570] = 16'b0000000000001000;
    assign weights1[16][571] = 16'b1111111111110111;
    assign weights1[16][572] = 16'b1111111111111011;
    assign weights1[16][573] = 16'b1111111111100111;
    assign weights1[16][574] = 16'b0000000000000110;
    assign weights1[16][575] = 16'b1111111111110110;
    assign weights1[16][576] = 16'b1111111111111110;
    assign weights1[16][577] = 16'b1111111111110000;
    assign weights1[16][578] = 16'b0000000000000001;
    assign weights1[16][579] = 16'b0000000000000101;
    assign weights1[16][580] = 16'b1111111111111010;
    assign weights1[16][581] = 16'b0000000000011101;
    assign weights1[16][582] = 16'b1111111111101001;
    assign weights1[16][583] = 16'b0000000000000100;
    assign weights1[16][584] = 16'b0000000000000111;
    assign weights1[16][585] = 16'b0000000000000100;
    assign weights1[16][586] = 16'b1111111111110111;
    assign weights1[16][587] = 16'b1111111111111011;
    assign weights1[16][588] = 16'b1111111111111110;
    assign weights1[16][589] = 16'b1111111111111110;
    assign weights1[16][590] = 16'b1111111111111001;
    assign weights1[16][591] = 16'b1111111111100011;
    assign weights1[16][592] = 16'b0000000000001101;
    assign weights1[16][593] = 16'b0000000000001111;
    assign weights1[16][594] = 16'b0000000000000101;
    assign weights1[16][595] = 16'b1111111111110111;
    assign weights1[16][596] = 16'b1111111111110101;
    assign weights1[16][597] = 16'b0000000000001111;
    assign weights1[16][598] = 16'b1111111111111111;
    assign weights1[16][599] = 16'b0000000000010010;
    assign weights1[16][600] = 16'b0000000000001100;
    assign weights1[16][601] = 16'b0000000000000000;
    assign weights1[16][602] = 16'b1111111111111110;
    assign weights1[16][603] = 16'b0000000000010111;
    assign weights1[16][604] = 16'b1111111111111001;
    assign weights1[16][605] = 16'b0000000000001000;
    assign weights1[16][606] = 16'b0000000000000010;
    assign weights1[16][607] = 16'b0000000000001000;
    assign weights1[16][608] = 16'b1111111111101011;
    assign weights1[16][609] = 16'b1111111111111000;
    assign weights1[16][610] = 16'b1111111111110111;
    assign weights1[16][611] = 16'b1111111111111001;
    assign weights1[16][612] = 16'b1111111111110100;
    assign weights1[16][613] = 16'b1111111111111100;
    assign weights1[16][614] = 16'b1111111111111101;
    assign weights1[16][615] = 16'b0000000000000010;
    assign weights1[16][616] = 16'b0000000000000010;
    assign weights1[16][617] = 16'b1111111111111111;
    assign weights1[16][618] = 16'b1111111111111111;
    assign weights1[16][619] = 16'b0000000000000100;
    assign weights1[16][620] = 16'b1111111111110011;
    assign weights1[16][621] = 16'b1111111111101111;
    assign weights1[16][622] = 16'b1111111111101000;
    assign weights1[16][623] = 16'b0000000000000000;
    assign weights1[16][624] = 16'b0000000000000010;
    assign weights1[16][625] = 16'b0000000000010100;
    assign weights1[16][626] = 16'b1111111111110111;
    assign weights1[16][627] = 16'b1111111111101000;
    assign weights1[16][628] = 16'b0000000000000010;
    assign weights1[16][629] = 16'b0000000000010111;
    assign weights1[16][630] = 16'b1111111111110110;
    assign weights1[16][631] = 16'b0000000000000001;
    assign weights1[16][632] = 16'b1111111111111111;
    assign weights1[16][633] = 16'b1111111111110101;
    assign weights1[16][634] = 16'b0000000000000111;
    assign weights1[16][635] = 16'b0000000000010101;
    assign weights1[16][636] = 16'b1111111111111001;
    assign weights1[16][637] = 16'b1111111111111010;
    assign weights1[16][638] = 16'b0000000000001000;
    assign weights1[16][639] = 16'b0000000000000100;
    assign weights1[16][640] = 16'b1111111111111111;
    assign weights1[16][641] = 16'b1111111111111001;
    assign weights1[16][642] = 16'b1111111111111010;
    assign weights1[16][643] = 16'b1111111111111100;
    assign weights1[16][644] = 16'b1111111111111011;
    assign weights1[16][645] = 16'b1111111111111111;
    assign weights1[16][646] = 16'b1111111111110111;
    assign weights1[16][647] = 16'b0000000000000000;
    assign weights1[16][648] = 16'b0000000000001001;
    assign weights1[16][649] = 16'b1111111111100111;
    assign weights1[16][650] = 16'b1111111111111101;
    assign weights1[16][651] = 16'b0000000000001001;
    assign weights1[16][652] = 16'b1111111111110010;
    assign weights1[16][653] = 16'b1111111111111010;
    assign weights1[16][654] = 16'b0000000000000000;
    assign weights1[16][655] = 16'b0000000000010001;
    assign weights1[16][656] = 16'b0000000000010111;
    assign weights1[16][657] = 16'b0000000000000010;
    assign weights1[16][658] = 16'b1111111111101110;
    assign weights1[16][659] = 16'b1111111111100011;
    assign weights1[16][660] = 16'b0000000000000110;
    assign weights1[16][661] = 16'b1111111111100010;
    assign weights1[16][662] = 16'b1111111111110111;
    assign weights1[16][663] = 16'b1111111111110011;
    assign weights1[16][664] = 16'b1111111111100111;
    assign weights1[16][665] = 16'b1111111111110111;
    assign weights1[16][666] = 16'b1111111111111001;
    assign weights1[16][667] = 16'b0000000000001111;
    assign weights1[16][668] = 16'b1111111111111101;
    assign weights1[16][669] = 16'b1111111111111000;
    assign weights1[16][670] = 16'b1111111111101110;
    assign weights1[16][671] = 16'b1111111111111111;
    assign weights1[16][672] = 16'b1111111111111011;
    assign weights1[16][673] = 16'b1111111111111111;
    assign weights1[16][674] = 16'b0000000000000101;
    assign weights1[16][675] = 16'b1111111111111100;
    assign weights1[16][676] = 16'b0000000000000010;
    assign weights1[16][677] = 16'b0000000000001011;
    assign weights1[16][678] = 16'b1111111111101011;
    assign weights1[16][679] = 16'b1111111111101010;
    assign weights1[16][680] = 16'b1111111111100110;
    assign weights1[16][681] = 16'b1111111111110111;
    assign weights1[16][682] = 16'b1111111111110111;
    assign weights1[16][683] = 16'b1111111111110110;
    assign weights1[16][684] = 16'b1111111111111011;
    assign weights1[16][685] = 16'b0000000000011100;
    assign weights1[16][686] = 16'b1111111111111101;
    assign weights1[16][687] = 16'b0000000000000010;
    assign weights1[16][688] = 16'b0000000000011000;
    assign weights1[16][689] = 16'b1111111111101100;
    assign weights1[16][690] = 16'b0000000000001101;
    assign weights1[16][691] = 16'b1111111111111100;
    assign weights1[16][692] = 16'b1111111111111110;
    assign weights1[16][693] = 16'b1111111111110110;
    assign weights1[16][694] = 16'b1111111111101001;
    assign weights1[16][695] = 16'b1111111111111011;
    assign weights1[16][696] = 16'b1111111111110101;
    assign weights1[16][697] = 16'b1111111111111010;
    assign weights1[16][698] = 16'b1111111111111010;
    assign weights1[16][699] = 16'b0000000000000010;
    assign weights1[16][700] = 16'b1111111111111000;
    assign weights1[16][701] = 16'b1111111111111000;
    assign weights1[16][702] = 16'b1111111111111100;
    assign weights1[16][703] = 16'b0000000000000000;
    assign weights1[16][704] = 16'b0000000000000100;
    assign weights1[16][705] = 16'b1111111111111110;
    assign weights1[16][706] = 16'b0000000000000011;
    assign weights1[16][707] = 16'b0000000000001001;
    assign weights1[16][708] = 16'b0000000000000011;
    assign weights1[16][709] = 16'b0000000000001110;
    assign weights1[16][710] = 16'b0000000000000010;
    assign weights1[16][711] = 16'b0000000000000101;
    assign weights1[16][712] = 16'b0000000000000000;
    assign weights1[16][713] = 16'b1111111111101110;
    assign weights1[16][714] = 16'b1111111111111010;
    assign weights1[16][715] = 16'b0000000000100011;
    assign weights1[16][716] = 16'b1111111111111110;
    assign weights1[16][717] = 16'b1111111111111010;
    assign weights1[16][718] = 16'b0000000000000000;
    assign weights1[16][719] = 16'b1111111111110000;
    assign weights1[16][720] = 16'b1111111111111110;
    assign weights1[16][721] = 16'b1111111111110000;
    assign weights1[16][722] = 16'b1111111111110000;
    assign weights1[16][723] = 16'b1111111111101100;
    assign weights1[16][724] = 16'b1111111111101101;
    assign weights1[16][725] = 16'b1111111111111001;
    assign weights1[16][726] = 16'b1111111111111100;
    assign weights1[16][727] = 16'b0000000000000101;
    assign weights1[16][728] = 16'b1111111111111111;
    assign weights1[16][729] = 16'b1111111111111101;
    assign weights1[16][730] = 16'b1111111111111100;
    assign weights1[16][731] = 16'b1111111111111101;
    assign weights1[16][732] = 16'b0000000000000100;
    assign weights1[16][733] = 16'b1111111111111000;
    assign weights1[16][734] = 16'b1111111111110110;
    assign weights1[16][735] = 16'b0000000000000010;
    assign weights1[16][736] = 16'b1111111111111111;
    assign weights1[16][737] = 16'b1111111111111101;
    assign weights1[16][738] = 16'b1111111111110100;
    assign weights1[16][739] = 16'b1111111111101010;
    assign weights1[16][740] = 16'b1111111111110011;
    assign weights1[16][741] = 16'b1111111111101110;
    assign weights1[16][742] = 16'b1111111111111101;
    assign weights1[16][743] = 16'b1111111111110110;
    assign weights1[16][744] = 16'b1111111111100010;
    assign weights1[16][745] = 16'b1111111111110101;
    assign weights1[16][746] = 16'b1111111111101110;
    assign weights1[16][747] = 16'b1111111111111100;
    assign weights1[16][748] = 16'b1111111111111000;
    assign weights1[16][749] = 16'b1111111111111010;
    assign weights1[16][750] = 16'b1111111111110110;
    assign weights1[16][751] = 16'b1111111111110100;
    assign weights1[16][752] = 16'b1111111111111101;
    assign weights1[16][753] = 16'b1111111111111101;
    assign weights1[16][754] = 16'b1111111111111111;
    assign weights1[16][755] = 16'b0000000000000100;
    assign weights1[16][756] = 16'b1111111111111110;
    assign weights1[16][757] = 16'b1111111111111101;
    assign weights1[16][758] = 16'b1111111111111110;
    assign weights1[16][759] = 16'b0000000000000011;
    assign weights1[16][760] = 16'b0000000000000010;
    assign weights1[16][761] = 16'b1111111111111100;
    assign weights1[16][762] = 16'b0000000000001011;
    assign weights1[16][763] = 16'b0000000000001000;
    assign weights1[16][764] = 16'b0000000000001000;
    assign weights1[16][765] = 16'b1111111111111010;
    assign weights1[16][766] = 16'b1111111111110010;
    assign weights1[16][767] = 16'b1111111111111010;
    assign weights1[16][768] = 16'b0000000000000111;
    assign weights1[16][769] = 16'b1111111111111100;
    assign weights1[16][770] = 16'b1111111111111111;
    assign weights1[16][771] = 16'b0000000000001000;
    assign weights1[16][772] = 16'b1111111111110011;
    assign weights1[16][773] = 16'b1111111111101111;
    assign weights1[16][774] = 16'b1111111111111111;
    assign weights1[16][775] = 16'b0000000000000001;
    assign weights1[16][776] = 16'b1111111111111011;
    assign weights1[16][777] = 16'b1111111111110001;
    assign weights1[16][778] = 16'b1111111111111011;
    assign weights1[16][779] = 16'b1111111111110110;
    assign weights1[16][780] = 16'b1111111111110110;
    assign weights1[16][781] = 16'b1111111111111010;
    assign weights1[16][782] = 16'b1111111111111111;
    assign weights1[16][783] = 16'b0000000000000001;
    assign weights1[17][0] = 16'b0000000000000000;
    assign weights1[17][1] = 16'b0000000000000000;
    assign weights1[17][2] = 16'b1111111111111110;
    assign weights1[17][3] = 16'b0000000000000000;
    assign weights1[17][4] = 16'b1111111111111111;
    assign weights1[17][5] = 16'b1111111111111111;
    assign weights1[17][6] = 16'b1111111111111111;
    assign weights1[17][7] = 16'b0000000000000000;
    assign weights1[17][8] = 16'b0000000000000010;
    assign weights1[17][9] = 16'b0000000000000011;
    assign weights1[17][10] = 16'b1111111111111010;
    assign weights1[17][11] = 16'b1111111111111110;
    assign weights1[17][12] = 16'b0000000000000000;
    assign weights1[17][13] = 16'b1111111111110110;
    assign weights1[17][14] = 16'b0000000000000101;
    assign weights1[17][15] = 16'b1111111111110001;
    assign weights1[17][16] = 16'b1111111111110000;
    assign weights1[17][17] = 16'b1111111111101111;
    assign weights1[17][18] = 16'b1111111111110101;
    assign weights1[17][19] = 16'b1111111111111001;
    assign weights1[17][20] = 16'b1111111111110001;
    assign weights1[17][21] = 16'b1111111111101100;
    assign weights1[17][22] = 16'b1111111111110011;
    assign weights1[17][23] = 16'b1111111111111001;
    assign weights1[17][24] = 16'b1111111111111010;
    assign weights1[17][25] = 16'b0000000000000000;
    assign weights1[17][26] = 16'b0000000000000000;
    assign weights1[17][27] = 16'b0000000000000000;
    assign weights1[17][28] = 16'b0000000000000000;
    assign weights1[17][29] = 16'b1111111111111111;
    assign weights1[17][30] = 16'b1111111111111111;
    assign weights1[17][31] = 16'b1111111111111110;
    assign weights1[17][32] = 16'b1111111111111100;
    assign weights1[17][33] = 16'b1111111111111100;
    assign weights1[17][34] = 16'b1111111111111000;
    assign weights1[17][35] = 16'b1111111111111000;
    assign weights1[17][36] = 16'b1111111111110111;
    assign weights1[17][37] = 16'b0000000000000011;
    assign weights1[17][38] = 16'b0000000000000010;
    assign weights1[17][39] = 16'b0000000000000001;
    assign weights1[17][40] = 16'b0000000000001101;
    assign weights1[17][41] = 16'b0000000000000011;
    assign weights1[17][42] = 16'b0000000000010110;
    assign weights1[17][43] = 16'b1111111111110101;
    assign weights1[17][44] = 16'b1111111111100001;
    assign weights1[17][45] = 16'b1111111111111010;
    assign weights1[17][46] = 16'b0000000000001010;
    assign weights1[17][47] = 16'b1111111111110001;
    assign weights1[17][48] = 16'b1111111111111110;
    assign weights1[17][49] = 16'b1111111111110010;
    assign weights1[17][50] = 16'b1111111111111010;
    assign weights1[17][51] = 16'b1111111111111011;
    assign weights1[17][52] = 16'b1111111111110110;
    assign weights1[17][53] = 16'b1111111111110110;
    assign weights1[17][54] = 16'b1111111111111110;
    assign weights1[17][55] = 16'b1111111111111100;
    assign weights1[17][56] = 16'b1111111111111110;
    assign weights1[17][57] = 16'b1111111111111110;
    assign weights1[17][58] = 16'b1111111111111001;
    assign weights1[17][59] = 16'b1111111111111001;
    assign weights1[17][60] = 16'b1111111111110100;
    assign weights1[17][61] = 16'b1111111111110001;
    assign weights1[17][62] = 16'b1111111111110110;
    assign weights1[17][63] = 16'b1111111111101111;
    assign weights1[17][64] = 16'b1111111111110100;
    assign weights1[17][65] = 16'b1111111111111100;
    assign weights1[17][66] = 16'b1111111111111110;
    assign weights1[17][67] = 16'b0000000000001001;
    assign weights1[17][68] = 16'b0000000000010010;
    assign weights1[17][69] = 16'b0000000000011001;
    assign weights1[17][70] = 16'b0000000000001001;
    assign weights1[17][71] = 16'b0000000000000000;
    assign weights1[17][72] = 16'b1111111111100110;
    assign weights1[17][73] = 16'b1111111111100001;
    assign weights1[17][74] = 16'b0000000000000001;
    assign weights1[17][75] = 16'b1111111111111101;
    assign weights1[17][76] = 16'b1111111111110011;
    assign weights1[17][77] = 16'b1111111111111010;
    assign weights1[17][78] = 16'b0000000000001001;
    assign weights1[17][79] = 16'b1111111111111101;
    assign weights1[17][80] = 16'b1111111111111001;
    assign weights1[17][81] = 16'b1111111111111000;
    assign weights1[17][82] = 16'b1111111111111011;
    assign weights1[17][83] = 16'b1111111111111100;
    assign weights1[17][84] = 16'b1111111111111011;
    assign weights1[17][85] = 16'b1111111111111010;
    assign weights1[17][86] = 16'b1111111111110110;
    assign weights1[17][87] = 16'b1111111111101101;
    assign weights1[17][88] = 16'b1111111111101111;
    assign weights1[17][89] = 16'b1111111111101010;
    assign weights1[17][90] = 16'b1111111111100100;
    assign weights1[17][91] = 16'b1111111111011101;
    assign weights1[17][92] = 16'b1111111111101000;
    assign weights1[17][93] = 16'b1111111111100110;
    assign weights1[17][94] = 16'b1111111111100100;
    assign weights1[17][95] = 16'b0000000000001001;
    assign weights1[17][96] = 16'b0000000000001001;
    assign weights1[17][97] = 16'b1111111111101100;
    assign weights1[17][98] = 16'b1111111111111011;
    assign weights1[17][99] = 16'b1111111111111111;
    assign weights1[17][100] = 16'b1111111111101000;
    assign weights1[17][101] = 16'b1111111111101111;
    assign weights1[17][102] = 16'b1111111111111111;
    assign weights1[17][103] = 16'b0000000000000101;
    assign weights1[17][104] = 16'b0000000000001111;
    assign weights1[17][105] = 16'b1111111111111010;
    assign weights1[17][106] = 16'b1111111111111101;
    assign weights1[17][107] = 16'b1111111111110001;
    assign weights1[17][108] = 16'b0000000000000000;
    assign weights1[17][109] = 16'b1111111111111010;
    assign weights1[17][110] = 16'b1111111111111000;
    assign weights1[17][111] = 16'b1111111111111011;
    assign weights1[17][112] = 16'b1111111111111001;
    assign weights1[17][113] = 16'b1111111111110111;
    assign weights1[17][114] = 16'b1111111111110000;
    assign weights1[17][115] = 16'b1111111111110001;
    assign weights1[17][116] = 16'b1111111111100110;
    assign weights1[17][117] = 16'b1111111111100001;
    assign weights1[17][118] = 16'b1111111111011100;
    assign weights1[17][119] = 16'b1111111111010110;
    assign weights1[17][120] = 16'b1111111111011010;
    assign weights1[17][121] = 16'b1111111110111111;
    assign weights1[17][122] = 16'b1111111111011100;
    assign weights1[17][123] = 16'b1111111111101010;
    assign weights1[17][124] = 16'b0000000000000111;
    assign weights1[17][125] = 16'b0000000000010010;
    assign weights1[17][126] = 16'b0000000000010110;
    assign weights1[17][127] = 16'b0000000000000011;
    assign weights1[17][128] = 16'b1111111111100000;
    assign weights1[17][129] = 16'b1111111111110001;
    assign weights1[17][130] = 16'b1111111111100111;
    assign weights1[17][131] = 16'b1111111111111010;
    assign weights1[17][132] = 16'b1111111111110101;
    assign weights1[17][133] = 16'b0000000000001001;
    assign weights1[17][134] = 16'b0000000000000110;
    assign weights1[17][135] = 16'b0000000000000100;
    assign weights1[17][136] = 16'b0000000000000000;
    assign weights1[17][137] = 16'b1111111111111101;
    assign weights1[17][138] = 16'b1111111111111010;
    assign weights1[17][139] = 16'b1111111111111110;
    assign weights1[17][140] = 16'b1111111111110110;
    assign weights1[17][141] = 16'b1111111111110000;
    assign weights1[17][142] = 16'b1111111111101011;
    assign weights1[17][143] = 16'b1111111111100010;
    assign weights1[17][144] = 16'b1111111111001101;
    assign weights1[17][145] = 16'b1111111111001000;
    assign weights1[17][146] = 16'b1111111111010000;
    assign weights1[17][147] = 16'b1111111111000101;
    assign weights1[17][148] = 16'b1111111111000111;
    assign weights1[17][149] = 16'b1111111111011000;
    assign weights1[17][150] = 16'b1111111111000101;
    assign weights1[17][151] = 16'b1111111111000111;
    assign weights1[17][152] = 16'b1111111111111010;
    assign weights1[17][153] = 16'b0000000000000110;
    assign weights1[17][154] = 16'b0000000000010010;
    assign weights1[17][155] = 16'b0000000000001011;
    assign weights1[17][156] = 16'b0000000000001110;
    assign weights1[17][157] = 16'b1111111111111100;
    assign weights1[17][158] = 16'b1111111111101101;
    assign weights1[17][159] = 16'b1111111111110100;
    assign weights1[17][160] = 16'b1111111111101101;
    assign weights1[17][161] = 16'b1111111111110111;
    assign weights1[17][162] = 16'b1111111111110100;
    assign weights1[17][163] = 16'b0000000000000000;
    assign weights1[17][164] = 16'b1111111111111011;
    assign weights1[17][165] = 16'b1111111111110001;
    assign weights1[17][166] = 16'b1111111111110110;
    assign weights1[17][167] = 16'b1111111111111110;
    assign weights1[17][168] = 16'b1111111111111011;
    assign weights1[17][169] = 16'b1111111111110001;
    assign weights1[17][170] = 16'b1111111111101010;
    assign weights1[17][171] = 16'b1111111111011110;
    assign weights1[17][172] = 16'b1111111111001110;
    assign weights1[17][173] = 16'b1111111111011110;
    assign weights1[17][174] = 16'b1111111111000110;
    assign weights1[17][175] = 16'b1111111111010100;
    assign weights1[17][176] = 16'b0000000000000001;
    assign weights1[17][177] = 16'b1111111111110011;
    assign weights1[17][178] = 16'b1111111111011110;
    assign weights1[17][179] = 16'b1111111111100010;
    assign weights1[17][180] = 16'b0000000000001111;
    assign weights1[17][181] = 16'b0000000000001100;
    assign weights1[17][182] = 16'b0000000000000100;
    assign weights1[17][183] = 16'b1111111111111101;
    assign weights1[17][184] = 16'b1111111111111110;
    assign weights1[17][185] = 16'b0000000000000001;
    assign weights1[17][186] = 16'b1111111111100100;
    assign weights1[17][187] = 16'b1111111111110001;
    assign weights1[17][188] = 16'b1111111111111110;
    assign weights1[17][189] = 16'b0000000000001000;
    assign weights1[17][190] = 16'b1111111111111111;
    assign weights1[17][191] = 16'b0000000000001101;
    assign weights1[17][192] = 16'b0000000000000111;
    assign weights1[17][193] = 16'b1111111111111001;
    assign weights1[17][194] = 16'b1111111111111100;
    assign weights1[17][195] = 16'b1111111111111101;
    assign weights1[17][196] = 16'b1111111111111001;
    assign weights1[17][197] = 16'b1111111111110011;
    assign weights1[17][198] = 16'b1111111111111000;
    assign weights1[17][199] = 16'b1111111111110001;
    assign weights1[17][200] = 16'b1111111111101011;
    assign weights1[17][201] = 16'b1111111111110100;
    assign weights1[17][202] = 16'b1111111111110111;
    assign weights1[17][203] = 16'b0000000000000011;
    assign weights1[17][204] = 16'b1111111111101000;
    assign weights1[17][205] = 16'b0000000000000101;
    assign weights1[17][206] = 16'b1111111111111010;
    assign weights1[17][207] = 16'b1111111111001111;
    assign weights1[17][208] = 16'b1111111111011101;
    assign weights1[17][209] = 16'b0000000000000010;
    assign weights1[17][210] = 16'b1111111111111000;
    assign weights1[17][211] = 16'b1111111111110110;
    assign weights1[17][212] = 16'b0000000000000010;
    assign weights1[17][213] = 16'b1111111111111100;
    assign weights1[17][214] = 16'b1111111111110101;
    assign weights1[17][215] = 16'b0000000000000000;
    assign weights1[17][216] = 16'b1111111111101110;
    assign weights1[17][217] = 16'b0000000000000111;
    assign weights1[17][218] = 16'b1111111111100111;
    assign weights1[17][219] = 16'b0000000000000101;
    assign weights1[17][220] = 16'b1111111111011101;
    assign weights1[17][221] = 16'b1111111111111011;
    assign weights1[17][222] = 16'b1111111111101110;
    assign weights1[17][223] = 16'b1111111111111001;
    assign weights1[17][224] = 16'b0000000000000010;
    assign weights1[17][225] = 16'b0000000000000011;
    assign weights1[17][226] = 16'b1111111111111010;
    assign weights1[17][227] = 16'b0000000000000011;
    assign weights1[17][228] = 16'b0000000000000111;
    assign weights1[17][229] = 16'b0000000000011010;
    assign weights1[17][230] = 16'b0000000000000100;
    assign weights1[17][231] = 16'b1111111111110100;
    assign weights1[17][232] = 16'b1111111111110010;
    assign weights1[17][233] = 16'b0000000000001000;
    assign weights1[17][234] = 16'b0000000000010011;
    assign weights1[17][235] = 16'b1111111111011100;
    assign weights1[17][236] = 16'b1111111111110101;
    assign weights1[17][237] = 16'b0000000000000111;
    assign weights1[17][238] = 16'b0000000000000110;
    assign weights1[17][239] = 16'b0000000000001010;
    assign weights1[17][240] = 16'b1111111111110111;
    assign weights1[17][241] = 16'b1111111111111111;
    assign weights1[17][242] = 16'b1111111111111110;
    assign weights1[17][243] = 16'b1111111111110001;
    assign weights1[17][244] = 16'b1111111111111111;
    assign weights1[17][245] = 16'b1111111111110000;
    assign weights1[17][246] = 16'b1111111111110111;
    assign weights1[17][247] = 16'b0000000000001000;
    assign weights1[17][248] = 16'b1111111111111111;
    assign weights1[17][249] = 16'b1111111111111110;
    assign weights1[17][250] = 16'b1111111111110101;
    assign weights1[17][251] = 16'b1111111111101110;
    assign weights1[17][252] = 16'b0000000000001000;
    assign weights1[17][253] = 16'b0000000000001110;
    assign weights1[17][254] = 16'b0000000000001111;
    assign weights1[17][255] = 16'b1111111111110100;
    assign weights1[17][256] = 16'b0000000000101110;
    assign weights1[17][257] = 16'b0000000000001011;
    assign weights1[17][258] = 16'b0000000000000101;
    assign weights1[17][259] = 16'b0000000000001001;
    assign weights1[17][260] = 16'b1111111111111110;
    assign weights1[17][261] = 16'b0000000000001000;
    assign weights1[17][262] = 16'b0000000000010001;
    assign weights1[17][263] = 16'b1111111111101111;
    assign weights1[17][264] = 16'b1111111111110011;
    assign weights1[17][265] = 16'b0000000000000111;
    assign weights1[17][266] = 16'b0000000000100100;
    assign weights1[17][267] = 16'b0000000000000100;
    assign weights1[17][268] = 16'b1111111111111110;
    assign weights1[17][269] = 16'b1111111111101111;
    assign weights1[17][270] = 16'b1111111111111111;
    assign weights1[17][271] = 16'b1111111111111101;
    assign weights1[17][272] = 16'b1111111111111110;
    assign weights1[17][273] = 16'b1111111111110101;
    assign weights1[17][274] = 16'b0000000000000110;
    assign weights1[17][275] = 16'b1111111111111010;
    assign weights1[17][276] = 16'b1111111111100000;
    assign weights1[17][277] = 16'b1111111111111101;
    assign weights1[17][278] = 16'b1111111111111101;
    assign weights1[17][279] = 16'b1111111111110000;
    assign weights1[17][280] = 16'b0000000000001111;
    assign weights1[17][281] = 16'b0000000000001110;
    assign weights1[17][282] = 16'b0000000000010010;
    assign weights1[17][283] = 16'b0000000000000110;
    assign weights1[17][284] = 16'b0000000000000001;
    assign weights1[17][285] = 16'b0000000000011111;
    assign weights1[17][286] = 16'b0000000000010001;
    assign weights1[17][287] = 16'b0000000000001101;
    assign weights1[17][288] = 16'b0000000000011110;
    assign weights1[17][289] = 16'b1111111111111111;
    assign weights1[17][290] = 16'b0000000000010000;
    assign weights1[17][291] = 16'b0000000000000011;
    assign weights1[17][292] = 16'b1111111111101001;
    assign weights1[17][293] = 16'b0000000000010100;
    assign weights1[17][294] = 16'b0000000000001110;
    assign weights1[17][295] = 16'b1111111111101100;
    assign weights1[17][296] = 16'b1111111111110101;
    assign weights1[17][297] = 16'b1111111111101101;
    assign weights1[17][298] = 16'b1111111111101111;
    assign weights1[17][299] = 16'b1111111111111000;
    assign weights1[17][300] = 16'b1111111111101001;
    assign weights1[17][301] = 16'b0000000000000001;
    assign weights1[17][302] = 16'b1111111111100110;
    assign weights1[17][303] = 16'b1111111111111011;
    assign weights1[17][304] = 16'b1111111111111100;
    assign weights1[17][305] = 16'b0000000000001010;
    assign weights1[17][306] = 16'b1111111111110111;
    assign weights1[17][307] = 16'b1111111111110001;
    assign weights1[17][308] = 16'b0000000000010010;
    assign weights1[17][309] = 16'b0000000000010011;
    assign weights1[17][310] = 16'b0000000000000101;
    assign weights1[17][311] = 16'b0000000000000100;
    assign weights1[17][312] = 16'b1111111111111011;
    assign weights1[17][313] = 16'b0000000000000110;
    assign weights1[17][314] = 16'b0000000000000000;
    assign weights1[17][315] = 16'b1111111111110101;
    assign weights1[17][316] = 16'b0000000000001000;
    assign weights1[17][317] = 16'b0000000000000110;
    assign weights1[17][318] = 16'b0000000000011010;
    assign weights1[17][319] = 16'b0000000000011010;
    assign weights1[17][320] = 16'b1111111111111011;
    assign weights1[17][321] = 16'b1111111111110011;
    assign weights1[17][322] = 16'b1111111111101100;
    assign weights1[17][323] = 16'b1111111111101110;
    assign weights1[17][324] = 16'b1111111111100010;
    assign weights1[17][325] = 16'b1111111111110011;
    assign weights1[17][326] = 16'b1111111111111010;
    assign weights1[17][327] = 16'b1111111111111110;
    assign weights1[17][328] = 16'b1111111111111010;
    assign weights1[17][329] = 16'b1111111111111010;
    assign weights1[17][330] = 16'b1111111111110111;
    assign weights1[17][331] = 16'b1111111111101110;
    assign weights1[17][332] = 16'b1111111111101111;
    assign weights1[17][333] = 16'b1111111111111101;
    assign weights1[17][334] = 16'b1111111111110010;
    assign weights1[17][335] = 16'b1111111111100010;
    assign weights1[17][336] = 16'b0000000000001100;
    assign weights1[17][337] = 16'b0000000000010011;
    assign weights1[17][338] = 16'b0000000000000110;
    assign weights1[17][339] = 16'b1111111111111011;
    assign weights1[17][340] = 16'b1111111111111101;
    assign weights1[17][341] = 16'b0000000000011001;
    assign weights1[17][342] = 16'b0000000000010000;
    assign weights1[17][343] = 16'b0000000000001001;
    assign weights1[17][344] = 16'b0000000000001100;
    assign weights1[17][345] = 16'b0000000000011010;
    assign weights1[17][346] = 16'b0000000000011011;
    assign weights1[17][347] = 16'b0000000000001110;
    assign weights1[17][348] = 16'b1111111111100111;
    assign weights1[17][349] = 16'b1111111110111011;
    assign weights1[17][350] = 16'b1111111111100101;
    assign weights1[17][351] = 16'b1111111111011110;
    assign weights1[17][352] = 16'b1111111111100111;
    assign weights1[17][353] = 16'b1111111111101100;
    assign weights1[17][354] = 16'b1111111111110110;
    assign weights1[17][355] = 16'b1111111111101100;
    assign weights1[17][356] = 16'b1111111111110111;
    assign weights1[17][357] = 16'b1111111111100110;
    assign weights1[17][358] = 16'b1111111111100100;
    assign weights1[17][359] = 16'b1111111111110100;
    assign weights1[17][360] = 16'b1111111111110011;
    assign weights1[17][361] = 16'b1111111111011010;
    assign weights1[17][362] = 16'b1111111111100011;
    assign weights1[17][363] = 16'b1111111111100011;
    assign weights1[17][364] = 16'b0000000000001000;
    assign weights1[17][365] = 16'b0000000000001011;
    assign weights1[17][366] = 16'b0000000000000000;
    assign weights1[17][367] = 16'b1111111111111001;
    assign weights1[17][368] = 16'b1111111111111111;
    assign weights1[17][369] = 16'b0000000000000111;
    assign weights1[17][370] = 16'b0000000000000110;
    assign weights1[17][371] = 16'b0000000000011101;
    assign weights1[17][372] = 16'b0000000000001100;
    assign weights1[17][373] = 16'b0000000000100000;
    assign weights1[17][374] = 16'b0000000000010000;
    assign weights1[17][375] = 16'b0000000000000110;
    assign weights1[17][376] = 16'b1111111110100001;
    assign weights1[17][377] = 16'b1111111111100101;
    assign weights1[17][378] = 16'b1111111111001111;
    assign weights1[17][379] = 16'b1111111111011001;
    assign weights1[17][380] = 16'b1111111111110100;
    assign weights1[17][381] = 16'b1111111111101011;
    assign weights1[17][382] = 16'b1111111111111010;
    assign weights1[17][383] = 16'b1111111111110010;
    assign weights1[17][384] = 16'b1111111111111100;
    assign weights1[17][385] = 16'b1111111111111010;
    assign weights1[17][386] = 16'b1111111111110111;
    assign weights1[17][387] = 16'b1111111111101000;
    assign weights1[17][388] = 16'b1111111111100010;
    assign weights1[17][389] = 16'b1111111111100101;
    assign weights1[17][390] = 16'b1111111111011001;
    assign weights1[17][391] = 16'b1111111111100111;
    assign weights1[17][392] = 16'b0000000000000111;
    assign weights1[17][393] = 16'b0000000000001101;
    assign weights1[17][394] = 16'b0000000000000101;
    assign weights1[17][395] = 16'b0000000000001101;
    assign weights1[17][396] = 16'b1111111111111000;
    assign weights1[17][397] = 16'b0000000000010010;
    assign weights1[17][398] = 16'b0000000000001011;
    assign weights1[17][399] = 16'b0000000000100001;
    assign weights1[17][400] = 16'b0000000000011011;
    assign weights1[17][401] = 16'b0000000000001001;
    assign weights1[17][402] = 16'b0000000000001000;
    assign weights1[17][403] = 16'b1111111110101101;
    assign weights1[17][404] = 16'b1111111101101101;
    assign weights1[17][405] = 16'b1111111111000111;
    assign weights1[17][406] = 16'b1111111111010010;
    assign weights1[17][407] = 16'b1111111111101101;
    assign weights1[17][408] = 16'b1111111111110010;
    assign weights1[17][409] = 16'b1111111111111010;
    assign weights1[17][410] = 16'b1111111111110010;
    assign weights1[17][411] = 16'b0000000000000010;
    assign weights1[17][412] = 16'b1111111111111010;
    assign weights1[17][413] = 16'b1111111111101111;
    assign weights1[17][414] = 16'b1111111111100100;
    assign weights1[17][415] = 16'b1111111111100110;
    assign weights1[17][416] = 16'b1111111111011110;
    assign weights1[17][417] = 16'b1111111111101101;
    assign weights1[17][418] = 16'b1111111111110101;
    assign weights1[17][419] = 16'b1111111111111000;
    assign weights1[17][420] = 16'b0000000000000011;
    assign weights1[17][421] = 16'b0000000000010000;
    assign weights1[17][422] = 16'b0000000000001110;
    assign weights1[17][423] = 16'b0000000000100111;
    assign weights1[17][424] = 16'b1111111111111010;
    assign weights1[17][425] = 16'b0000000000101100;
    assign weights1[17][426] = 16'b0000000000100001;
    assign weights1[17][427] = 16'b0000000000000000;
    assign weights1[17][428] = 16'b0000000000101101;
    assign weights1[17][429] = 16'b1111111111111111;
    assign weights1[17][430] = 16'b1111111110011011;
    assign weights1[17][431] = 16'b1111111101000000;
    assign weights1[17][432] = 16'b1111111110000101;
    assign weights1[17][433] = 16'b1111111111100111;
    assign weights1[17][434] = 16'b1111111111100101;
    assign weights1[17][435] = 16'b0000000000000000;
    assign weights1[17][436] = 16'b1111111111100101;
    assign weights1[17][437] = 16'b1111111111110100;
    assign weights1[17][438] = 16'b1111111111111011;
    assign weights1[17][439] = 16'b1111111111110011;
    assign weights1[17][440] = 16'b1111111111111110;
    assign weights1[17][441] = 16'b1111111111101110;
    assign weights1[17][442] = 16'b0000000000000001;
    assign weights1[17][443] = 16'b1111111111110000;
    assign weights1[17][444] = 16'b0000000000001011;
    assign weights1[17][445] = 16'b1111111111101001;
    assign weights1[17][446] = 16'b1111111111101100;
    assign weights1[17][447] = 16'b1111111111111000;
    assign weights1[17][448] = 16'b0000000000000000;
    assign weights1[17][449] = 16'b0000000000000111;
    assign weights1[17][450] = 16'b0000000000010001;
    assign weights1[17][451] = 16'b0000000000010110;
    assign weights1[17][452] = 16'b0000000000100000;
    assign weights1[17][453] = 16'b0000000000010101;
    assign weights1[17][454] = 16'b0000000000001110;
    assign weights1[17][455] = 16'b0000000000011100;
    assign weights1[17][456] = 16'b1111111111101011;
    assign weights1[17][457] = 16'b1111111110101001;
    assign weights1[17][458] = 16'b1111111100010000;
    assign weights1[17][459] = 16'b1111111101011111;
    assign weights1[17][460] = 16'b1111111111100010;
    assign weights1[17][461] = 16'b1111111111111110;
    assign weights1[17][462] = 16'b0000000000000001;
    assign weights1[17][463] = 16'b0000000000010110;
    assign weights1[17][464] = 16'b1111111111111011;
    assign weights1[17][465] = 16'b0000000000001100;
    assign weights1[17][466] = 16'b0000000000001010;
    assign weights1[17][467] = 16'b0000000000000100;
    assign weights1[17][468] = 16'b0000000000000111;
    assign weights1[17][469] = 16'b0000000000100011;
    assign weights1[17][470] = 16'b0000000000000010;
    assign weights1[17][471] = 16'b0000000000001100;
    assign weights1[17][472] = 16'b1111111111110011;
    assign weights1[17][473] = 16'b1111111111111000;
    assign weights1[17][474] = 16'b1111111111110111;
    assign weights1[17][475] = 16'b0000000000010100;
    assign weights1[17][476] = 16'b1111111111110000;
    assign weights1[17][477] = 16'b0000000000001001;
    assign weights1[17][478] = 16'b1111111111101111;
    assign weights1[17][479] = 16'b1111111111110000;
    assign weights1[17][480] = 16'b0000000000011011;
    assign weights1[17][481] = 16'b0000000000000100;
    assign weights1[17][482] = 16'b1111111111011101;
    assign weights1[17][483] = 16'b1111111111001111;
    assign weights1[17][484] = 16'b1111111101111010;
    assign weights1[17][485] = 16'b1111111100101001;
    assign weights1[17][486] = 16'b1111111101001110;
    assign weights1[17][487] = 16'b1111111111001100;
    assign weights1[17][488] = 16'b0000000000001101;
    assign weights1[17][489] = 16'b0000000000001001;
    assign weights1[17][490] = 16'b1111111111111101;
    assign weights1[17][491] = 16'b1111111111110001;
    assign weights1[17][492] = 16'b0000000000000010;
    assign weights1[17][493] = 16'b0000000000000110;
    assign weights1[17][494] = 16'b0000000000011001;
    assign weights1[17][495] = 16'b0000000000000100;
    assign weights1[17][496] = 16'b1111111111101110;
    assign weights1[17][497] = 16'b1111111111110000;
    assign weights1[17][498] = 16'b1111111111111110;
    assign weights1[17][499] = 16'b1111111111111100;
    assign weights1[17][500] = 16'b0000000000000000;
    assign weights1[17][501] = 16'b0000000000011111;
    assign weights1[17][502] = 16'b0000000000011111;
    assign weights1[17][503] = 16'b0000000000011010;
    assign weights1[17][504] = 16'b1111111111101110;
    assign weights1[17][505] = 16'b1111111111110101;
    assign weights1[17][506] = 16'b1111111111101100;
    assign weights1[17][507] = 16'b1111111111010000;
    assign weights1[17][508] = 16'b1111111111100000;
    assign weights1[17][509] = 16'b1111111111011011;
    assign weights1[17][510] = 16'b1111111110110000;
    assign weights1[17][511] = 16'b1111111110001010;
    assign weights1[17][512] = 16'b1111111100101101;
    assign weights1[17][513] = 16'b1111111101010101;
    assign weights1[17][514] = 16'b1111111111010101;
    assign weights1[17][515] = 16'b0000000000000011;
    assign weights1[17][516] = 16'b0000000000001100;
    assign weights1[17][517] = 16'b0000000000010001;
    assign weights1[17][518] = 16'b0000000000011101;
    assign weights1[17][519] = 16'b0000000000010100;
    assign weights1[17][520] = 16'b1111111111111001;
    assign weights1[17][521] = 16'b0000000000010111;
    assign weights1[17][522] = 16'b0000000000001000;
    assign weights1[17][523] = 16'b0000000000010101;
    assign weights1[17][524] = 16'b0000000000001100;
    assign weights1[17][525] = 16'b0000000000000111;
    assign weights1[17][526] = 16'b0000000000010111;
    assign weights1[17][527] = 16'b1111111111111110;
    assign weights1[17][528] = 16'b0000000000000000;
    assign weights1[17][529] = 16'b0000000000100001;
    assign weights1[17][530] = 16'b0000000000011001;
    assign weights1[17][531] = 16'b0000000000101101;
    assign weights1[17][532] = 16'b1111111111100101;
    assign weights1[17][533] = 16'b1111111111101001;
    assign weights1[17][534] = 16'b1111111111010101;
    assign weights1[17][535] = 16'b1111111111010100;
    assign weights1[17][536] = 16'b1111111111001010;
    assign weights1[17][537] = 16'b1111111110101010;
    assign weights1[17][538] = 16'b1111111110000010;
    assign weights1[17][539] = 16'b1111111101010101;
    assign weights1[17][540] = 16'b1111111101101011;
    assign weights1[17][541] = 16'b1111111111001000;
    assign weights1[17][542] = 16'b1111111111111111;
    assign weights1[17][543] = 16'b1111111111110101;
    assign weights1[17][544] = 16'b1111111111111000;
    assign weights1[17][545] = 16'b0000000000000110;
    assign weights1[17][546] = 16'b1111111111111001;
    assign weights1[17][547] = 16'b0000000000001011;
    assign weights1[17][548] = 16'b0000000000000000;
    assign weights1[17][549] = 16'b0000000000001000;
    assign weights1[17][550] = 16'b0000000000001010;
    assign weights1[17][551] = 16'b0000000000001000;
    assign weights1[17][552] = 16'b0000000000011000;
    assign weights1[17][553] = 16'b0000000000000111;
    assign weights1[17][554] = 16'b1111111111111001;
    assign weights1[17][555] = 16'b0000000000010100;
    assign weights1[17][556] = 16'b0000000000100001;
    assign weights1[17][557] = 16'b0000000000001001;
    assign weights1[17][558] = 16'b0000000000011111;
    assign weights1[17][559] = 16'b0000000000101011;
    assign weights1[17][560] = 16'b1111111111011011;
    assign weights1[17][561] = 16'b1111111111010100;
    assign weights1[17][562] = 16'b1111111111000001;
    assign weights1[17][563] = 16'b1111111110111111;
    assign weights1[17][564] = 16'b1111111110100010;
    assign weights1[17][565] = 16'b1111111101111011;
    assign weights1[17][566] = 16'b1111111101110000;
    assign weights1[17][567] = 16'b1111111110001110;
    assign weights1[17][568] = 16'b1111111111011100;
    assign weights1[17][569] = 16'b0000000000000101;
    assign weights1[17][570] = 16'b0000000000001010;
    assign weights1[17][571] = 16'b0000000000001111;
    assign weights1[17][572] = 16'b0000000000010101;
    assign weights1[17][573] = 16'b0000000000000010;
    assign weights1[17][574] = 16'b0000000000010100;
    assign weights1[17][575] = 16'b0000000000010110;
    assign weights1[17][576] = 16'b0000000000000010;
    assign weights1[17][577] = 16'b0000000000000100;
    assign weights1[17][578] = 16'b0000000000001000;
    assign weights1[17][579] = 16'b1111111111111101;
    assign weights1[17][580] = 16'b0000000000001010;
    assign weights1[17][581] = 16'b0000000000001010;
    assign weights1[17][582] = 16'b0000000000000100;
    assign weights1[17][583] = 16'b0000000000001001;
    assign weights1[17][584] = 16'b0000000000011010;
    assign weights1[17][585] = 16'b0000000000000111;
    assign weights1[17][586] = 16'b0000000000010011;
    assign weights1[17][587] = 16'b0000000000011011;
    assign weights1[17][588] = 16'b1111111111011111;
    assign weights1[17][589] = 16'b1111111111010010;
    assign weights1[17][590] = 16'b1111111111000000;
    assign weights1[17][591] = 16'b1111111110110011;
    assign weights1[17][592] = 16'b1111111110010100;
    assign weights1[17][593] = 16'b1111111110010010;
    assign weights1[17][594] = 16'b1111111110100110;
    assign weights1[17][595] = 16'b1111111111011101;
    assign weights1[17][596] = 16'b0000000000001010;
    assign weights1[17][597] = 16'b0000000000010100;
    assign weights1[17][598] = 16'b0000000000001101;
    assign weights1[17][599] = 16'b0000000000010110;
    assign weights1[17][600] = 16'b0000000000001110;
    assign weights1[17][601] = 16'b0000000000011000;
    assign weights1[17][602] = 16'b0000000000001000;
    assign weights1[17][603] = 16'b0000000000010110;
    assign weights1[17][604] = 16'b0000000000010110;
    assign weights1[17][605] = 16'b0000000000010011;
    assign weights1[17][606] = 16'b0000000000000001;
    assign weights1[17][607] = 16'b0000000000000100;
    assign weights1[17][608] = 16'b0000000000000101;
    assign weights1[17][609] = 16'b0000000000000001;
    assign weights1[17][610] = 16'b0000000000010011;
    assign weights1[17][611] = 16'b0000000000011000;
    assign weights1[17][612] = 16'b0000000000001110;
    assign weights1[17][613] = 16'b0000000000011011;
    assign weights1[17][614] = 16'b0000000000011011;
    assign weights1[17][615] = 16'b0000000000101101;
    assign weights1[17][616] = 16'b1111111111010110;
    assign weights1[17][617] = 16'b1111111111001110;
    assign weights1[17][618] = 16'b1111111111001101;
    assign weights1[17][619] = 16'b1111111110111010;
    assign weights1[17][620] = 16'b1111111110011100;
    assign weights1[17][621] = 16'b1111111110110001;
    assign weights1[17][622] = 16'b1111111111101100;
    assign weights1[17][623] = 16'b0000000000100010;
    assign weights1[17][624] = 16'b0000000000010111;
    assign weights1[17][625] = 16'b0000000000011011;
    assign weights1[17][626] = 16'b0000000000001011;
    assign weights1[17][627] = 16'b0000000000001111;
    assign weights1[17][628] = 16'b0000000000011011;
    assign weights1[17][629] = 16'b0000000000001111;
    assign weights1[17][630] = 16'b0000000000011011;
    assign weights1[17][631] = 16'b0000000000010000;
    assign weights1[17][632] = 16'b1111111111110101;
    assign weights1[17][633] = 16'b0000000000000101;
    assign weights1[17][634] = 16'b1111111111110100;
    assign weights1[17][635] = 16'b1111111111110001;
    assign weights1[17][636] = 16'b1111111111111011;
    assign weights1[17][637] = 16'b0000000000001010;
    assign weights1[17][638] = 16'b0000000000001110;
    assign weights1[17][639] = 16'b0000000000011101;
    assign weights1[17][640] = 16'b0000000000011010;
    assign weights1[17][641] = 16'b0000000000001111;
    assign weights1[17][642] = 16'b0000000000001110;
    assign weights1[17][643] = 16'b0000000000011001;
    assign weights1[17][644] = 16'b1111111111011100;
    assign weights1[17][645] = 16'b1111111111001010;
    assign weights1[17][646] = 16'b1111111111001010;
    assign weights1[17][647] = 16'b1111111111001010;
    assign weights1[17][648] = 16'b1111111111010001;
    assign weights1[17][649] = 16'b1111111111111110;
    assign weights1[17][650] = 16'b0000000000000111;
    assign weights1[17][651] = 16'b0000000000011110;
    assign weights1[17][652] = 16'b1111111111111000;
    assign weights1[17][653] = 16'b0000000000001011;
    assign weights1[17][654] = 16'b0000000000011101;
    assign weights1[17][655] = 16'b0000000000010001;
    assign weights1[17][656] = 16'b0000000000001000;
    assign weights1[17][657] = 16'b0000000000000100;
    assign weights1[17][658] = 16'b0000000000001110;
    assign weights1[17][659] = 16'b0000000000010111;
    assign weights1[17][660] = 16'b0000000000001001;
    assign weights1[17][661] = 16'b0000000000001101;
    assign weights1[17][662] = 16'b0000000000000011;
    assign weights1[17][663] = 16'b0000000000001101;
    assign weights1[17][664] = 16'b0000000000000000;
    assign weights1[17][665] = 16'b0000000000010111;
    assign weights1[17][666] = 16'b1111111111111110;
    assign weights1[17][667] = 16'b0000000000001101;
    assign weights1[17][668] = 16'b0000000000100011;
    assign weights1[17][669] = 16'b0000000000010110;
    assign weights1[17][670] = 16'b0000000000010100;
    assign weights1[17][671] = 16'b0000000000010110;
    assign weights1[17][672] = 16'b1111111111100110;
    assign weights1[17][673] = 16'b1111111111011010;
    assign weights1[17][674] = 16'b1111111111000011;
    assign weights1[17][675] = 16'b1111111111011011;
    assign weights1[17][676] = 16'b1111111111100110;
    assign weights1[17][677] = 16'b1111111111110001;
    assign weights1[17][678] = 16'b0000000000101001;
    assign weights1[17][679] = 16'b0000000000010011;
    assign weights1[17][680] = 16'b0000000000000110;
    assign weights1[17][681] = 16'b0000000000010001;
    assign weights1[17][682] = 16'b1111111111111100;
    assign weights1[17][683] = 16'b0000000000000110;
    assign weights1[17][684] = 16'b1111111111110011;
    assign weights1[17][685] = 16'b1111111111111111;
    assign weights1[17][686] = 16'b0000000000001100;
    assign weights1[17][687] = 16'b1111111111110111;
    assign weights1[17][688] = 16'b1111111111111110;
    assign weights1[17][689] = 16'b0000000000010010;
    assign weights1[17][690] = 16'b0000000000010000;
    assign weights1[17][691] = 16'b0000000000000101;
    assign weights1[17][692] = 16'b0000000000000110;
    assign weights1[17][693] = 16'b1111111111111100;
    assign weights1[17][694] = 16'b0000000000001011;
    assign weights1[17][695] = 16'b0000000000010010;
    assign weights1[17][696] = 16'b0000000000010111;
    assign weights1[17][697] = 16'b0000000000001011;
    assign weights1[17][698] = 16'b0000000000001100;
    assign weights1[17][699] = 16'b0000000000010011;
    assign weights1[17][700] = 16'b1111111111110101;
    assign weights1[17][701] = 16'b1111111111100110;
    assign weights1[17][702] = 16'b1111111111011111;
    assign weights1[17][703] = 16'b1111111111100101;
    assign weights1[17][704] = 16'b1111111111100111;
    assign weights1[17][705] = 16'b1111111111111111;
    assign weights1[17][706] = 16'b0000000000001111;
    assign weights1[17][707] = 16'b0000000000001010;
    assign weights1[17][708] = 16'b0000000000001110;
    assign weights1[17][709] = 16'b0000000000011110;
    assign weights1[17][710] = 16'b0000000000000001;
    assign weights1[17][711] = 16'b0000000000011101;
    assign weights1[17][712] = 16'b0000000000010101;
    assign weights1[17][713] = 16'b1111111111111101;
    assign weights1[17][714] = 16'b1111111111111011;
    assign weights1[17][715] = 16'b1111111111110101;
    assign weights1[17][716] = 16'b1111111111111111;
    assign weights1[17][717] = 16'b0000000000000011;
    assign weights1[17][718] = 16'b0000000000001101;
    assign weights1[17][719] = 16'b0000000000001010;
    assign weights1[17][720] = 16'b1111111111111010;
    assign weights1[17][721] = 16'b0000000000010101;
    assign weights1[17][722] = 16'b0000000000000000;
    assign weights1[17][723] = 16'b1111111111111101;
    assign weights1[17][724] = 16'b0000000000001010;
    assign weights1[17][725] = 16'b0000000000001111;
    assign weights1[17][726] = 16'b0000000000000100;
    assign weights1[17][727] = 16'b0000000000000111;
    assign weights1[17][728] = 16'b1111111111111110;
    assign weights1[17][729] = 16'b1111111111111110;
    assign weights1[17][730] = 16'b1111111111110111;
    assign weights1[17][731] = 16'b0000000000000001;
    assign weights1[17][732] = 16'b0000000000010001;
    assign weights1[17][733] = 16'b1111111111111101;
    assign weights1[17][734] = 16'b0000000000001000;
    assign weights1[17][735] = 16'b0000000000001101;
    assign weights1[17][736] = 16'b0000000000100100;
    assign weights1[17][737] = 16'b0000000000001100;
    assign weights1[17][738] = 16'b1111111111111011;
    assign weights1[17][739] = 16'b0000000000010111;
    assign weights1[17][740] = 16'b0000000000000011;
    assign weights1[17][741] = 16'b0000000000001011;
    assign weights1[17][742] = 16'b1111111111111110;
    assign weights1[17][743] = 16'b0000000000000011;
    assign weights1[17][744] = 16'b0000000000001001;
    assign weights1[17][745] = 16'b0000000000000101;
    assign weights1[17][746] = 16'b0000000000000000;
    assign weights1[17][747] = 16'b0000000000001101;
    assign weights1[17][748] = 16'b0000000000000001;
    assign weights1[17][749] = 16'b0000000000001100;
    assign weights1[17][750] = 16'b1111111111111100;
    assign weights1[17][751] = 16'b0000000000000000;
    assign weights1[17][752] = 16'b0000000000000100;
    assign weights1[17][753] = 16'b0000000000000111;
    assign weights1[17][754] = 16'b0000000000001101;
    assign weights1[17][755] = 16'b0000000000000101;
    assign weights1[17][756] = 16'b1111111111111111;
    assign weights1[17][757] = 16'b0000000000000011;
    assign weights1[17][758] = 16'b0000000000001101;
    assign weights1[17][759] = 16'b0000000000010100;
    assign weights1[17][760] = 16'b0000000000001100;
    assign weights1[17][761] = 16'b0000000000001110;
    assign weights1[17][762] = 16'b0000000000010011;
    assign weights1[17][763] = 16'b0000000000010100;
    assign weights1[17][764] = 16'b0000000000010000;
    assign weights1[17][765] = 16'b0000000000010000;
    assign weights1[17][766] = 16'b0000000000101011;
    assign weights1[17][767] = 16'b0000000000001000;
    assign weights1[17][768] = 16'b0000000000000110;
    assign weights1[17][769] = 16'b1111111111111011;
    assign weights1[17][770] = 16'b0000000000000001;
    assign weights1[17][771] = 16'b1111111111110001;
    assign weights1[17][772] = 16'b1111111111110101;
    assign weights1[17][773] = 16'b1111111111111000;
    assign weights1[17][774] = 16'b0000000000000100;
    assign weights1[17][775] = 16'b1111111111110110;
    assign weights1[17][776] = 16'b0000000000000111;
    assign weights1[17][777] = 16'b0000000000000010;
    assign weights1[17][778] = 16'b1111111111110111;
    assign weights1[17][779] = 16'b0000000000001001;
    assign weights1[17][780] = 16'b1111111111111011;
    assign weights1[17][781] = 16'b1111111111111110;
    assign weights1[17][782] = 16'b0000000000000010;
    assign weights1[17][783] = 16'b0000000000000010;
    assign weights1[18][0] = 16'b0000000000000000;
    assign weights1[18][1] = 16'b0000000000000000;
    assign weights1[18][2] = 16'b0000000000000001;
    assign weights1[18][3] = 16'b0000000000000010;
    assign weights1[18][4] = 16'b1111111111111110;
    assign weights1[18][5] = 16'b0000000000000100;
    assign weights1[18][6] = 16'b0000000000000000;
    assign weights1[18][7] = 16'b1111111111111101;
    assign weights1[18][8] = 16'b0000000000001000;
    assign weights1[18][9] = 16'b1111111111111100;
    assign weights1[18][10] = 16'b1111111111111111;
    assign weights1[18][11] = 16'b0000000000010011;
    assign weights1[18][12] = 16'b0000000000010111;
    assign weights1[18][13] = 16'b0000000000001010;
    assign weights1[18][14] = 16'b0000000000001101;
    assign weights1[18][15] = 16'b0000000000000110;
    assign weights1[18][16] = 16'b1111111111110110;
    assign weights1[18][17] = 16'b1111111111111101;
    assign weights1[18][18] = 16'b1111111111101101;
    assign weights1[18][19] = 16'b0000000000001000;
    assign weights1[18][20] = 16'b0000000000001011;
    assign weights1[18][21] = 16'b0000000000000110;
    assign weights1[18][22] = 16'b0000000000000100;
    assign weights1[18][23] = 16'b1111111111110110;
    assign weights1[18][24] = 16'b1111111111111111;
    assign weights1[18][25] = 16'b0000000000000010;
    assign weights1[18][26] = 16'b0000000000000011;
    assign weights1[18][27] = 16'b1111111111111110;
    assign weights1[18][28] = 16'b0000000000000000;
    assign weights1[18][29] = 16'b0000000000000000;
    assign weights1[18][30] = 16'b0000000000000001;
    assign weights1[18][31] = 16'b0000000000000101;
    assign weights1[18][32] = 16'b0000000000000101;
    assign weights1[18][33] = 16'b0000000000000110;
    assign weights1[18][34] = 16'b0000000000000010;
    assign weights1[18][35] = 16'b1111111111110100;
    assign weights1[18][36] = 16'b0000000000000101;
    assign weights1[18][37] = 16'b1111111111110011;
    assign weights1[18][38] = 16'b1111111111110111;
    assign weights1[18][39] = 16'b1111111111111110;
    assign weights1[18][40] = 16'b0000000000000011;
    assign weights1[18][41] = 16'b0000000000000101;
    assign weights1[18][42] = 16'b1111111111110010;
    assign weights1[18][43] = 16'b0000000000001011;
    assign weights1[18][44] = 16'b0000000000001010;
    assign weights1[18][45] = 16'b0000000000001011;
    assign weights1[18][46] = 16'b0000000000000110;
    assign weights1[18][47] = 16'b1111111111111000;
    assign weights1[18][48] = 16'b1111111111111010;
    assign weights1[18][49] = 16'b1111111111111111;
    assign weights1[18][50] = 16'b0000000000000010;
    assign weights1[18][51] = 16'b1111111111111010;
    assign weights1[18][52] = 16'b1111111111111101;
    assign weights1[18][53] = 16'b1111111111111100;
    assign weights1[18][54] = 16'b1111111111110111;
    assign weights1[18][55] = 16'b1111111111111111;
    assign weights1[18][56] = 16'b1111111111111111;
    assign weights1[18][57] = 16'b0000000000000001;
    assign weights1[18][58] = 16'b0000000000000011;
    assign weights1[18][59] = 16'b0000000000001001;
    assign weights1[18][60] = 16'b0000000000001000;
    assign weights1[18][61] = 16'b0000000000000101;
    assign weights1[18][62] = 16'b0000000000001100;
    assign weights1[18][63] = 16'b1111111111101010;
    assign weights1[18][64] = 16'b0000000000000000;
    assign weights1[18][65] = 16'b1111111111101110;
    assign weights1[18][66] = 16'b1111111111100110;
    assign weights1[18][67] = 16'b1111111111011101;
    assign weights1[18][68] = 16'b1111111111011111;
    assign weights1[18][69] = 16'b1111111111111101;
    assign weights1[18][70] = 16'b0000000000000101;
    assign weights1[18][71] = 16'b1111111111110010;
    assign weights1[18][72] = 16'b1111111111111111;
    assign weights1[18][73] = 16'b0000000000000011;
    assign weights1[18][74] = 16'b0000000000000100;
    assign weights1[18][75] = 16'b0000000000001111;
    assign weights1[18][76] = 16'b0000000000000111;
    assign weights1[18][77] = 16'b0000000000000001;
    assign weights1[18][78] = 16'b0000000000001011;
    assign weights1[18][79] = 16'b1111111111111010;
    assign weights1[18][80] = 16'b0000000000001011;
    assign weights1[18][81] = 16'b0000000000000001;
    assign weights1[18][82] = 16'b0000000000000001;
    assign weights1[18][83] = 16'b1111111111111111;
    assign weights1[18][84] = 16'b0000000000000001;
    assign weights1[18][85] = 16'b0000000000000011;
    assign weights1[18][86] = 16'b0000000000000010;
    assign weights1[18][87] = 16'b0000000000000110;
    assign weights1[18][88] = 16'b1111111111111111;
    assign weights1[18][89] = 16'b0000000000010000;
    assign weights1[18][90] = 16'b0000000000001111;
    assign weights1[18][91] = 16'b0000000000011000;
    assign weights1[18][92] = 16'b0000000000011101;
    assign weights1[18][93] = 16'b0000000000000100;
    assign weights1[18][94] = 16'b0000000000001100;
    assign weights1[18][95] = 16'b1111111111111110;
    assign weights1[18][96] = 16'b0000000000000100;
    assign weights1[18][97] = 16'b0000000000000100;
    assign weights1[18][98] = 16'b0000000000001101;
    assign weights1[18][99] = 16'b0000000000001000;
    assign weights1[18][100] = 16'b0000000000000111;
    assign weights1[18][101] = 16'b0000000000001111;
    assign weights1[18][102] = 16'b1111111111101010;
    assign weights1[18][103] = 16'b0000000000000010;
    assign weights1[18][104] = 16'b0000000000000000;
    assign weights1[18][105] = 16'b0000000000010000;
    assign weights1[18][106] = 16'b1111111111111110;
    assign weights1[18][107] = 16'b1111111111110111;
    assign weights1[18][108] = 16'b0000000000000011;
    assign weights1[18][109] = 16'b1111111111110001;
    assign weights1[18][110] = 16'b1111111111111001;
    assign weights1[18][111] = 16'b0000000000000111;
    assign weights1[18][112] = 16'b0000000000001000;
    assign weights1[18][113] = 16'b0000000000001001;
    assign weights1[18][114] = 16'b0000000000000100;
    assign weights1[18][115] = 16'b1111111111111001;
    assign weights1[18][116] = 16'b0000000000011000;
    assign weights1[18][117] = 16'b0000000000100000;
    assign weights1[18][118] = 16'b0000000000010110;
    assign weights1[18][119] = 16'b0000000000100111;
    assign weights1[18][120] = 16'b0000000000010001;
    assign weights1[18][121] = 16'b0000000000101110;
    assign weights1[18][122] = 16'b0000000000100110;
    assign weights1[18][123] = 16'b0000000000011011;
    assign weights1[18][124] = 16'b0000000000011001;
    assign weights1[18][125] = 16'b0000000000000100;
    assign weights1[18][126] = 16'b1111111111101100;
    assign weights1[18][127] = 16'b1111111111101110;
    assign weights1[18][128] = 16'b1111111111101111;
    assign weights1[18][129] = 16'b1111111111110111;
    assign weights1[18][130] = 16'b0000000000010000;
    assign weights1[18][131] = 16'b1111111111111111;
    assign weights1[18][132] = 16'b1111111111111010;
    assign weights1[18][133] = 16'b1111111111101111;
    assign weights1[18][134] = 16'b0000000000001001;
    assign weights1[18][135] = 16'b0000000000000010;
    assign weights1[18][136] = 16'b0000000000001110;
    assign weights1[18][137] = 16'b1111111111110010;
    assign weights1[18][138] = 16'b0000000000000100;
    assign weights1[18][139] = 16'b1111111111111111;
    assign weights1[18][140] = 16'b0000000000001000;
    assign weights1[18][141] = 16'b0000000000001101;
    assign weights1[18][142] = 16'b0000000000000101;
    assign weights1[18][143] = 16'b0000000000100001;
    assign weights1[18][144] = 16'b0000000000110000;
    assign weights1[18][145] = 16'b0000000000100011;
    assign weights1[18][146] = 16'b0000000000010110;
    assign weights1[18][147] = 16'b0000000000010111;
    assign weights1[18][148] = 16'b0000000000010001;
    assign weights1[18][149] = 16'b0000000000010110;
    assign weights1[18][150] = 16'b1111111111111100;
    assign weights1[18][151] = 16'b1111111111101011;
    assign weights1[18][152] = 16'b0000000000000011;
    assign weights1[18][153] = 16'b1111111111111010;
    assign weights1[18][154] = 16'b0000000000001010;
    assign weights1[18][155] = 16'b1111111111111101;
    assign weights1[18][156] = 16'b0000000000010101;
    assign weights1[18][157] = 16'b0000000000001010;
    assign weights1[18][158] = 16'b1111111111110111;
    assign weights1[18][159] = 16'b1111111111110101;
    assign weights1[18][160] = 16'b0000000000001101;
    assign weights1[18][161] = 16'b1111111111111110;
    assign weights1[18][162] = 16'b0000000000010011;
    assign weights1[18][163] = 16'b1111111111111110;
    assign weights1[18][164] = 16'b1111111111110001;
    assign weights1[18][165] = 16'b1111111111111111;
    assign weights1[18][166] = 16'b1111111111110110;
    assign weights1[18][167] = 16'b1111111111110000;
    assign weights1[18][168] = 16'b0000000000000100;
    assign weights1[18][169] = 16'b0000000000001110;
    assign weights1[18][170] = 16'b0000000000011001;
    assign weights1[18][171] = 16'b0000000000101100;
    assign weights1[18][172] = 16'b0000000000111100;
    assign weights1[18][173] = 16'b0000000000010111;
    assign weights1[18][174] = 16'b0000000000010011;
    assign weights1[18][175] = 16'b0000000000011001;
    assign weights1[18][176] = 16'b0000000000001011;
    assign weights1[18][177] = 16'b0000000000011010;
    assign weights1[18][178] = 16'b0000000000011100;
    assign weights1[18][179] = 16'b0000000000010111;
    assign weights1[18][180] = 16'b0000000000011000;
    assign weights1[18][181] = 16'b1111111111110101;
    assign weights1[18][182] = 16'b0000000000100111;
    assign weights1[18][183] = 16'b1111111111111101;
    assign weights1[18][184] = 16'b0000000000000101;
    assign weights1[18][185] = 16'b1111111111110011;
    assign weights1[18][186] = 16'b0000000000010001;
    assign weights1[18][187] = 16'b0000000000010000;
    assign weights1[18][188] = 16'b1111111111111110;
    assign weights1[18][189] = 16'b1111111111101110;
    assign weights1[18][190] = 16'b0000000000010000;
    assign weights1[18][191] = 16'b0000000000000110;
    assign weights1[18][192] = 16'b1111111111101000;
    assign weights1[18][193] = 16'b1111111111111110;
    assign weights1[18][194] = 16'b1111111111111111;
    assign weights1[18][195] = 16'b1111111111111100;
    assign weights1[18][196] = 16'b0000000000000100;
    assign weights1[18][197] = 16'b0000000000010101;
    assign weights1[18][198] = 16'b0000000000100101;
    assign weights1[18][199] = 16'b0000000000111000;
    assign weights1[18][200] = 16'b0000000001000001;
    assign weights1[18][201] = 16'b0000000000110111;
    assign weights1[18][202] = 16'b0000000001100111;
    assign weights1[18][203] = 16'b0000000000110010;
    assign weights1[18][204] = 16'b0000000000100101;
    assign weights1[18][205] = 16'b0000000000110000;
    assign weights1[18][206] = 16'b0000000000111001;
    assign weights1[18][207] = 16'b0000000000110000;
    assign weights1[18][208] = 16'b0000000000010001;
    assign weights1[18][209] = 16'b0000000000100110;
    assign weights1[18][210] = 16'b0000000000010010;
    assign weights1[18][211] = 16'b0000000000010001;
    assign weights1[18][212] = 16'b0000000000001111;
    assign weights1[18][213] = 16'b0000000000010110;
    assign weights1[18][214] = 16'b0000000000000110;
    assign weights1[18][215] = 16'b1111111111111111;
    assign weights1[18][216] = 16'b0000000000000111;
    assign weights1[18][217] = 16'b0000000000000111;
    assign weights1[18][218] = 16'b0000000000000111;
    assign weights1[18][219] = 16'b1111111111101110;
    assign weights1[18][220] = 16'b0000000000001100;
    assign weights1[18][221] = 16'b1111111111110011;
    assign weights1[18][222] = 16'b0000000000000010;
    assign weights1[18][223] = 16'b0000000000000000;
    assign weights1[18][224] = 16'b0000000000000111;
    assign weights1[18][225] = 16'b0000000000001010;
    assign weights1[18][226] = 16'b0000000000010111;
    assign weights1[18][227] = 16'b0000000000101111;
    assign weights1[18][228] = 16'b0000000001001111;
    assign weights1[18][229] = 16'b0000000000110111;
    assign weights1[18][230] = 16'b0000000001010110;
    assign weights1[18][231] = 16'b0000000001000000;
    assign weights1[18][232] = 16'b0000000001011111;
    assign weights1[18][233] = 16'b0000000000111011;
    assign weights1[18][234] = 16'b0000000001000001;
    assign weights1[18][235] = 16'b0000000001000001;
    assign weights1[18][236] = 16'b0000000000101100;
    assign weights1[18][237] = 16'b0000000000110010;
    assign weights1[18][238] = 16'b0000000000100110;
    assign weights1[18][239] = 16'b0000000000010111;
    assign weights1[18][240] = 16'b0000000000001101;
    assign weights1[18][241] = 16'b0000000000011010;
    assign weights1[18][242] = 16'b0000000000001111;
    assign weights1[18][243] = 16'b0000000000001000;
    assign weights1[18][244] = 16'b0000000000010110;
    assign weights1[18][245] = 16'b0000000000000101;
    assign weights1[18][246] = 16'b0000000000000100;
    assign weights1[18][247] = 16'b1111111111101001;
    assign weights1[18][248] = 16'b0000000000001011;
    assign weights1[18][249] = 16'b0000000000001010;
    assign weights1[18][250] = 16'b0000000000000101;
    assign weights1[18][251] = 16'b0000000000001010;
    assign weights1[18][252] = 16'b0000000000000000;
    assign weights1[18][253] = 16'b1111111111101111;
    assign weights1[18][254] = 16'b1111111111111001;
    assign weights1[18][255] = 16'b0000000000001001;
    assign weights1[18][256] = 16'b0000000000011011;
    assign weights1[18][257] = 16'b0000000000001110;
    assign weights1[18][258] = 16'b0000000000010011;
    assign weights1[18][259] = 16'b0000000000100001;
    assign weights1[18][260] = 16'b0000000000110111;
    assign weights1[18][261] = 16'b0000000000001111;
    assign weights1[18][262] = 16'b0000000000011011;
    assign weights1[18][263] = 16'b0000000000101111;
    assign weights1[18][264] = 16'b0000000000100100;
    assign weights1[18][265] = 16'b0000000000010000;
    assign weights1[18][266] = 16'b0000000000001010;
    assign weights1[18][267] = 16'b0000000000010001;
    assign weights1[18][268] = 16'b0000000000000001;
    assign weights1[18][269] = 16'b1111111111110111;
    assign weights1[18][270] = 16'b0000000000000101;
    assign weights1[18][271] = 16'b0000000000000010;
    assign weights1[18][272] = 16'b1111111111111001;
    assign weights1[18][273] = 16'b0000000000010000;
    assign weights1[18][274] = 16'b0000000000010010;
    assign weights1[18][275] = 16'b1111111111111100;
    assign weights1[18][276] = 16'b0000000000000010;
    assign weights1[18][277] = 16'b0000000000000110;
    assign weights1[18][278] = 16'b0000000000001110;
    assign weights1[18][279] = 16'b0000000000001001;
    assign weights1[18][280] = 16'b1111111111101011;
    assign weights1[18][281] = 16'b1111111111001001;
    assign weights1[18][282] = 16'b1111111110111011;
    assign weights1[18][283] = 16'b1111111110111000;
    assign weights1[18][284] = 16'b1111111110101100;
    assign weights1[18][285] = 16'b1111111110111100;
    assign weights1[18][286] = 16'b1111111111000010;
    assign weights1[18][287] = 16'b1111111110111001;
    assign weights1[18][288] = 16'b1111111110111001;
    assign weights1[18][289] = 16'b1111111111001001;
    assign weights1[18][290] = 16'b1111111110111010;
    assign weights1[18][291] = 16'b1111111110011100;
    assign weights1[18][292] = 16'b1111111110111100;
    assign weights1[18][293] = 16'b1111111110110111;
    assign weights1[18][294] = 16'b1111111110111000;
    assign weights1[18][295] = 16'b1111111110111100;
    assign weights1[18][296] = 16'b1111111111110000;
    assign weights1[18][297] = 16'b1111111111110001;
    assign weights1[18][298] = 16'b1111111111101101;
    assign weights1[18][299] = 16'b1111111111110100;
    assign weights1[18][300] = 16'b1111111111111111;
    assign weights1[18][301] = 16'b1111111111110110;
    assign weights1[18][302] = 16'b1111111111110001;
    assign weights1[18][303] = 16'b0000000000000111;
    assign weights1[18][304] = 16'b1111111111101100;
    assign weights1[18][305] = 16'b0000000000010011;
    assign weights1[18][306] = 16'b1111111111111111;
    assign weights1[18][307] = 16'b0000000000010000;
    assign weights1[18][308] = 16'b1111111111000010;
    assign weights1[18][309] = 16'b1111111110010101;
    assign weights1[18][310] = 16'b1111111110000110;
    assign weights1[18][311] = 16'b1111111101111011;
    assign weights1[18][312] = 16'b1111111101010001;
    assign weights1[18][313] = 16'b1111111101001000;
    assign weights1[18][314] = 16'b1111111101001000;
    assign weights1[18][315] = 16'b1111111100110110;
    assign weights1[18][316] = 16'b1111111100000011;
    assign weights1[18][317] = 16'b1111111100001101;
    assign weights1[18][318] = 16'b1111111100101111;
    assign weights1[18][319] = 16'b1111111101100001;
    assign weights1[18][320] = 16'b1111111101111110;
    assign weights1[18][321] = 16'b1111111110011101;
    assign weights1[18][322] = 16'b1111111111010001;
    assign weights1[18][323] = 16'b1111111111001101;
    assign weights1[18][324] = 16'b1111111111100011;
    assign weights1[18][325] = 16'b1111111111110010;
    assign weights1[18][326] = 16'b1111111111100101;
    assign weights1[18][327] = 16'b1111111111110101;
    assign weights1[18][328] = 16'b1111111111111011;
    assign weights1[18][329] = 16'b1111111111100111;
    assign weights1[18][330] = 16'b1111111111111101;
    assign weights1[18][331] = 16'b1111111111111110;
    assign weights1[18][332] = 16'b0000000000000100;
    assign weights1[18][333] = 16'b0000000000001010;
    assign weights1[18][334] = 16'b0000000000000100;
    assign weights1[18][335] = 16'b1111111111110110;
    assign weights1[18][336] = 16'b1111111110110100;
    assign weights1[18][337] = 16'b1111111110001011;
    assign weights1[18][338] = 16'b1111111101110001;
    assign weights1[18][339] = 16'b1111111101001100;
    assign weights1[18][340] = 16'b1111111100110000;
    assign weights1[18][341] = 16'b1111111100001000;
    assign weights1[18][342] = 16'b1111111011101101;
    assign weights1[18][343] = 16'b1111111011010010;
    assign weights1[18][344] = 16'b1111111100000101;
    assign weights1[18][345] = 16'b1111111101100000;
    assign weights1[18][346] = 16'b1111111110101001;
    assign weights1[18][347] = 16'b1111111111000000;
    assign weights1[18][348] = 16'b1111111111100101;
    assign weights1[18][349] = 16'b1111111111101100;
    assign weights1[18][350] = 16'b1111111111111011;
    assign weights1[18][351] = 16'b1111111111111010;
    assign weights1[18][352] = 16'b0000000000001110;
    assign weights1[18][353] = 16'b1111111111110101;
    assign weights1[18][354] = 16'b0000000000001101;
    assign weights1[18][355] = 16'b1111111111111110;
    assign weights1[18][356] = 16'b0000000000001011;
    assign weights1[18][357] = 16'b0000000000000100;
    assign weights1[18][358] = 16'b0000000000000011;
    assign weights1[18][359] = 16'b0000000000000010;
    assign weights1[18][360] = 16'b1111111111111000;
    assign weights1[18][361] = 16'b0000000000001101;
    assign weights1[18][362] = 16'b1111111111110110;
    assign weights1[18][363] = 16'b1111111111111011;
    assign weights1[18][364] = 16'b1111111110110000;
    assign weights1[18][365] = 16'b1111111110010001;
    assign weights1[18][366] = 16'b1111111110000000;
    assign weights1[18][367] = 16'b1111111101101001;
    assign weights1[18][368] = 16'b1111111101011001;
    assign weights1[18][369] = 16'b1111111101110011;
    assign weights1[18][370] = 16'b1111111110001010;
    assign weights1[18][371] = 16'b1111111111001001;
    assign weights1[18][372] = 16'b0000000000001001;
    assign weights1[18][373] = 16'b0000000000001101;
    assign weights1[18][374] = 16'b0000000000011000;
    assign weights1[18][375] = 16'b0000000000011001;
    assign weights1[18][376] = 16'b0000000000010100;
    assign weights1[18][377] = 16'b0000000000010001;
    assign weights1[18][378] = 16'b0000000000001011;
    assign weights1[18][379] = 16'b0000000000000110;
    assign weights1[18][380] = 16'b0000000000001110;
    assign weights1[18][381] = 16'b1111111111110011;
    assign weights1[18][382] = 16'b1111111111111100;
    assign weights1[18][383] = 16'b0000000000000000;
    assign weights1[18][384] = 16'b1111111111110110;
    assign weights1[18][385] = 16'b0000000000011001;
    assign weights1[18][386] = 16'b0000000000000101;
    assign weights1[18][387] = 16'b0000000000000011;
    assign weights1[18][388] = 16'b1111111111111010;
    assign weights1[18][389] = 16'b0000000000001100;
    assign weights1[18][390] = 16'b1111111111111111;
    assign weights1[18][391] = 16'b0000000000000011;
    assign weights1[18][392] = 16'b1111111111000111;
    assign weights1[18][393] = 16'b1111111110101011;
    assign weights1[18][394] = 16'b1111111110110011;
    assign weights1[18][395] = 16'b1111111110111111;
    assign weights1[18][396] = 16'b1111111111011100;
    assign weights1[18][397] = 16'b0000000000010011;
    assign weights1[18][398] = 16'b0000000001000000;
    assign weights1[18][399] = 16'b0000000001001110;
    assign weights1[18][400] = 16'b0000000000111000;
    assign weights1[18][401] = 16'b0000000000111001;
    assign weights1[18][402] = 16'b0000000000101010;
    assign weights1[18][403] = 16'b0000000000100110;
    assign weights1[18][404] = 16'b0000000000011100;
    assign weights1[18][405] = 16'b0000000000001011;
    assign weights1[18][406] = 16'b0000000000011010;
    assign weights1[18][407] = 16'b0000000000000011;
    assign weights1[18][408] = 16'b0000000000000100;
    assign weights1[18][409] = 16'b0000000000000011;
    assign weights1[18][410] = 16'b0000000000001000;
    assign weights1[18][411] = 16'b0000000000000110;
    assign weights1[18][412] = 16'b0000000000001001;
    assign weights1[18][413] = 16'b1111111111111111;
    assign weights1[18][414] = 16'b0000000000000110;
    assign weights1[18][415] = 16'b0000000000000011;
    assign weights1[18][416] = 16'b1111111111111000;
    assign weights1[18][417] = 16'b1111111111111100;
    assign weights1[18][418] = 16'b1111111111110111;
    assign weights1[18][419] = 16'b1111111111111010;
    assign weights1[18][420] = 16'b1111111111011000;
    assign weights1[18][421] = 16'b1111111111010111;
    assign weights1[18][422] = 16'b1111111111100101;
    assign weights1[18][423] = 16'b1111111111110110;
    assign weights1[18][424] = 16'b0000000000100001;
    assign weights1[18][425] = 16'b0000000000111101;
    assign weights1[18][426] = 16'b0000000000111011;
    assign weights1[18][427] = 16'b0000000000111111;
    assign weights1[18][428] = 16'b0000000000100000;
    assign weights1[18][429] = 16'b0000000000010010;
    assign weights1[18][430] = 16'b0000000000001001;
    assign weights1[18][431] = 16'b0000000000011111;
    assign weights1[18][432] = 16'b0000000000000010;
    assign weights1[18][433] = 16'b1111111111111111;
    assign weights1[18][434] = 16'b1111111111111000;
    assign weights1[18][435] = 16'b0000000000001011;
    assign weights1[18][436] = 16'b0000000000010010;
    assign weights1[18][437] = 16'b0000000000001100;
    assign weights1[18][438] = 16'b0000000000000000;
    assign weights1[18][439] = 16'b0000000000000100;
    assign weights1[18][440] = 16'b1111111111110010;
    assign weights1[18][441] = 16'b1111111111110101;
    assign weights1[18][442] = 16'b0000000000000001;
    assign weights1[18][443] = 16'b0000000000000000;
    assign weights1[18][444] = 16'b0000000000000000;
    assign weights1[18][445] = 16'b0000000000000010;
    assign weights1[18][446] = 16'b0000000000000110;
    assign weights1[18][447] = 16'b0000000000010011;
    assign weights1[18][448] = 16'b1111111111110110;
    assign weights1[18][449] = 16'b0000000000000010;
    assign weights1[18][450] = 16'b0000000000010010;
    assign weights1[18][451] = 16'b0000000000011010;
    assign weights1[18][452] = 16'b0000000000111111;
    assign weights1[18][453] = 16'b0000000000000100;
    assign weights1[18][454] = 16'b0000000000100100;
    assign weights1[18][455] = 16'b0000000000011101;
    assign weights1[18][456] = 16'b0000000000010001;
    assign weights1[18][457] = 16'b0000000000001100;
    assign weights1[18][458] = 16'b0000000000000001;
    assign weights1[18][459] = 16'b1111111111110100;
    assign weights1[18][460] = 16'b0000000000000100;
    assign weights1[18][461] = 16'b1111111111111011;
    assign weights1[18][462] = 16'b0000000000000101;
    assign weights1[18][463] = 16'b1111111111110111;
    assign weights1[18][464] = 16'b0000000000000010;
    assign weights1[18][465] = 16'b1111111111110100;
    assign weights1[18][466] = 16'b0000000000001010;
    assign weights1[18][467] = 16'b0000000000001100;
    assign weights1[18][468] = 16'b0000000000010000;
    assign weights1[18][469] = 16'b1111111111111101;
    assign weights1[18][470] = 16'b0000000000001000;
    assign weights1[18][471] = 16'b0000000000001001;
    assign weights1[18][472] = 16'b0000000000001100;
    assign weights1[18][473] = 16'b0000000000010101;
    assign weights1[18][474] = 16'b0000000000010111;
    assign weights1[18][475] = 16'b0000000000001000;
    assign weights1[18][476] = 16'b0000000000001101;
    assign weights1[18][477] = 16'b0000000000100000;
    assign weights1[18][478] = 16'b0000000000010011;
    assign weights1[18][479] = 16'b1111111111111111;
    assign weights1[18][480] = 16'b0000000000010011;
    assign weights1[18][481] = 16'b1111111111111101;
    assign weights1[18][482] = 16'b1111111111110000;
    assign weights1[18][483] = 16'b1111111111111100;
    assign weights1[18][484] = 16'b1111111111101111;
    assign weights1[18][485] = 16'b0000000000000000;
    assign weights1[18][486] = 16'b1111111111111100;
    assign weights1[18][487] = 16'b0000000000001101;
    assign weights1[18][488] = 16'b1111111111110101;
    assign weights1[18][489] = 16'b0000000000000011;
    assign weights1[18][490] = 16'b0000000000000001;
    assign weights1[18][491] = 16'b1111111111110110;
    assign weights1[18][492] = 16'b0000000000000101;
    assign weights1[18][493] = 16'b1111111111110111;
    assign weights1[18][494] = 16'b1111111111111101;
    assign weights1[18][495] = 16'b1111111111110101;
    assign weights1[18][496] = 16'b0000000000000111;
    assign weights1[18][497] = 16'b0000000000001011;
    assign weights1[18][498] = 16'b0000000000000101;
    assign weights1[18][499] = 16'b0000000000000110;
    assign weights1[18][500] = 16'b1111111111111100;
    assign weights1[18][501] = 16'b0000000000000011;
    assign weights1[18][502] = 16'b0000000000000000;
    assign weights1[18][503] = 16'b1111111111111110;
    assign weights1[18][504] = 16'b0000000000100100;
    assign weights1[18][505] = 16'b0000000000010000;
    assign weights1[18][506] = 16'b0000000000011000;
    assign weights1[18][507] = 16'b0000000000001011;
    assign weights1[18][508] = 16'b0000000000010111;
    assign weights1[18][509] = 16'b0000000000000101;
    assign weights1[18][510] = 16'b0000000000011011;
    assign weights1[18][511] = 16'b0000000000011110;
    assign weights1[18][512] = 16'b0000000000000011;
    assign weights1[18][513] = 16'b0000000000010110;
    assign weights1[18][514] = 16'b0000000000000001;
    assign weights1[18][515] = 16'b1111111111110011;
    assign weights1[18][516] = 16'b0000000000000011;
    assign weights1[18][517] = 16'b1111111111111010;
    assign weights1[18][518] = 16'b1111111111111100;
    assign weights1[18][519] = 16'b1111111111111000;
    assign weights1[18][520] = 16'b1111111111110011;
    assign weights1[18][521] = 16'b1111111111110111;
    assign weights1[18][522] = 16'b1111111111110110;
    assign weights1[18][523] = 16'b1111111111111111;
    assign weights1[18][524] = 16'b1111111111111001;
    assign weights1[18][525] = 16'b1111111111101101;
    assign weights1[18][526] = 16'b1111111111101010;
    assign weights1[18][527] = 16'b0000000000000000;
    assign weights1[18][528] = 16'b1111111111110111;
    assign weights1[18][529] = 16'b0000000000000110;
    assign weights1[18][530] = 16'b0000000000000011;
    assign weights1[18][531] = 16'b1111111111111111;
    assign weights1[18][532] = 16'b0000000000010110;
    assign weights1[18][533] = 16'b0000000000001011;
    assign weights1[18][534] = 16'b0000000000001110;
    assign weights1[18][535] = 16'b1111111111111110;
    assign weights1[18][536] = 16'b0000000000000011;
    assign weights1[18][537] = 16'b1111111111101101;
    assign weights1[18][538] = 16'b1111111111101110;
    assign weights1[18][539] = 16'b0000000000001001;
    assign weights1[18][540] = 16'b1111111111110001;
    assign weights1[18][541] = 16'b1111111111110001;
    assign weights1[18][542] = 16'b1111111111111001;
    assign weights1[18][543] = 16'b0000000000001011;
    assign weights1[18][544] = 16'b1111111111101111;
    assign weights1[18][545] = 16'b0000000000001010;
    assign weights1[18][546] = 16'b0000000000001101;
    assign weights1[18][547] = 16'b1111111111111101;
    assign weights1[18][548] = 16'b0000000000001001;
    assign weights1[18][549] = 16'b1111111111111110;
    assign weights1[18][550] = 16'b1111111111111000;
    assign weights1[18][551] = 16'b0000000000000001;
    assign weights1[18][552] = 16'b1111111111111111;
    assign weights1[18][553] = 16'b1111111111111110;
    assign weights1[18][554] = 16'b0000000000000111;
    assign weights1[18][555] = 16'b0000000000000001;
    assign weights1[18][556] = 16'b1111111111111010;
    assign weights1[18][557] = 16'b1111111111110110;
    assign weights1[18][558] = 16'b1111111111111111;
    assign weights1[18][559] = 16'b0000000000000001;
    assign weights1[18][560] = 16'b0000000000001001;
    assign weights1[18][561] = 16'b0000000000010100;
    assign weights1[18][562] = 16'b1111111111111001;
    assign weights1[18][563] = 16'b0000000000010001;
    assign weights1[18][564] = 16'b0000000000001010;
    assign weights1[18][565] = 16'b0000000000001111;
    assign weights1[18][566] = 16'b0000000000001100;
    assign weights1[18][567] = 16'b1111111111111101;
    assign weights1[18][568] = 16'b1111111111111110;
    assign weights1[18][569] = 16'b0000000000001000;
    assign weights1[18][570] = 16'b0000000000000000;
    assign weights1[18][571] = 16'b0000000000001010;
    assign weights1[18][572] = 16'b1111111111111101;
    assign weights1[18][573] = 16'b1111111111110100;
    assign weights1[18][574] = 16'b1111111111111100;
    assign weights1[18][575] = 16'b1111111111110110;
    assign weights1[18][576] = 16'b0000000000001001;
    assign weights1[18][577] = 16'b1111111111111111;
    assign weights1[18][578] = 16'b1111111111110100;
    assign weights1[18][579] = 16'b1111111111111000;
    assign weights1[18][580] = 16'b1111111111111000;
    assign weights1[18][581] = 16'b1111111111101000;
    assign weights1[18][582] = 16'b1111111111101010;
    assign weights1[18][583] = 16'b1111111111101001;
    assign weights1[18][584] = 16'b1111111111101110;
    assign weights1[18][585] = 16'b1111111111110010;
    assign weights1[18][586] = 16'b1111111111110011;
    assign weights1[18][587] = 16'b1111111111111000;
    assign weights1[18][588] = 16'b0000000000000001;
    assign weights1[18][589] = 16'b1111111111111010;
    assign weights1[18][590] = 16'b1111111111110110;
    assign weights1[18][591] = 16'b0000000000001000;
    assign weights1[18][592] = 16'b0000000000000011;
    assign weights1[18][593] = 16'b1111111111110101;
    assign weights1[18][594] = 16'b1111111111110000;
    assign weights1[18][595] = 16'b1111111111111111;
    assign weights1[18][596] = 16'b0000000000010011;
    assign weights1[18][597] = 16'b0000000000001110;
    assign weights1[18][598] = 16'b0000000000010100;
    assign weights1[18][599] = 16'b0000000000001101;
    assign weights1[18][600] = 16'b0000000000001010;
    assign weights1[18][601] = 16'b0000000000001001;
    assign weights1[18][602] = 16'b0000000000000100;
    assign weights1[18][603] = 16'b1111111111110101;
    assign weights1[18][604] = 16'b1111111111110100;
    assign weights1[18][605] = 16'b1111111111111010;
    assign weights1[18][606] = 16'b1111111111111111;
    assign weights1[18][607] = 16'b0000000000000011;
    assign weights1[18][608] = 16'b0000000000010101;
    assign weights1[18][609] = 16'b0000000000000010;
    assign weights1[18][610] = 16'b1111111111110011;
    assign weights1[18][611] = 16'b0000000000001100;
    assign weights1[18][612] = 16'b1111111111111001;
    assign weights1[18][613] = 16'b1111111111110101;
    assign weights1[18][614] = 16'b1111111111101110;
    assign weights1[18][615] = 16'b0000000000000001;
    assign weights1[18][616] = 16'b1111111111111001;
    assign weights1[18][617] = 16'b1111111111101111;
    assign weights1[18][618] = 16'b1111111111101110;
    assign weights1[18][619] = 16'b1111111111111011;
    assign weights1[18][620] = 16'b1111111111110100;
    assign weights1[18][621] = 16'b0000000000000011;
    assign weights1[18][622] = 16'b1111111111111101;
    assign weights1[18][623] = 16'b0000000000000010;
    assign weights1[18][624] = 16'b1111111111111101;
    assign weights1[18][625] = 16'b1111111111101001;
    assign weights1[18][626] = 16'b1111111111110000;
    assign weights1[18][627] = 16'b1111111111110100;
    assign weights1[18][628] = 16'b1111111111111110;
    assign weights1[18][629] = 16'b0000000000000000;
    assign weights1[18][630] = 16'b1111111111110100;
    assign weights1[18][631] = 16'b0000000000000111;
    assign weights1[18][632] = 16'b0000000000000011;
    assign weights1[18][633] = 16'b1111111111111001;
    assign weights1[18][634] = 16'b1111111111111100;
    assign weights1[18][635] = 16'b0000000000001110;
    assign weights1[18][636] = 16'b0000000000000011;
    assign weights1[18][637] = 16'b0000000000000011;
    assign weights1[18][638] = 16'b0000000000000100;
    assign weights1[18][639] = 16'b1111111111111100;
    assign weights1[18][640] = 16'b0000000000001001;
    assign weights1[18][641] = 16'b0000000000001000;
    assign weights1[18][642] = 16'b1111111111110101;
    assign weights1[18][643] = 16'b1111111111111110;
    assign weights1[18][644] = 16'b1111111111110101;
    assign weights1[18][645] = 16'b1111111111101111;
    assign weights1[18][646] = 16'b1111111111110001;
    assign weights1[18][647] = 16'b1111111111101110;
    assign weights1[18][648] = 16'b1111111111111011;
    assign weights1[18][649] = 16'b1111111111111001;
    assign weights1[18][650] = 16'b0000000000000010;
    assign weights1[18][651] = 16'b1111111111111010;
    assign weights1[18][652] = 16'b0000000000001010;
    assign weights1[18][653] = 16'b0000000000001111;
    assign weights1[18][654] = 16'b1111111111110101;
    assign weights1[18][655] = 16'b0000000000000100;
    assign weights1[18][656] = 16'b1111111111111000;
    assign weights1[18][657] = 16'b1111111111110110;
    assign weights1[18][658] = 16'b0000000000001100;
    assign weights1[18][659] = 16'b0000000000000001;
    assign weights1[18][660] = 16'b1111111111110111;
    assign weights1[18][661] = 16'b1111111111110010;
    assign weights1[18][662] = 16'b1111111111101100;
    assign weights1[18][663] = 16'b1111111111110101;
    assign weights1[18][664] = 16'b1111111111111010;
    assign weights1[18][665] = 16'b0000000000001110;
    assign weights1[18][666] = 16'b1111111111111110;
    assign weights1[18][667] = 16'b1111111111110011;
    assign weights1[18][668] = 16'b0000000000000101;
    assign weights1[18][669] = 16'b1111111111111111;
    assign weights1[18][670] = 16'b1111111111111100;
    assign weights1[18][671] = 16'b0000000000000101;
    assign weights1[18][672] = 16'b1111111111111001;
    assign weights1[18][673] = 16'b1111111111101011;
    assign weights1[18][674] = 16'b1111111111110011;
    assign weights1[18][675] = 16'b1111111111111010;
    assign weights1[18][676] = 16'b0000000000000000;
    assign weights1[18][677] = 16'b0000000000001010;
    assign weights1[18][678] = 16'b1111111111110110;
    assign weights1[18][679] = 16'b1111111111110111;
    assign weights1[18][680] = 16'b1111111111110101;
    assign weights1[18][681] = 16'b1111111111110100;
    assign weights1[18][682] = 16'b0000000000000100;
    assign weights1[18][683] = 16'b0000000000001110;
    assign weights1[18][684] = 16'b1111111111110101;
    assign weights1[18][685] = 16'b0000000000000001;
    assign weights1[18][686] = 16'b1111111111101010;
    assign weights1[18][687] = 16'b0000000000001100;
    assign weights1[18][688] = 16'b1111111111111000;
    assign weights1[18][689] = 16'b0000000000000000;
    assign weights1[18][690] = 16'b0000000000000010;
    assign weights1[18][691] = 16'b1111111111110110;
    assign weights1[18][692] = 16'b0000000000001001;
    assign weights1[18][693] = 16'b0000000000000011;
    assign weights1[18][694] = 16'b0000000000010010;
    assign weights1[18][695] = 16'b1111111111111100;
    assign weights1[18][696] = 16'b0000000000000010;
    assign weights1[18][697] = 16'b0000000000000100;
    assign weights1[18][698] = 16'b0000000000000110;
    assign weights1[18][699] = 16'b0000000000000011;
    assign weights1[18][700] = 16'b1111111111111110;
    assign weights1[18][701] = 16'b1111111111101101;
    assign weights1[18][702] = 16'b1111111111110011;
    assign weights1[18][703] = 16'b1111111111111001;
    assign weights1[18][704] = 16'b1111111111111101;
    assign weights1[18][705] = 16'b0000000000000100;
    assign weights1[18][706] = 16'b1111111111111101;
    assign weights1[18][707] = 16'b1111111111111011;
    assign weights1[18][708] = 16'b1111111111111101;
    assign weights1[18][709] = 16'b0000000000010101;
    assign weights1[18][710] = 16'b1111111111111100;
    assign weights1[18][711] = 16'b1111111111110111;
    assign weights1[18][712] = 16'b0000000000001011;
    assign weights1[18][713] = 16'b1111111111111011;
    assign weights1[18][714] = 16'b0000000000001000;
    assign weights1[18][715] = 16'b0000000000000101;
    assign weights1[18][716] = 16'b1111111111111111;
    assign weights1[18][717] = 16'b0000000000010000;
    assign weights1[18][718] = 16'b1111111111110001;
    assign weights1[18][719] = 16'b1111111111110101;
    assign weights1[18][720] = 16'b1111111111111110;
    assign weights1[18][721] = 16'b1111111111110111;
    assign weights1[18][722] = 16'b0000000000001111;
    assign weights1[18][723] = 16'b0000000000001000;
    assign weights1[18][724] = 16'b0000000000010001;
    assign weights1[18][725] = 16'b0000000000001001;
    assign weights1[18][726] = 16'b0000000000001001;
    assign weights1[18][727] = 16'b0000000000000001;
    assign weights1[18][728] = 16'b0000000000000000;
    assign weights1[18][729] = 16'b0000000000000010;
    assign weights1[18][730] = 16'b1111111111110101;
    assign weights1[18][731] = 16'b1111111111110001;
    assign weights1[18][732] = 16'b1111111111110010;
    assign weights1[18][733] = 16'b1111111111101110;
    assign weights1[18][734] = 16'b1111111111110001;
    assign weights1[18][735] = 16'b1111111111110111;
    assign weights1[18][736] = 16'b1111111111110010;
    assign weights1[18][737] = 16'b1111111111101110;
    assign weights1[18][738] = 16'b1111111111110110;
    assign weights1[18][739] = 16'b1111111111111000;
    assign weights1[18][740] = 16'b1111111111110110;
    assign weights1[18][741] = 16'b1111111111111010;
    assign weights1[18][742] = 16'b1111111111101101;
    assign weights1[18][743] = 16'b1111111111110100;
    assign weights1[18][744] = 16'b0000000000000001;
    assign weights1[18][745] = 16'b0000000000000010;
    assign weights1[18][746] = 16'b0000000000000110;
    assign weights1[18][747] = 16'b0000000000001011;
    assign weights1[18][748] = 16'b0000000000000100;
    assign weights1[18][749] = 16'b0000000000001001;
    assign weights1[18][750] = 16'b1111111111111101;
    assign weights1[18][751] = 16'b0000000000000001;
    assign weights1[18][752] = 16'b0000000000000110;
    assign weights1[18][753] = 16'b0000000000000110;
    assign weights1[18][754] = 16'b0000000000000100;
    assign weights1[18][755] = 16'b0000000000000000;
    assign weights1[18][756] = 16'b1111111111111110;
    assign weights1[18][757] = 16'b0000000000000000;
    assign weights1[18][758] = 16'b1111111111111001;
    assign weights1[18][759] = 16'b1111111111110111;
    assign weights1[18][760] = 16'b1111111111111001;
    assign weights1[18][761] = 16'b0000000000000100;
    assign weights1[18][762] = 16'b1111111111111100;
    assign weights1[18][763] = 16'b1111111111110001;
    assign weights1[18][764] = 16'b1111111111110110;
    assign weights1[18][765] = 16'b0000000000000110;
    assign weights1[18][766] = 16'b0000000000001100;
    assign weights1[18][767] = 16'b0000000000000111;
    assign weights1[18][768] = 16'b0000000000000001;
    assign weights1[18][769] = 16'b1111111111110110;
    assign weights1[18][770] = 16'b1111111111111100;
    assign weights1[18][771] = 16'b0000000000001010;
    assign weights1[18][772] = 16'b0000000000001101;
    assign weights1[18][773] = 16'b0000000000001001;
    assign weights1[18][774] = 16'b0000000000001001;
    assign weights1[18][775] = 16'b0000000000000111;
    assign weights1[18][776] = 16'b0000000000001000;
    assign weights1[18][777] = 16'b0000000000000111;
    assign weights1[18][778] = 16'b1111111111111011;
    assign weights1[18][779] = 16'b0000000000000110;
    assign weights1[18][780] = 16'b0000000000001010;
    assign weights1[18][781] = 16'b0000000000001011;
    assign weights1[18][782] = 16'b0000000000000010;
    assign weights1[18][783] = 16'b1111111111111111;
    assign weights1[19][0] = 16'b0000000000000000;
    assign weights1[19][1] = 16'b0000000000000000;
    assign weights1[19][2] = 16'b1111111111111111;
    assign weights1[19][3] = 16'b1111111111111111;
    assign weights1[19][4] = 16'b0000000000000000;
    assign weights1[19][5] = 16'b1111111111111101;
    assign weights1[19][6] = 16'b1111111111111100;
    assign weights1[19][7] = 16'b1111111111111110;
    assign weights1[19][8] = 16'b0000000000000010;
    assign weights1[19][9] = 16'b0000000000000001;
    assign weights1[19][10] = 16'b0000000000000111;
    assign weights1[19][11] = 16'b0000000000011101;
    assign weights1[19][12] = 16'b0000000000110001;
    assign weights1[19][13] = 16'b0000000000011101;
    assign weights1[19][14] = 16'b0000000000100001;
    assign weights1[19][15] = 16'b0000000000011011;
    assign weights1[19][16] = 16'b0000000000000110;
    assign weights1[19][17] = 16'b0000000000010010;
    assign weights1[19][18] = 16'b0000000000000101;
    assign weights1[19][19] = 16'b1111111111111001;
    assign weights1[19][20] = 16'b1111111111110000;
    assign weights1[19][21] = 16'b1111111111110101;
    assign weights1[19][22] = 16'b1111111111110010;
    assign weights1[19][23] = 16'b1111111111101101;
    assign weights1[19][24] = 16'b1111111111111000;
    assign weights1[19][25] = 16'b1111111111111100;
    assign weights1[19][26] = 16'b1111111111111010;
    assign weights1[19][27] = 16'b1111111111111101;
    assign weights1[19][28] = 16'b0000000000000000;
    assign weights1[19][29] = 16'b1111111111111111;
    assign weights1[19][30] = 16'b1111111111111101;
    assign weights1[19][31] = 16'b1111111111111110;
    assign weights1[19][32] = 16'b1111111111111011;
    assign weights1[19][33] = 16'b1111111111101111;
    assign weights1[19][34] = 16'b1111111111100111;
    assign weights1[19][35] = 16'b1111111111100110;
    assign weights1[19][36] = 16'b1111111111101001;
    assign weights1[19][37] = 16'b1111111111110101;
    assign weights1[19][38] = 16'b0000000000001011;
    assign weights1[19][39] = 16'b0000000000011111;
    assign weights1[19][40] = 16'b0000000000101011;
    assign weights1[19][41] = 16'b0000000000100111;
    assign weights1[19][42] = 16'b0000000000101111;
    assign weights1[19][43] = 16'b0000000000100011;
    assign weights1[19][44] = 16'b0000000000010010;
    assign weights1[19][45] = 16'b0000000000010111;
    assign weights1[19][46] = 16'b0000000000000101;
    assign weights1[19][47] = 16'b1111111111111101;
    assign weights1[19][48] = 16'b1111111111111101;
    assign weights1[19][49] = 16'b1111111111111010;
    assign weights1[19][50] = 16'b1111111111111000;
    assign weights1[19][51] = 16'b1111111111110110;
    assign weights1[19][52] = 16'b1111111111110001;
    assign weights1[19][53] = 16'b1111111111110010;
    assign weights1[19][54] = 16'b1111111111110111;
    assign weights1[19][55] = 16'b1111111111111011;
    assign weights1[19][56] = 16'b0000000000000000;
    assign weights1[19][57] = 16'b1111111111111111;
    assign weights1[19][58] = 16'b1111111111111010;
    assign weights1[19][59] = 16'b1111111111110100;
    assign weights1[19][60] = 16'b1111111111101001;
    assign weights1[19][61] = 16'b1111111111100010;
    assign weights1[19][62] = 16'b1111111111011010;
    assign weights1[19][63] = 16'b1111111111001110;
    assign weights1[19][64] = 16'b1111111111010000;
    assign weights1[19][65] = 16'b1111111111010101;
    assign weights1[19][66] = 16'b1111111111100000;
    assign weights1[19][67] = 16'b1111111111110011;
    assign weights1[19][68] = 16'b0000000000000100;
    assign weights1[19][69] = 16'b0000000000011101;
    assign weights1[19][70] = 16'b0000000000100111;
    assign weights1[19][71] = 16'b0000000000101001;
    assign weights1[19][72] = 16'b0000000000100110;
    assign weights1[19][73] = 16'b0000000000100001;
    assign weights1[19][74] = 16'b0000000000011111;
    assign weights1[19][75] = 16'b0000000000010000;
    assign weights1[19][76] = 16'b0000000000000011;
    assign weights1[19][77] = 16'b0000000000001011;
    assign weights1[19][78] = 16'b1111111111111100;
    assign weights1[19][79] = 16'b1111111111110000;
    assign weights1[19][80] = 16'b1111111111110100;
    assign weights1[19][81] = 16'b1111111111110001;
    assign weights1[19][82] = 16'b1111111111110101;
    assign weights1[19][83] = 16'b1111111111111001;
    assign weights1[19][84] = 16'b1111111111111101;
    assign weights1[19][85] = 16'b1111111111111101;
    assign weights1[19][86] = 16'b1111111111110110;
    assign weights1[19][87] = 16'b1111111111101000;
    assign weights1[19][88] = 16'b1111111111010111;
    assign weights1[19][89] = 16'b1111111111001001;
    assign weights1[19][90] = 16'b1111111111000000;
    assign weights1[19][91] = 16'b1111111110110010;
    assign weights1[19][92] = 16'b1111111111000101;
    assign weights1[19][93] = 16'b1111111110111000;
    assign weights1[19][94] = 16'b1111111111000001;
    assign weights1[19][95] = 16'b1111111111000101;
    assign weights1[19][96] = 16'b1111111111011000;
    assign weights1[19][97] = 16'b1111111111101000;
    assign weights1[19][98] = 16'b1111111111101000;
    assign weights1[19][99] = 16'b0000000000000010;
    assign weights1[19][100] = 16'b0000000000001010;
    assign weights1[19][101] = 16'b0000000000010110;
    assign weights1[19][102] = 16'b0000000000011001;
    assign weights1[19][103] = 16'b0000000000010011;
    assign weights1[19][104] = 16'b0000000000000110;
    assign weights1[19][105] = 16'b0000000000000110;
    assign weights1[19][106] = 16'b0000000000000111;
    assign weights1[19][107] = 16'b0000000000000001;
    assign weights1[19][108] = 16'b1111111111111100;
    assign weights1[19][109] = 16'b1111111111100110;
    assign weights1[19][110] = 16'b1111111111101001;
    assign weights1[19][111] = 16'b1111111111110110;
    assign weights1[19][112] = 16'b1111111111111110;
    assign weights1[19][113] = 16'b1111111111110110;
    assign weights1[19][114] = 16'b1111111111101001;
    assign weights1[19][115] = 16'b1111111111011110;
    assign weights1[19][116] = 16'b1111111111000111;
    assign weights1[19][117] = 16'b1111111110111011;
    assign weights1[19][118] = 16'b1111111110110000;
    assign weights1[19][119] = 16'b1111111110110001;
    assign weights1[19][120] = 16'b1111111110101100;
    assign weights1[19][121] = 16'b1111111110011001;
    assign weights1[19][122] = 16'b1111111110010110;
    assign weights1[19][123] = 16'b1111111110010010;
    assign weights1[19][124] = 16'b1111111110100000;
    assign weights1[19][125] = 16'b1111111110111111;
    assign weights1[19][126] = 16'b1111111111001001;
    assign weights1[19][127] = 16'b1111111111010011;
    assign weights1[19][128] = 16'b1111111111001010;
    assign weights1[19][129] = 16'b1111111111010111;
    assign weights1[19][130] = 16'b1111111111111000;
    assign weights1[19][131] = 16'b0000000000000010;
    assign weights1[19][132] = 16'b0000000000001000;
    assign weights1[19][133] = 16'b0000000000010001;
    assign weights1[19][134] = 16'b0000000000010101;
    assign weights1[19][135] = 16'b0000000000001100;
    assign weights1[19][136] = 16'b1111111111110011;
    assign weights1[19][137] = 16'b1111111111110000;
    assign weights1[19][138] = 16'b1111111111110010;
    assign weights1[19][139] = 16'b1111111111110101;
    assign weights1[19][140] = 16'b1111111111111100;
    assign weights1[19][141] = 16'b1111111111110101;
    assign weights1[19][142] = 16'b1111111111100111;
    assign weights1[19][143] = 16'b1111111111010001;
    assign weights1[19][144] = 16'b1111111110111111;
    assign weights1[19][145] = 16'b1111111111000010;
    assign weights1[19][146] = 16'b1111111111001101;
    assign weights1[19][147] = 16'b1111111110111011;
    assign weights1[19][148] = 16'b1111111110011111;
    assign weights1[19][149] = 16'b1111111110001101;
    assign weights1[19][150] = 16'b1111111101111001;
    assign weights1[19][151] = 16'b1111111110001011;
    assign weights1[19][152] = 16'b1111111101111111;
    assign weights1[19][153] = 16'b1111111110100010;
    assign weights1[19][154] = 16'b1111111111010010;
    assign weights1[19][155] = 16'b1111111111110101;
    assign weights1[19][156] = 16'b1111111111111011;
    assign weights1[19][157] = 16'b1111111111101110;
    assign weights1[19][158] = 16'b1111111111110111;
    assign weights1[19][159] = 16'b0000000000001000;
    assign weights1[19][160] = 16'b0000000000000000;
    assign weights1[19][161] = 16'b1111111111111010;
    assign weights1[19][162] = 16'b1111111111111101;
    assign weights1[19][163] = 16'b0000000000001011;
    assign weights1[19][164] = 16'b1111111111111010;
    assign weights1[19][165] = 16'b1111111111110011;
    assign weights1[19][166] = 16'b1111111111101000;
    assign weights1[19][167] = 16'b1111111111101100;
    assign weights1[19][168] = 16'b1111111111111100;
    assign weights1[19][169] = 16'b1111111111110100;
    assign weights1[19][170] = 16'b1111111111110000;
    assign weights1[19][171] = 16'b1111111111100000;
    assign weights1[19][172] = 16'b1111111111101110;
    assign weights1[19][173] = 16'b1111111111101110;
    assign weights1[19][174] = 16'b1111111111011010;
    assign weights1[19][175] = 16'b1111111111001000;
    assign weights1[19][176] = 16'b1111111111101010;
    assign weights1[19][177] = 16'b1111111111100101;
    assign weights1[19][178] = 16'b1111111111000010;
    assign weights1[19][179] = 16'b1111111111010111;
    assign weights1[19][180] = 16'b1111111111010000;
    assign weights1[19][181] = 16'b1111111111011010;
    assign weights1[19][182] = 16'b1111111111010101;
    assign weights1[19][183] = 16'b1111111111001111;
    assign weights1[19][184] = 16'b1111111111101110;
    assign weights1[19][185] = 16'b0000000000000000;
    assign weights1[19][186] = 16'b1111111111111000;
    assign weights1[19][187] = 16'b0000000000000110;
    assign weights1[19][188] = 16'b1111111111101010;
    assign weights1[19][189] = 16'b0000000000010110;
    assign weights1[19][190] = 16'b1111111111101110;
    assign weights1[19][191] = 16'b1111111111111011;
    assign weights1[19][192] = 16'b0000000000000101;
    assign weights1[19][193] = 16'b1111111111110101;
    assign weights1[19][194] = 16'b1111111111110100;
    assign weights1[19][195] = 16'b1111111111111000;
    assign weights1[19][196] = 16'b1111111111111110;
    assign weights1[19][197] = 16'b1111111111111111;
    assign weights1[19][198] = 16'b1111111111111100;
    assign weights1[19][199] = 16'b1111111111111000;
    assign weights1[19][200] = 16'b0000000000001100;
    assign weights1[19][201] = 16'b0000000000100100;
    assign weights1[19][202] = 16'b0000000000110011;
    assign weights1[19][203] = 16'b0000000000100000;
    assign weights1[19][204] = 16'b0000000000000010;
    assign weights1[19][205] = 16'b0000000000010111;
    assign weights1[19][206] = 16'b0000000000010111;
    assign weights1[19][207] = 16'b1111111111100100;
    assign weights1[19][208] = 16'b1111111111101100;
    assign weights1[19][209] = 16'b1111111111111110;
    assign weights1[19][210] = 16'b1111111111110011;
    assign weights1[19][211] = 16'b1111111111110001;
    assign weights1[19][212] = 16'b1111111111101001;
    assign weights1[19][213] = 16'b0000000000000011;
    assign weights1[19][214] = 16'b0000000000000110;
    assign weights1[19][215] = 16'b1111111111111001;
    assign weights1[19][216] = 16'b0000000000001110;
    assign weights1[19][217] = 16'b0000000000000111;
    assign weights1[19][218] = 16'b0000000000001001;
    assign weights1[19][219] = 16'b1111111111110010;
    assign weights1[19][220] = 16'b1111111111101011;
    assign weights1[19][221] = 16'b1111111111111010;
    assign weights1[19][222] = 16'b1111111111111100;
    assign weights1[19][223] = 16'b1111111111111010;
    assign weights1[19][224] = 16'b0000000000000110;
    assign weights1[19][225] = 16'b0000000000001010;
    assign weights1[19][226] = 16'b0000000000000110;
    assign weights1[19][227] = 16'b0000000000010111;
    assign weights1[19][228] = 16'b0000000001001010;
    assign weights1[19][229] = 16'b0000000000100110;
    assign weights1[19][230] = 16'b0000000000100101;
    assign weights1[19][231] = 16'b0000000000110101;
    assign weights1[19][232] = 16'b0000000001001001;
    assign weights1[19][233] = 16'b0000000000001101;
    assign weights1[19][234] = 16'b0000000000100110;
    assign weights1[19][235] = 16'b0000000000010001;
    assign weights1[19][236] = 16'b0000000000000110;
    assign weights1[19][237] = 16'b1111111111111100;
    assign weights1[19][238] = 16'b0000000000000000;
    assign weights1[19][239] = 16'b1111111111111100;
    assign weights1[19][240] = 16'b0000000000000010;
    assign weights1[19][241] = 16'b1111111111111111;
    assign weights1[19][242] = 16'b0000000000000000;
    assign weights1[19][243] = 16'b0000000000000000;
    assign weights1[19][244] = 16'b1111111111111010;
    assign weights1[19][245] = 16'b1111111111111100;
    assign weights1[19][246] = 16'b1111111111111111;
    assign weights1[19][247] = 16'b0000000000010000;
    assign weights1[19][248] = 16'b1111111111101001;
    assign weights1[19][249] = 16'b1111111111110110;
    assign weights1[19][250] = 16'b1111111111111111;
    assign weights1[19][251] = 16'b1111111111110000;
    assign weights1[19][252] = 16'b0000000000001100;
    assign weights1[19][253] = 16'b0000000000001010;
    assign weights1[19][254] = 16'b0000000000011001;
    assign weights1[19][255] = 16'b0000000000010110;
    assign weights1[19][256] = 16'b0000000000100000;
    assign weights1[19][257] = 16'b0000000000110110;
    assign weights1[19][258] = 16'b0000000000010011;
    assign weights1[19][259] = 16'b0000000000100100;
    assign weights1[19][260] = 16'b0000000000000000;
    assign weights1[19][261] = 16'b0000000000100101;
    assign weights1[19][262] = 16'b0000000000011101;
    assign weights1[19][263] = 16'b0000000000011000;
    assign weights1[19][264] = 16'b0000000000010100;
    assign weights1[19][265] = 16'b0000000000011101;
    assign weights1[19][266] = 16'b0000000000100010;
    assign weights1[19][267] = 16'b0000000000001010;
    assign weights1[19][268] = 16'b1111111111110001;
    assign weights1[19][269] = 16'b0000000000001001;
    assign weights1[19][270] = 16'b1111111111101001;
    assign weights1[19][271] = 16'b1111111111101110;
    assign weights1[19][272] = 16'b0000000000001110;
    assign weights1[19][273] = 16'b1111111111111100;
    assign weights1[19][274] = 16'b1111111111111101;
    assign weights1[19][275] = 16'b1111111111110101;
    assign weights1[19][276] = 16'b0000000000000010;
    assign weights1[19][277] = 16'b1111111111110111;
    assign weights1[19][278] = 16'b0000000000001000;
    assign weights1[19][279] = 16'b1111111111101000;
    assign weights1[19][280] = 16'b0000000000010011;
    assign weights1[19][281] = 16'b0000000000010111;
    assign weights1[19][282] = 16'b0000000000011011;
    assign weights1[19][283] = 16'b0000000000000100;
    assign weights1[19][284] = 16'b0000000000011111;
    assign weights1[19][285] = 16'b0000000000100000;
    assign weights1[19][286] = 16'b0000000000010111;
    assign weights1[19][287] = 16'b0000000000100110;
    assign weights1[19][288] = 16'b0000000000011001;
    assign weights1[19][289] = 16'b0000000000111010;
    assign weights1[19][290] = 16'b0000000000100110;
    assign weights1[19][291] = 16'b0000000000110001;
    assign weights1[19][292] = 16'b0000000000110101;
    assign weights1[19][293] = 16'b0000000000011011;
    assign weights1[19][294] = 16'b0000000000100010;
    assign weights1[19][295] = 16'b0000000000011000;
    assign weights1[19][296] = 16'b0000000000000110;
    assign weights1[19][297] = 16'b0000000000001111;
    assign weights1[19][298] = 16'b0000000000001000;
    assign weights1[19][299] = 16'b0000000000001001;
    assign weights1[19][300] = 16'b0000000000000001;
    assign weights1[19][301] = 16'b1111111111110101;
    assign weights1[19][302] = 16'b1111111111110111;
    assign weights1[19][303] = 16'b1111111111101001;
    assign weights1[19][304] = 16'b1111111111111100;
    assign weights1[19][305] = 16'b1111111111111100;
    assign weights1[19][306] = 16'b1111111111111011;
    assign weights1[19][307] = 16'b1111111111110110;
    assign weights1[19][308] = 16'b0000000000011010;
    assign weights1[19][309] = 16'b0000000000100010;
    assign weights1[19][310] = 16'b0000000000010010;
    assign weights1[19][311] = 16'b0000000000001011;
    assign weights1[19][312] = 16'b0000000000011111;
    assign weights1[19][313] = 16'b0000000000000111;
    assign weights1[19][314] = 16'b0000000000001101;
    assign weights1[19][315] = 16'b0000000000111000;
    assign weights1[19][316] = 16'b1111111111110110;
    assign weights1[19][317] = 16'b0000000000011011;
    assign weights1[19][318] = 16'b0000000000111111;
    assign weights1[19][319] = 16'b0000000000011111;
    assign weights1[19][320] = 16'b0000000000011101;
    assign weights1[19][321] = 16'b0000000000000001;
    assign weights1[19][322] = 16'b0000000000000011;
    assign weights1[19][323] = 16'b0000000000000011;
    assign weights1[19][324] = 16'b0000000000001100;
    assign weights1[19][325] = 16'b1111111111111010;
    assign weights1[19][326] = 16'b0000000000000011;
    assign weights1[19][327] = 16'b1111111111110111;
    assign weights1[19][328] = 16'b0000000000000011;
    assign weights1[19][329] = 16'b1111111111111011;
    assign weights1[19][330] = 16'b0000000000010000;
    assign weights1[19][331] = 16'b0000000000000000;
    assign weights1[19][332] = 16'b1111111111111101;
    assign weights1[19][333] = 16'b1111111111111111;
    assign weights1[19][334] = 16'b1111111111111110;
    assign weights1[19][335] = 16'b1111111111100100;
    assign weights1[19][336] = 16'b0000000000001111;
    assign weights1[19][337] = 16'b0000000000001111;
    assign weights1[19][338] = 16'b0000000000010001;
    assign weights1[19][339] = 16'b0000000000010101;
    assign weights1[19][340] = 16'b0000000000100101;
    assign weights1[19][341] = 16'b0000000000010001;
    assign weights1[19][342] = 16'b0000000000010101;
    assign weights1[19][343] = 16'b0000000000101111;
    assign weights1[19][344] = 16'b0000000000010110;
    assign weights1[19][345] = 16'b0000000000010110;
    assign weights1[19][346] = 16'b0000000000000010;
    assign weights1[19][347] = 16'b1111111111101100;
    assign weights1[19][348] = 16'b1111111111111010;
    assign weights1[19][349] = 16'b1111111111100110;
    assign weights1[19][350] = 16'b1111111111101111;
    assign weights1[19][351] = 16'b1111111111110001;
    assign weights1[19][352] = 16'b1111111111011111;
    assign weights1[19][353] = 16'b0000000000001101;
    assign weights1[19][354] = 16'b1111111111111011;
    assign weights1[19][355] = 16'b0000000000011011;
    assign weights1[19][356] = 16'b1111111111111100;
    assign weights1[19][357] = 16'b0000000000000001;
    assign weights1[19][358] = 16'b0000000000010000;
    assign weights1[19][359] = 16'b1111111111101110;
    assign weights1[19][360] = 16'b1111111111110111;
    assign weights1[19][361] = 16'b0000000000010011;
    assign weights1[19][362] = 16'b0000000000001010;
    assign weights1[19][363] = 16'b1111111111110111;
    assign weights1[19][364] = 16'b0000000000001010;
    assign weights1[19][365] = 16'b1111111111111001;
    assign weights1[19][366] = 16'b0000000000010010;
    assign weights1[19][367] = 16'b0000000000010111;
    assign weights1[19][368] = 16'b0000000000001011;
    assign weights1[19][369] = 16'b0000000000001111;
    assign weights1[19][370] = 16'b0000000000011010;
    assign weights1[19][371] = 16'b0000000000001011;
    assign weights1[19][372] = 16'b0000000000000111;
    assign weights1[19][373] = 16'b1111111111010001;
    assign weights1[19][374] = 16'b1111111110111011;
    assign weights1[19][375] = 16'b1111111110101001;
    assign weights1[19][376] = 16'b1111111110100000;
    assign weights1[19][377] = 16'b1111111111000010;
    assign weights1[19][378] = 16'b1111111111010100;
    assign weights1[19][379] = 16'b1111111111100100;
    assign weights1[19][380] = 16'b1111111111110101;
    assign weights1[19][381] = 16'b1111111111111110;
    assign weights1[19][382] = 16'b1111111111111111;
    assign weights1[19][383] = 16'b1111111111101011;
    assign weights1[19][384] = 16'b1111111111111010;
    assign weights1[19][385] = 16'b1111111111111000;
    assign weights1[19][386] = 16'b0000000000000010;
    assign weights1[19][387] = 16'b0000000000001000;
    assign weights1[19][388] = 16'b0000000000001000;
    assign weights1[19][389] = 16'b1111111111110001;
    assign weights1[19][390] = 16'b0000000000010011;
    assign weights1[19][391] = 16'b1111111111101010;
    assign weights1[19][392] = 16'b1111111111101011;
    assign weights1[19][393] = 16'b1111111111011000;
    assign weights1[19][394] = 16'b1111111111101101;
    assign weights1[19][395] = 16'b1111111111111000;
    assign weights1[19][396] = 16'b1111111111111111;
    assign weights1[19][397] = 16'b0000000000000001;
    assign weights1[19][398] = 16'b1111111111000110;
    assign weights1[19][399] = 16'b1111111110110011;
    assign weights1[19][400] = 16'b1111111101111101;
    assign weights1[19][401] = 16'b1111111100011110;
    assign weights1[19][402] = 16'b1111111101111100;
    assign weights1[19][403] = 16'b1111111110011110;
    assign weights1[19][404] = 16'b1111111111011001;
    assign weights1[19][405] = 16'b1111111111001101;
    assign weights1[19][406] = 16'b1111111111100101;
    assign weights1[19][407] = 16'b1111111111111000;
    assign weights1[19][408] = 16'b1111111111111000;
    assign weights1[19][409] = 16'b1111111111111110;
    assign weights1[19][410] = 16'b1111111111101110;
    assign weights1[19][411] = 16'b0000000000000010;
    assign weights1[19][412] = 16'b1111111111111000;
    assign weights1[19][413] = 16'b1111111111111111;
    assign weights1[19][414] = 16'b1111111111110110;
    assign weights1[19][415] = 16'b0000000000011000;
    assign weights1[19][416] = 16'b1111111111101001;
    assign weights1[19][417] = 16'b1111111111111100;
    assign weights1[19][418] = 16'b1111111111111111;
    assign weights1[19][419] = 16'b1111111111110111;
    assign weights1[19][420] = 16'b1111111111011001;
    assign weights1[19][421] = 16'b1111111110111101;
    assign weights1[19][422] = 16'b1111111111000010;
    assign weights1[19][423] = 16'b1111111110111111;
    assign weights1[19][424] = 16'b1111111110100100;
    assign weights1[19][425] = 16'b1111111110011001;
    assign weights1[19][426] = 16'b1111111101100100;
    assign weights1[19][427] = 16'b1111111100000110;
    assign weights1[19][428] = 16'b1111111100010011;
    assign weights1[19][429] = 16'b1111111110000111;
    assign weights1[19][430] = 16'b1111111111011101;
    assign weights1[19][431] = 16'b0000000000000000;
    assign weights1[19][432] = 16'b0000000000000000;
    assign weights1[19][433] = 16'b0000000000000110;
    assign weights1[19][434] = 16'b0000000000001110;
    assign weights1[19][435] = 16'b0000000000000111;
    assign weights1[19][436] = 16'b0000000000001101;
    assign weights1[19][437] = 16'b0000000000010001;
    assign weights1[19][438] = 16'b0000000000000101;
    assign weights1[19][439] = 16'b0000000000000000;
    assign weights1[19][440] = 16'b0000000000011010;
    assign weights1[19][441] = 16'b0000000000010001;
    assign weights1[19][442] = 16'b0000000000000100;
    assign weights1[19][443] = 16'b0000000000001111;
    assign weights1[19][444] = 16'b0000000000001001;
    assign weights1[19][445] = 16'b0000000000000010;
    assign weights1[19][446] = 16'b0000000000000011;
    assign weights1[19][447] = 16'b0000000000000101;
    assign weights1[19][448] = 16'b1111111111000001;
    assign weights1[19][449] = 16'b1111111110110100;
    assign weights1[19][450] = 16'b1111111110101011;
    assign weights1[19][451] = 16'b1111111110001111;
    assign weights1[19][452] = 16'b1111111101010110;
    assign weights1[19][453] = 16'b1111111100111001;
    assign weights1[19][454] = 16'b1111111100100010;
    assign weights1[19][455] = 16'b1111111101010101;
    assign weights1[19][456] = 16'b1111111111110010;
    assign weights1[19][457] = 16'b0000000000010100;
    assign weights1[19][458] = 16'b0000000000001101;
    assign weights1[19][459] = 16'b0000000000001110;
    assign weights1[19][460] = 16'b0000000000100000;
    assign weights1[19][461] = 16'b0000000000001010;
    assign weights1[19][462] = 16'b0000000000000001;
    assign weights1[19][463] = 16'b0000000000000011;
    assign weights1[19][464] = 16'b0000000000010011;
    assign weights1[19][465] = 16'b0000000000010001;
    assign weights1[19][466] = 16'b0000000000010000;
    assign weights1[19][467] = 16'b0000000000000010;
    assign weights1[19][468] = 16'b0000000000000011;
    assign weights1[19][469] = 16'b0000000000000000;
    assign weights1[19][470] = 16'b0000000000001010;
    assign weights1[19][471] = 16'b0000000000000011;
    assign weights1[19][472] = 16'b1111111111111111;
    assign weights1[19][473] = 16'b0000000000011000;
    assign weights1[19][474] = 16'b1111111111111001;
    assign weights1[19][475] = 16'b0000000000000101;
    assign weights1[19][476] = 16'b1111111110111110;
    assign weights1[19][477] = 16'b1111111110110100;
    assign weights1[19][478] = 16'b1111111110100001;
    assign weights1[19][479] = 16'b1111111110001100;
    assign weights1[19][480] = 16'b1111111110000010;
    assign weights1[19][481] = 16'b1111111110010110;
    assign weights1[19][482] = 16'b1111111110101001;
    assign weights1[19][483] = 16'b0000000000001011;
    assign weights1[19][484] = 16'b0000000000000111;
    assign weights1[19][485] = 16'b0000000000011001;
    assign weights1[19][486] = 16'b0000000000010100;
    assign weights1[19][487] = 16'b0000000000011011;
    assign weights1[19][488] = 16'b0000000000001101;
    assign weights1[19][489] = 16'b0000000000001110;
    assign weights1[19][490] = 16'b0000000000001101;
    assign weights1[19][491] = 16'b0000000000000000;
    assign weights1[19][492] = 16'b1111111111111000;
    assign weights1[19][493] = 16'b0000000000000000;
    assign weights1[19][494] = 16'b0000000000001100;
    assign weights1[19][495] = 16'b0000000000000000;
    assign weights1[19][496] = 16'b0000000000011111;
    assign weights1[19][497] = 16'b1111111111111111;
    assign weights1[19][498] = 16'b1111111111110110;
    assign weights1[19][499] = 16'b0000000000001000;
    assign weights1[19][500] = 16'b0000000000000101;
    assign weights1[19][501] = 16'b1111111111111010;
    assign weights1[19][502] = 16'b1111111111110001;
    assign weights1[19][503] = 16'b1111111111110100;
    assign weights1[19][504] = 16'b1111111111000101;
    assign weights1[19][505] = 16'b1111111110111100;
    assign weights1[19][506] = 16'b1111111110101001;
    assign weights1[19][507] = 16'b1111111110101001;
    assign weights1[19][508] = 16'b1111111111001100;
    assign weights1[19][509] = 16'b1111111111110010;
    assign weights1[19][510] = 16'b0000000000000100;
    assign weights1[19][511] = 16'b0000000000101010;
    assign weights1[19][512] = 16'b0000000000110000;
    assign weights1[19][513] = 16'b0000000000001100;
    assign weights1[19][514] = 16'b0000000000011001;
    assign weights1[19][515] = 16'b0000000000010001;
    assign weights1[19][516] = 16'b1111111111111011;
    assign weights1[19][517] = 16'b0000000000000010;
    assign weights1[19][518] = 16'b0000000000000100;
    assign weights1[19][519] = 16'b0000000000001110;
    assign weights1[19][520] = 16'b0000000000000010;
    assign weights1[19][521] = 16'b1111111111111010;
    assign weights1[19][522] = 16'b1111111111111111;
    assign weights1[19][523] = 16'b0000000000000100;
    assign weights1[19][524] = 16'b0000000000000010;
    assign weights1[19][525] = 16'b0000000000000011;
    assign weights1[19][526] = 16'b0000000000001111;
    assign weights1[19][527] = 16'b1111111111110110;
    assign weights1[19][528] = 16'b1111111111110000;
    assign weights1[19][529] = 16'b1111111111111011;
    assign weights1[19][530] = 16'b0000000000001001;
    assign weights1[19][531] = 16'b0000000000100000;
    assign weights1[19][532] = 16'b1111111111010111;
    assign weights1[19][533] = 16'b1111111111010001;
    assign weights1[19][534] = 16'b1111111111001110;
    assign weights1[19][535] = 16'b1111111111001111;
    assign weights1[19][536] = 16'b1111111111101111;
    assign weights1[19][537] = 16'b0000000000100000;
    assign weights1[19][538] = 16'b0000000000000101;
    assign weights1[19][539] = 16'b0000000000010001;
    assign weights1[19][540] = 16'b0000000000000011;
    assign weights1[19][541] = 16'b0000000000000000;
    assign weights1[19][542] = 16'b1111111111111100;
    assign weights1[19][543] = 16'b1111111111111100;
    assign weights1[19][544] = 16'b0000000000000111;
    assign weights1[19][545] = 16'b1111111111111001;
    assign weights1[19][546] = 16'b0000000000000111;
    assign weights1[19][547] = 16'b0000000000000011;
    assign weights1[19][548] = 16'b0000000000001011;
    assign weights1[19][549] = 16'b1111111111111101;
    assign weights1[19][550] = 16'b1111111111101011;
    assign weights1[19][551] = 16'b0000000000000101;
    assign weights1[19][552] = 16'b0000000000000000;
    assign weights1[19][553] = 16'b0000000000000010;
    assign weights1[19][554] = 16'b0000000000000011;
    assign weights1[19][555] = 16'b0000000000010100;
    assign weights1[19][556] = 16'b1111111111111010;
    assign weights1[19][557] = 16'b1111111111111111;
    assign weights1[19][558] = 16'b1111111111111111;
    assign weights1[19][559] = 16'b0000000000010110;
    assign weights1[19][560] = 16'b1111111111101111;
    assign weights1[19][561] = 16'b1111111111101011;
    assign weights1[19][562] = 16'b1111111111111001;
    assign weights1[19][563] = 16'b1111111111111011;
    assign weights1[19][564] = 16'b0000000000100001;
    assign weights1[19][565] = 16'b1111111111111001;
    assign weights1[19][566] = 16'b1111111111101010;
    assign weights1[19][567] = 16'b1111111111111100;
    assign weights1[19][568] = 16'b0000000000001000;
    assign weights1[19][569] = 16'b0000000000010101;
    assign weights1[19][570] = 16'b1111111111101101;
    assign weights1[19][571] = 16'b0000000000001100;
    assign weights1[19][572] = 16'b1111111111111001;
    assign weights1[19][573] = 16'b1111111111111101;
    assign weights1[19][574] = 16'b0000000000000010;
    assign weights1[19][575] = 16'b1111111111111001;
    assign weights1[19][576] = 16'b0000000000000001;
    assign weights1[19][577] = 16'b1111111111111101;
    assign weights1[19][578] = 16'b0000000000001110;
    assign weights1[19][579] = 16'b0000000000000110;
    assign weights1[19][580] = 16'b1111111111111110;
    assign weights1[19][581] = 16'b1111111111110011;
    assign weights1[19][582] = 16'b0000000000000110;
    assign weights1[19][583] = 16'b0000000000000101;
    assign weights1[19][584] = 16'b1111111111111111;
    assign weights1[19][585] = 16'b1111111111111001;
    assign weights1[19][586] = 16'b1111111111111111;
    assign weights1[19][587] = 16'b0000000000000001;
    assign weights1[19][588] = 16'b1111111111111010;
    assign weights1[19][589] = 16'b1111111111111100;
    assign weights1[19][590] = 16'b0000000000001111;
    assign weights1[19][591] = 16'b0000000000001011;
    assign weights1[19][592] = 16'b0000000000000011;
    assign weights1[19][593] = 16'b1111111111111101;
    assign weights1[19][594] = 16'b1111111111111011;
    assign weights1[19][595] = 16'b0000000000000100;
    assign weights1[19][596] = 16'b1111111111111010;
    assign weights1[19][597] = 16'b1111111111110110;
    assign weights1[19][598] = 16'b0000000000010000;
    assign weights1[19][599] = 16'b1111111111101000;
    assign weights1[19][600] = 16'b0000000000010000;
    assign weights1[19][601] = 16'b0000000000000001;
    assign weights1[19][602] = 16'b0000000000000001;
    assign weights1[19][603] = 16'b1111111111111011;
    assign weights1[19][604] = 16'b1111111111111101;
    assign weights1[19][605] = 16'b1111111111110001;
    assign weights1[19][606] = 16'b1111111111111001;
    assign weights1[19][607] = 16'b1111111111111000;
    assign weights1[19][608] = 16'b1111111111111100;
    assign weights1[19][609] = 16'b1111111111111000;
    assign weights1[19][610] = 16'b0000000000000000;
    assign weights1[19][611] = 16'b0000000000001000;
    assign weights1[19][612] = 16'b1111111111111010;
    assign weights1[19][613] = 16'b0000000000000101;
    assign weights1[19][614] = 16'b1111111111111011;
    assign weights1[19][615] = 16'b1111111111111110;
    assign weights1[19][616] = 16'b0000000000001001;
    assign weights1[19][617] = 16'b1111111111111111;
    assign weights1[19][618] = 16'b0000000000001110;
    assign weights1[19][619] = 16'b0000000000010001;
    assign weights1[19][620] = 16'b0000000000001010;
    assign weights1[19][621] = 16'b1111111111111011;
    assign weights1[19][622] = 16'b0000000000011100;
    assign weights1[19][623] = 16'b1111111111111011;
    assign weights1[19][624] = 16'b1111111111111111;
    assign weights1[19][625] = 16'b1111111111111111;
    assign weights1[19][626] = 16'b0000000000011011;
    assign weights1[19][627] = 16'b1111111111110011;
    assign weights1[19][628] = 16'b0000000000000110;
    assign weights1[19][629] = 16'b1111111111111010;
    assign weights1[19][630] = 16'b1111111111111000;
    assign weights1[19][631] = 16'b1111111111110000;
    assign weights1[19][632] = 16'b1111111111110001;
    assign weights1[19][633] = 16'b0000000000001010;
    assign weights1[19][634] = 16'b1111111111101100;
    assign weights1[19][635] = 16'b0000000000001001;
    assign weights1[19][636] = 16'b0000000000001001;
    assign weights1[19][637] = 16'b1111111111111100;
    assign weights1[19][638] = 16'b0000000000000101;
    assign weights1[19][639] = 16'b0000000000000001;
    assign weights1[19][640] = 16'b1111111111111101;
    assign weights1[19][641] = 16'b1111111111111110;
    assign weights1[19][642] = 16'b0000000000000001;
    assign weights1[19][643] = 16'b0000000000000011;
    assign weights1[19][644] = 16'b0000000000000011;
    assign weights1[19][645] = 16'b0000000000000001;
    assign weights1[19][646] = 16'b0000000000010001;
    assign weights1[19][647] = 16'b0000000000001100;
    assign weights1[19][648] = 16'b1111111111111110;
    assign weights1[19][649] = 16'b0000000000011010;
    assign weights1[19][650] = 16'b0000000000010010;
    assign weights1[19][651] = 16'b0000000000011100;
    assign weights1[19][652] = 16'b1111111111111100;
    assign weights1[19][653] = 16'b0000000000000101;
    assign weights1[19][654] = 16'b1111111111111110;
    assign weights1[19][655] = 16'b0000000000001011;
    assign weights1[19][656] = 16'b0000000000000000;
    assign weights1[19][657] = 16'b1111111111110111;
    assign weights1[19][658] = 16'b0000000000000010;
    assign weights1[19][659] = 16'b0000000000010000;
    assign weights1[19][660] = 16'b0000000000000110;
    assign weights1[19][661] = 16'b1111111111110110;
    assign weights1[19][662] = 16'b0000000000010100;
    assign weights1[19][663] = 16'b1111111111101111;
    assign weights1[19][664] = 16'b0000000000000111;
    assign weights1[19][665] = 16'b1111111111110100;
    assign weights1[19][666] = 16'b0000000000000001;
    assign weights1[19][667] = 16'b0000000000000111;
    assign weights1[19][668] = 16'b0000000000000001;
    assign weights1[19][669] = 16'b1111111111111011;
    assign weights1[19][670] = 16'b1111111111111101;
    assign weights1[19][671] = 16'b0000000000000111;
    assign weights1[19][672] = 16'b0000000000000001;
    assign weights1[19][673] = 16'b0000000000000011;
    assign weights1[19][674] = 16'b0000000000001110;
    assign weights1[19][675] = 16'b0000000000000101;
    assign weights1[19][676] = 16'b0000000000000001;
    assign weights1[19][677] = 16'b0000000000001001;
    assign weights1[19][678] = 16'b1111111111101110;
    assign weights1[19][679] = 16'b0000000000001100;
    assign weights1[19][680] = 16'b1111111111011010;
    assign weights1[19][681] = 16'b0000000000011100;
    assign weights1[19][682] = 16'b1111111111111111;
    assign weights1[19][683] = 16'b0000000000010110;
    assign weights1[19][684] = 16'b0000000000000110;
    assign weights1[19][685] = 16'b1111111111110110;
    assign weights1[19][686] = 16'b0000000000010110;
    assign weights1[19][687] = 16'b0000000000000001;
    assign weights1[19][688] = 16'b1111111111111111;
    assign weights1[19][689] = 16'b0000000000001110;
    assign weights1[19][690] = 16'b0000000000001010;
    assign weights1[19][691] = 16'b1111111111111111;
    assign weights1[19][692] = 16'b0000000000000010;
    assign weights1[19][693] = 16'b0000000000001011;
    assign weights1[19][694] = 16'b1111111111111010;
    assign weights1[19][695] = 16'b1111111111110010;
    assign weights1[19][696] = 16'b1111111111110111;
    assign weights1[19][697] = 16'b0000000000000000;
    assign weights1[19][698] = 16'b1111111111110001;
    assign weights1[19][699] = 16'b0000000000000001;
    assign weights1[19][700] = 16'b1111111111111111;
    assign weights1[19][701] = 16'b0000000000000011;
    assign weights1[19][702] = 16'b0000000000001100;
    assign weights1[19][703] = 16'b1111111111111000;
    assign weights1[19][704] = 16'b0000000000000110;
    assign weights1[19][705] = 16'b1111111111110011;
    assign weights1[19][706] = 16'b1111111111110011;
    assign weights1[19][707] = 16'b0000000000000101;
    assign weights1[19][708] = 16'b0000000000010010;
    assign weights1[19][709] = 16'b0000000000001011;
    assign weights1[19][710] = 16'b1111111111010110;
    assign weights1[19][711] = 16'b1111111111111000;
    assign weights1[19][712] = 16'b0000000000000111;
    assign weights1[19][713] = 16'b0000000000001100;
    assign weights1[19][714] = 16'b0000000000001100;
    assign weights1[19][715] = 16'b1111111111110010;
    assign weights1[19][716] = 16'b0000000000000010;
    assign weights1[19][717] = 16'b1111111111111000;
    assign weights1[19][718] = 16'b0000000000000101;
    assign weights1[19][719] = 16'b1111111111111100;
    assign weights1[19][720] = 16'b0000000000010010;
    assign weights1[19][721] = 16'b1111111111111111;
    assign weights1[19][722] = 16'b0000000000000000;
    assign weights1[19][723] = 16'b1111111111111001;
    assign weights1[19][724] = 16'b1111111111101101;
    assign weights1[19][725] = 16'b1111111111110110;
    assign weights1[19][726] = 16'b1111111111110000;
    assign weights1[19][727] = 16'b0000000000000011;
    assign weights1[19][728] = 16'b0000000000000010;
    assign weights1[19][729] = 16'b1111111111111110;
    assign weights1[19][730] = 16'b0000000000001000;
    assign weights1[19][731] = 16'b1111111111111100;
    assign weights1[19][732] = 16'b1111111111111011;
    assign weights1[19][733] = 16'b1111111111011110;
    assign weights1[19][734] = 16'b1111111111110100;
    assign weights1[19][735] = 16'b0000000000001011;
    assign weights1[19][736] = 16'b0000000000000000;
    assign weights1[19][737] = 16'b0000000000000101;
    assign weights1[19][738] = 16'b0000000000010001;
    assign weights1[19][739] = 16'b0000000000000011;
    assign weights1[19][740] = 16'b0000000000001000;
    assign weights1[19][741] = 16'b1111111111110111;
    assign weights1[19][742] = 16'b0000000000000001;
    assign weights1[19][743] = 16'b1111111111111101;
    assign weights1[19][744] = 16'b1111111111111000;
    assign weights1[19][745] = 16'b1111111111111110;
    assign weights1[19][746] = 16'b1111111111101011;
    assign weights1[19][747] = 16'b0000000000000011;
    assign weights1[19][748] = 16'b1111111111111000;
    assign weights1[19][749] = 16'b0000000000001001;
    assign weights1[19][750] = 16'b0000000000000101;
    assign weights1[19][751] = 16'b1111111111111110;
    assign weights1[19][752] = 16'b1111111111110101;
    assign weights1[19][753] = 16'b1111111111111101;
    assign weights1[19][754] = 16'b0000000000000001;
    assign weights1[19][755] = 16'b0000000000000001;
    assign weights1[19][756] = 16'b0000000000000010;
    assign weights1[19][757] = 16'b1111111111111111;
    assign weights1[19][758] = 16'b0000000000001010;
    assign weights1[19][759] = 16'b0000000000010001;
    assign weights1[19][760] = 16'b0000000000001110;
    assign weights1[19][761] = 16'b0000000000000011;
    assign weights1[19][762] = 16'b0000000000001111;
    assign weights1[19][763] = 16'b0000000000001101;
    assign weights1[19][764] = 16'b0000000000000111;
    assign weights1[19][765] = 16'b1111111111111011;
    assign weights1[19][766] = 16'b0000000000001000;
    assign weights1[19][767] = 16'b0000000000001010;
    assign weights1[19][768] = 16'b1111111111111001;
    assign weights1[19][769] = 16'b0000000000001001;
    assign weights1[19][770] = 16'b0000000000000010;
    assign weights1[19][771] = 16'b1111111111111011;
    assign weights1[19][772] = 16'b1111111111111111;
    assign weights1[19][773] = 16'b0000000000010100;
    assign weights1[19][774] = 16'b1111111111110011;
    assign weights1[19][775] = 16'b1111111111110111;
    assign weights1[19][776] = 16'b1111111111111001;
    assign weights1[19][777] = 16'b1111111111111001;
    assign weights1[19][778] = 16'b1111111111110000;
    assign weights1[19][779] = 16'b1111111111111110;
    assign weights1[19][780] = 16'b1111111111111011;
    assign weights1[19][781] = 16'b1111111111111110;
    assign weights1[19][782] = 16'b0000000000000011;
    assign weights1[19][783] = 16'b0000000000000011;
    assign weights1[20][0] = 16'b0000000000000000;
    assign weights1[20][1] = 16'b0000000000000000;
    assign weights1[20][2] = 16'b0000000000000000;
    assign weights1[20][3] = 16'b0000000000000000;
    assign weights1[20][4] = 16'b0000000000000000;
    assign weights1[20][5] = 16'b1111111111111111;
    assign weights1[20][6] = 16'b1111111111111101;
    assign weights1[20][7] = 16'b1111111111111101;
    assign weights1[20][8] = 16'b1111111111111101;
    assign weights1[20][9] = 16'b1111111111111010;
    assign weights1[20][10] = 16'b1111111111111011;
    assign weights1[20][11] = 16'b1111111111110101;
    assign weights1[20][12] = 16'b1111111111101110;
    assign weights1[20][13] = 16'b1111111111110010;
    assign weights1[20][14] = 16'b1111111111110100;
    assign weights1[20][15] = 16'b1111111111110110;
    assign weights1[20][16] = 16'b1111111111110110;
    assign weights1[20][17] = 16'b1111111111110011;
    assign weights1[20][18] = 16'b1111111111110110;
    assign weights1[20][19] = 16'b1111111111110110;
    assign weights1[20][20] = 16'b1111111111111011;
    assign weights1[20][21] = 16'b1111111111111011;
    assign weights1[20][22] = 16'b1111111111111101;
    assign weights1[20][23] = 16'b1111111111111111;
    assign weights1[20][24] = 16'b1111111111111110;
    assign weights1[20][25] = 16'b0000000000000000;
    assign weights1[20][26] = 16'b0000000000000000;
    assign weights1[20][27] = 16'b0000000000000000;
    assign weights1[20][28] = 16'b0000000000000000;
    assign weights1[20][29] = 16'b0000000000000000;
    assign weights1[20][30] = 16'b0000000000000000;
    assign weights1[20][31] = 16'b1111111111111110;
    assign weights1[20][32] = 16'b1111111111111110;
    assign weights1[20][33] = 16'b1111111111111010;
    assign weights1[20][34] = 16'b1111111111111000;
    assign weights1[20][35] = 16'b1111111111111001;
    assign weights1[20][36] = 16'b1111111111111000;
    assign weights1[20][37] = 16'b1111111111110101;
    assign weights1[20][38] = 16'b1111111111101101;
    assign weights1[20][39] = 16'b1111111111110000;
    assign weights1[20][40] = 16'b1111111111101110;
    assign weights1[20][41] = 16'b1111111111101110;
    assign weights1[20][42] = 16'b1111111111101101;
    assign weights1[20][43] = 16'b1111111111110001;
    assign weights1[20][44] = 16'b1111111111101100;
    assign weights1[20][45] = 16'b1111111111101110;
    assign weights1[20][46] = 16'b1111111111101101;
    assign weights1[20][47] = 16'b1111111111101111;
    assign weights1[20][48] = 16'b1111111111101110;
    assign weights1[20][49] = 16'b1111111111100101;
    assign weights1[20][50] = 16'b1111111111101100;
    assign weights1[20][51] = 16'b1111111111110111;
    assign weights1[20][52] = 16'b1111111111111110;
    assign weights1[20][53] = 16'b1111111111111111;
    assign weights1[20][54] = 16'b0000000000000001;
    assign weights1[20][55] = 16'b0000000000000000;
    assign weights1[20][56] = 16'b0000000000000000;
    assign weights1[20][57] = 16'b0000000000000000;
    assign weights1[20][58] = 16'b0000000000000000;
    assign weights1[20][59] = 16'b1111111111111101;
    assign weights1[20][60] = 16'b1111111111111010;
    assign weights1[20][61] = 16'b1111111111110101;
    assign weights1[20][62] = 16'b1111111111110101;
    assign weights1[20][63] = 16'b1111111111110010;
    assign weights1[20][64] = 16'b1111111111101110;
    assign weights1[20][65] = 16'b1111111111101110;
    assign weights1[20][66] = 16'b1111111111100011;
    assign weights1[20][67] = 16'b1111111111100101;
    assign weights1[20][68] = 16'b1111111111100101;
    assign weights1[20][69] = 16'b1111111111100100;
    assign weights1[20][70] = 16'b1111111111100100;
    assign weights1[20][71] = 16'b1111111111100111;
    assign weights1[20][72] = 16'b1111111111011110;
    assign weights1[20][73] = 16'b1111111111100010;
    assign weights1[20][74] = 16'b1111111111011111;
    assign weights1[20][75] = 16'b1111111111100111;
    assign weights1[20][76] = 16'b1111111111100101;
    assign weights1[20][77] = 16'b1111111111100101;
    assign weights1[20][78] = 16'b1111111111100000;
    assign weights1[20][79] = 16'b1111111111101111;
    assign weights1[20][80] = 16'b1111111111110101;
    assign weights1[20][81] = 16'b1111111111111011;
    assign weights1[20][82] = 16'b1111111111111100;
    assign weights1[20][83] = 16'b1111111111111110;
    assign weights1[20][84] = 16'b0000000000000000;
    assign weights1[20][85] = 16'b0000000000000000;
    assign weights1[20][86] = 16'b1111111111111100;
    assign weights1[20][87] = 16'b1111111111111001;
    assign weights1[20][88] = 16'b1111111111110100;
    assign weights1[20][89] = 16'b1111111111110000;
    assign weights1[20][90] = 16'b1111111111100011;
    assign weights1[20][91] = 16'b1111111111100011;
    assign weights1[20][92] = 16'b1111111111011111;
    assign weights1[20][93] = 16'b1111111111011000;
    assign weights1[20][94] = 16'b1111111111011000;
    assign weights1[20][95] = 16'b1111111111100001;
    assign weights1[20][96] = 16'b1111111111011100;
    assign weights1[20][97] = 16'b1111111111011001;
    assign weights1[20][98] = 16'b1111111111011101;
    assign weights1[20][99] = 16'b1111111111011100;
    assign weights1[20][100] = 16'b1111111111011100;
    assign weights1[20][101] = 16'b1111111111011010;
    assign weights1[20][102] = 16'b1111111111100101;
    assign weights1[20][103] = 16'b1111111111100010;
    assign weights1[20][104] = 16'b1111111111011110;
    assign weights1[20][105] = 16'b1111111111011000;
    assign weights1[20][106] = 16'b1111111111100110;
    assign weights1[20][107] = 16'b1111111111101011;
    assign weights1[20][108] = 16'b1111111111110000;
    assign weights1[20][109] = 16'b1111111111110101;
    assign weights1[20][110] = 16'b1111111111111001;
    assign weights1[20][111] = 16'b1111111111111110;
    assign weights1[20][112] = 16'b0000000000000000;
    assign weights1[20][113] = 16'b1111111111111110;
    assign weights1[20][114] = 16'b1111111111110101;
    assign weights1[20][115] = 16'b1111111111101110;
    assign weights1[20][116] = 16'b1111111111101000;
    assign weights1[20][117] = 16'b1111111111100001;
    assign weights1[20][118] = 16'b1111111111100000;
    assign weights1[20][119] = 16'b1111111111011100;
    assign weights1[20][120] = 16'b1111111111011011;
    assign weights1[20][121] = 16'b1111111111001101;
    assign weights1[20][122] = 16'b1111111111010101;
    assign weights1[20][123] = 16'b1111111111010111;
    assign weights1[20][124] = 16'b1111111111010110;
    assign weights1[20][125] = 16'b1111111111010100;
    assign weights1[20][126] = 16'b1111111111001111;
    assign weights1[20][127] = 16'b1111111111010011;
    assign weights1[20][128] = 16'b1111111111010101;
    assign weights1[20][129] = 16'b1111111111010111;
    assign weights1[20][130] = 16'b1111111111011101;
    assign weights1[20][131] = 16'b1111111111100011;
    assign weights1[20][132] = 16'b1111111111011000;
    assign weights1[20][133] = 16'b1111111111010011;
    assign weights1[20][134] = 16'b1111111111011011;
    assign weights1[20][135] = 16'b1111111111101000;
    assign weights1[20][136] = 16'b1111111111101100;
    assign weights1[20][137] = 16'b1111111111101101;
    assign weights1[20][138] = 16'b1111111111110001;
    assign weights1[20][139] = 16'b1111111111110110;
    assign weights1[20][140] = 16'b0000000000000001;
    assign weights1[20][141] = 16'b1111111111111001;
    assign weights1[20][142] = 16'b1111111111101011;
    assign weights1[20][143] = 16'b1111111111011101;
    assign weights1[20][144] = 16'b1111111111010011;
    assign weights1[20][145] = 16'b1111111111001100;
    assign weights1[20][146] = 16'b1111111111001010;
    assign weights1[20][147] = 16'b1111111111000110;
    assign weights1[20][148] = 16'b1111111111000000;
    assign weights1[20][149] = 16'b1111111110110001;
    assign weights1[20][150] = 16'b1111111111000001;
    assign weights1[20][151] = 16'b1111111111001101;
    assign weights1[20][152] = 16'b1111111111000111;
    assign weights1[20][153] = 16'b1111111111001100;
    assign weights1[20][154] = 16'b1111111111001111;
    assign weights1[20][155] = 16'b1111111111001110;
    assign weights1[20][156] = 16'b1111111111000100;
    assign weights1[20][157] = 16'b1111111111001010;
    assign weights1[20][158] = 16'b1111111111010011;
    assign weights1[20][159] = 16'b1111111111010011;
    assign weights1[20][160] = 16'b1111111111001001;
    assign weights1[20][161] = 16'b1111111111001000;
    assign weights1[20][162] = 16'b1111111111011000;
    assign weights1[20][163] = 16'b1111111111011101;
    assign weights1[20][164] = 16'b1111111111011111;
    assign weights1[20][165] = 16'b1111111111101001;
    assign weights1[20][166] = 16'b1111111111101011;
    assign weights1[20][167] = 16'b1111111111110001;
    assign weights1[20][168] = 16'b1111111111111110;
    assign weights1[20][169] = 16'b1111111111110110;
    assign weights1[20][170] = 16'b1111111111101101;
    assign weights1[20][171] = 16'b1111111111010101;
    assign weights1[20][172] = 16'b1111111111000010;
    assign weights1[20][173] = 16'b1111111110110101;
    assign weights1[20][174] = 16'b1111111110101001;
    assign weights1[20][175] = 16'b1111111110011101;
    assign weights1[20][176] = 16'b1111111110100110;
    assign weights1[20][177] = 16'b1111111110010100;
    assign weights1[20][178] = 16'b1111111110011000;
    assign weights1[20][179] = 16'b1111111110100000;
    assign weights1[20][180] = 16'b1111111110101011;
    assign weights1[20][181] = 16'b1111111110011101;
    assign weights1[20][182] = 16'b1111111110101010;
    assign weights1[20][183] = 16'b1111111110011011;
    assign weights1[20][184] = 16'b1111111110111000;
    assign weights1[20][185] = 16'b1111111110110001;
    assign weights1[20][186] = 16'b1111111110101110;
    assign weights1[20][187] = 16'b1111111110111010;
    assign weights1[20][188] = 16'b1111111110111011;
    assign weights1[20][189] = 16'b1111111110111111;
    assign weights1[20][190] = 16'b1111111111001101;
    assign weights1[20][191] = 16'b1111111111011011;
    assign weights1[20][192] = 16'b1111111111011110;
    assign weights1[20][193] = 16'b1111111111011110;
    assign weights1[20][194] = 16'b1111111111100110;
    assign weights1[20][195] = 16'b1111111111110000;
    assign weights1[20][196] = 16'b1111111111111101;
    assign weights1[20][197] = 16'b1111111111110100;
    assign weights1[20][198] = 16'b1111111111100110;
    assign weights1[20][199] = 16'b1111111111000111;
    assign weights1[20][200] = 16'b1111111110110011;
    assign weights1[20][201] = 16'b1111111110011111;
    assign weights1[20][202] = 16'b1111111110000000;
    assign weights1[20][203] = 16'b1111111110000111;
    assign weights1[20][204] = 16'b1111111110100110;
    assign weights1[20][205] = 16'b1111111110010000;
    assign weights1[20][206] = 16'b1111111110001010;
    assign weights1[20][207] = 16'b1111111110010000;
    assign weights1[20][208] = 16'b1111111110010111;
    assign weights1[20][209] = 16'b1111111110010011;
    assign weights1[20][210] = 16'b1111111110011111;
    assign weights1[20][211] = 16'b1111111110100101;
    assign weights1[20][212] = 16'b1111111110111011;
    assign weights1[20][213] = 16'b1111111110010111;
    assign weights1[20][214] = 16'b1111111110010101;
    assign weights1[20][215] = 16'b1111111110100101;
    assign weights1[20][216] = 16'b1111111110010101;
    assign weights1[20][217] = 16'b1111111110101100;
    assign weights1[20][218] = 16'b1111111110111100;
    assign weights1[20][219] = 16'b1111111111001011;
    assign weights1[20][220] = 16'b1111111111001101;
    assign weights1[20][221] = 16'b1111111111011101;
    assign weights1[20][222] = 16'b1111111111011101;
    assign weights1[20][223] = 16'b1111111111101101;
    assign weights1[20][224] = 16'b1111111111111100;
    assign weights1[20][225] = 16'b1111111111110101;
    assign weights1[20][226] = 16'b1111111111100100;
    assign weights1[20][227] = 16'b1111111111001101;
    assign weights1[20][228] = 16'b1111111110111100;
    assign weights1[20][229] = 16'b1111111110101010;
    assign weights1[20][230] = 16'b1111111110111010;
    assign weights1[20][231] = 16'b1111111111001101;
    assign weights1[20][232] = 16'b1111111110110000;
    assign weights1[20][233] = 16'b1111111110101110;
    assign weights1[20][234] = 16'b1111111110111010;
    assign weights1[20][235] = 16'b1111111111000100;
    assign weights1[20][236] = 16'b1111111111001000;
    assign weights1[20][237] = 16'b1111111111011010;
    assign weights1[20][238] = 16'b1111111111001010;
    assign weights1[20][239] = 16'b1111111111010110;
    assign weights1[20][240] = 16'b1111111110111110;
    assign weights1[20][241] = 16'b1111111110111111;
    assign weights1[20][242] = 16'b1111111111000110;
    assign weights1[20][243] = 16'b1111111111010011;
    assign weights1[20][244] = 16'b1111111111001111;
    assign weights1[20][245] = 16'b1111111111100010;
    assign weights1[20][246] = 16'b1111111110111111;
    assign weights1[20][247] = 16'b1111111110111101;
    assign weights1[20][248] = 16'b1111111111000110;
    assign weights1[20][249] = 16'b1111111111100001;
    assign weights1[20][250] = 16'b1111111111110000;
    assign weights1[20][251] = 16'b1111111111111000;
    assign weights1[20][252] = 16'b0000000000000111;
    assign weights1[20][253] = 16'b1111111111111100;
    assign weights1[20][254] = 16'b1111111111101010;
    assign weights1[20][255] = 16'b1111111111101000;
    assign weights1[20][256] = 16'b1111111111101100;
    assign weights1[20][257] = 16'b1111111111101101;
    assign weights1[20][258] = 16'b1111111111110001;
    assign weights1[20][259] = 16'b1111111111110011;
    assign weights1[20][260] = 16'b1111111111111011;
    assign weights1[20][261] = 16'b1111111111011100;
    assign weights1[20][262] = 16'b1111111111001111;
    assign weights1[20][263] = 16'b1111111111011001;
    assign weights1[20][264] = 16'b1111111111011100;
    assign weights1[20][265] = 16'b1111111111011111;
    assign weights1[20][266] = 16'b1111111111001100;
    assign weights1[20][267] = 16'b1111111111100000;
    assign weights1[20][268] = 16'b1111111111010111;
    assign weights1[20][269] = 16'b1111111111101010;
    assign weights1[20][270] = 16'b1111111111010011;
    assign weights1[20][271] = 16'b1111111111011100;
    assign weights1[20][272] = 16'b1111111111100010;
    assign weights1[20][273] = 16'b1111111111110111;
    assign weights1[20][274] = 16'b1111111111010110;
    assign weights1[20][275] = 16'b1111111111101110;
    assign weights1[20][276] = 16'b1111111111101111;
    assign weights1[20][277] = 16'b1111111111111000;
    assign weights1[20][278] = 16'b1111111111111000;
    assign weights1[20][279] = 16'b0000000000001110;
    assign weights1[20][280] = 16'b0000000000001010;
    assign weights1[20][281] = 16'b0000000000000110;
    assign weights1[20][282] = 16'b1111111111110010;
    assign weights1[20][283] = 16'b1111111111111011;
    assign weights1[20][284] = 16'b1111111111111101;
    assign weights1[20][285] = 16'b0000000000000000;
    assign weights1[20][286] = 16'b0000000000000011;
    assign weights1[20][287] = 16'b0000000000100100;
    assign weights1[20][288] = 16'b0000000000000100;
    assign weights1[20][289] = 16'b0000000000100000;
    assign weights1[20][290] = 16'b0000000000000000;
    assign weights1[20][291] = 16'b1111111111110100;
    assign weights1[20][292] = 16'b1111111111010111;
    assign weights1[20][293] = 16'b1111111111010101;
    assign weights1[20][294] = 16'b1111111111011010;
    assign weights1[20][295] = 16'b1111111111100011;
    assign weights1[20][296] = 16'b1111111111100101;
    assign weights1[20][297] = 16'b1111111111111101;
    assign weights1[20][298] = 16'b1111111111101000;
    assign weights1[20][299] = 16'b1111111111100101;
    assign weights1[20][300] = 16'b0000000000000000;
    assign weights1[20][301] = 16'b1111111111110000;
    assign weights1[20][302] = 16'b0000000000011001;
    assign weights1[20][303] = 16'b1111111111110010;
    assign weights1[20][304] = 16'b1111111111110000;
    assign weights1[20][305] = 16'b0000000000010001;
    assign weights1[20][306] = 16'b1111111111111101;
    assign weights1[20][307] = 16'b1111111111111100;
    assign weights1[20][308] = 16'b0000000000000101;
    assign weights1[20][309] = 16'b0000000000000010;
    assign weights1[20][310] = 16'b0000000000001001;
    assign weights1[20][311] = 16'b0000000000001000;
    assign weights1[20][312] = 16'b0000000000100001;
    assign weights1[20][313] = 16'b0000000000010100;
    assign weights1[20][314] = 16'b0000000000011011;
    assign weights1[20][315] = 16'b0000000000011101;
    assign weights1[20][316] = 16'b0000000000100001;
    assign weights1[20][317] = 16'b0000000000001100;
    assign weights1[20][318] = 16'b0000000000001001;
    assign weights1[20][319] = 16'b0000000000010101;
    assign weights1[20][320] = 16'b0000000000100001;
    assign weights1[20][321] = 16'b0000000000010011;
    assign weights1[20][322] = 16'b1111111111111110;
    assign weights1[20][323] = 16'b1111111111111110;
    assign weights1[20][324] = 16'b1111111111111011;
    assign weights1[20][325] = 16'b1111111111110001;
    assign weights1[20][326] = 16'b0000000000000011;
    assign weights1[20][327] = 16'b1111111111111111;
    assign weights1[20][328] = 16'b0000000000000010;
    assign weights1[20][329] = 16'b0000000000000001;
    assign weights1[20][330] = 16'b0000000000000010;
    assign weights1[20][331] = 16'b1111111111100110;
    assign weights1[20][332] = 16'b1111111111111011;
    assign weights1[20][333] = 16'b0000000000000001;
    assign weights1[20][334] = 16'b1111111111111010;
    assign weights1[20][335] = 16'b1111111111111110;
    assign weights1[20][336] = 16'b0000000000001011;
    assign weights1[20][337] = 16'b0000000000001000;
    assign weights1[20][338] = 16'b0000000000000000;
    assign weights1[20][339] = 16'b0000000000010011;
    assign weights1[20][340] = 16'b0000000000000011;
    assign weights1[20][341] = 16'b0000000000001101;
    assign weights1[20][342] = 16'b1111111111110110;
    assign weights1[20][343] = 16'b0000000000011100;
    assign weights1[20][344] = 16'b0000000000101111;
    assign weights1[20][345] = 16'b0000000000011110;
    assign weights1[20][346] = 16'b0000000000101000;
    assign weights1[20][347] = 16'b0000000000100011;
    assign weights1[20][348] = 16'b0000000000100101;
    assign weights1[20][349] = 16'b0000000000101010;
    assign weights1[20][350] = 16'b0000000000010111;
    assign weights1[20][351] = 16'b0000000000011001;
    assign weights1[20][352] = 16'b0000000000001010;
    assign weights1[20][353] = 16'b0000000000011110;
    assign weights1[20][354] = 16'b0000000000001001;
    assign weights1[20][355] = 16'b0000000000001110;
    assign weights1[20][356] = 16'b1111111111111111;
    assign weights1[20][357] = 16'b1111111111111111;
    assign weights1[20][358] = 16'b1111111111111101;
    assign weights1[20][359] = 16'b0000000000001010;
    assign weights1[20][360] = 16'b1111111111111101;
    assign weights1[20][361] = 16'b0000000000000001;
    assign weights1[20][362] = 16'b0000000000000100;
    assign weights1[20][363] = 16'b0000000000000110;
    assign weights1[20][364] = 16'b0000000000010001;
    assign weights1[20][365] = 16'b0000000000010110;
    assign weights1[20][366] = 16'b0000000000011010;
    assign weights1[20][367] = 16'b0000000000011011;
    assign weights1[20][368] = 16'b0000000000010101;
    assign weights1[20][369] = 16'b0000000000010011;
    assign weights1[20][370] = 16'b0000000000000011;
    assign weights1[20][371] = 16'b0000000000011010;
    assign weights1[20][372] = 16'b0000000000011000;
    assign weights1[20][373] = 16'b0000000000100001;
    assign weights1[20][374] = 16'b0000000000100101;
    assign weights1[20][375] = 16'b0000000000110000;
    assign weights1[20][376] = 16'b0000000000101110;
    assign weights1[20][377] = 16'b0000000000011011;
    assign weights1[20][378] = 16'b0000000000100010;
    assign weights1[20][379] = 16'b0000000000011000;
    assign weights1[20][380] = 16'b0000000000011000;
    assign weights1[20][381] = 16'b0000000000010110;
    assign weights1[20][382] = 16'b0000000000010110;
    assign weights1[20][383] = 16'b0000000000001010;
    assign weights1[20][384] = 16'b0000000000010111;
    assign weights1[20][385] = 16'b0000000000010001;
    assign weights1[20][386] = 16'b0000000000011101;
    assign weights1[20][387] = 16'b1111111111111010;
    assign weights1[20][388] = 16'b0000000000001101;
    assign weights1[20][389] = 16'b0000000000010110;
    assign weights1[20][390] = 16'b0000000000010011;
    assign weights1[20][391] = 16'b0000000000010111;
    assign weights1[20][392] = 16'b0000000000011100;
    assign weights1[20][393] = 16'b0000000000101100;
    assign weights1[20][394] = 16'b0000000000010001;
    assign weights1[20][395] = 16'b0000000000010111;
    assign weights1[20][396] = 16'b0000000000000011;
    assign weights1[20][397] = 16'b0000000000001010;
    assign weights1[20][398] = 16'b0000000000010110;
    assign weights1[20][399] = 16'b0000000000000111;
    assign weights1[20][400] = 16'b0000000000011011;
    assign weights1[20][401] = 16'b0000000000001100;
    assign weights1[20][402] = 16'b0000000000001110;
    assign weights1[20][403] = 16'b0000000000100000;
    assign weights1[20][404] = 16'b0000000000001000;
    assign weights1[20][405] = 16'b0000000000101001;
    assign weights1[20][406] = 16'b0000000000011011;
    assign weights1[20][407] = 16'b0000000000011100;
    assign weights1[20][408] = 16'b0000000000010110;
    assign weights1[20][409] = 16'b0000000000000100;
    assign weights1[20][410] = 16'b0000000000011010;
    assign weights1[20][411] = 16'b0000000000000110;
    assign weights1[20][412] = 16'b0000000000000000;
    assign weights1[20][413] = 16'b0000000000001011;
    assign weights1[20][414] = 16'b0000000000000110;
    assign weights1[20][415] = 16'b0000000000010111;
    assign weights1[20][416] = 16'b0000000000000111;
    assign weights1[20][417] = 16'b1111111111111100;
    assign weights1[20][418] = 16'b0000000000001110;
    assign weights1[20][419] = 16'b0000000000011000;
    assign weights1[20][420] = 16'b0000000000011100;
    assign weights1[20][421] = 16'b0000000000011110;
    assign weights1[20][422] = 16'b0000000000000111;
    assign weights1[20][423] = 16'b0000000000001110;
    assign weights1[20][424] = 16'b0000000000001000;
    assign weights1[20][425] = 16'b0000000000001001;
    assign weights1[20][426] = 16'b0000000000010110;
    assign weights1[20][427] = 16'b1111111111111100;
    assign weights1[20][428] = 16'b0000000000010001;
    assign weights1[20][429] = 16'b0000000000000011;
    assign weights1[20][430] = 16'b0000000000000100;
    assign weights1[20][431] = 16'b0000000000001001;
    assign weights1[20][432] = 16'b0000000000001011;
    assign weights1[20][433] = 16'b0000000000000100;
    assign weights1[20][434] = 16'b0000000000001100;
    assign weights1[20][435] = 16'b0000000000010010;
    assign weights1[20][436] = 16'b0000000000001000;
    assign weights1[20][437] = 16'b0000000000000100;
    assign weights1[20][438] = 16'b0000000000010001;
    assign weights1[20][439] = 16'b0000000000001001;
    assign weights1[20][440] = 16'b0000000000010100;
    assign weights1[20][441] = 16'b0000000000000010;
    assign weights1[20][442] = 16'b0000000000001111;
    assign weights1[20][443] = 16'b0000000000000011;
    assign weights1[20][444] = 16'b0000000000001011;
    assign weights1[20][445] = 16'b1111111111111111;
    assign weights1[20][446] = 16'b0000000000001110;
    assign weights1[20][447] = 16'b0000000000001110;
    assign weights1[20][448] = 16'b0000000000100000;
    assign weights1[20][449] = 16'b0000000000100100;
    assign weights1[20][450] = 16'b0000000000001000;
    assign weights1[20][451] = 16'b0000000000001011;
    assign weights1[20][452] = 16'b0000000000000111;
    assign weights1[20][453] = 16'b1111111111110101;
    assign weights1[20][454] = 16'b0000000000010000;
    assign weights1[20][455] = 16'b0000000000010011;
    assign weights1[20][456] = 16'b1111111111110110;
    assign weights1[20][457] = 16'b0000000000000101;
    assign weights1[20][458] = 16'b1111111111101001;
    assign weights1[20][459] = 16'b1111111111110110;
    assign weights1[20][460] = 16'b1111111111111001;
    assign weights1[20][461] = 16'b1111111111111101;
    assign weights1[20][462] = 16'b0000000000000000;
    assign weights1[20][463] = 16'b0000000000001011;
    assign weights1[20][464] = 16'b1111111111110000;
    assign weights1[20][465] = 16'b1111111111111111;
    assign weights1[20][466] = 16'b1111111111111111;
    assign weights1[20][467] = 16'b1111111111110001;
    assign weights1[20][468] = 16'b1111111111111111;
    assign weights1[20][469] = 16'b0000000000000101;
    assign weights1[20][470] = 16'b1111111111111100;
    assign weights1[20][471] = 16'b0000000000010000;
    assign weights1[20][472] = 16'b0000000000010111;
    assign weights1[20][473] = 16'b0000000000011000;
    assign weights1[20][474] = 16'b0000000000011110;
    assign weights1[20][475] = 16'b0000000000001100;
    assign weights1[20][476] = 16'b0000000000000111;
    assign weights1[20][477] = 16'b0000000000011000;
    assign weights1[20][478] = 16'b0000000000001001;
    assign weights1[20][479] = 16'b0000000000001010;
    assign weights1[20][480] = 16'b0000000000000101;
    assign weights1[20][481] = 16'b0000000000011011;
    assign weights1[20][482] = 16'b0000000000001111;
    assign weights1[20][483] = 16'b0000000000000001;
    assign weights1[20][484] = 16'b0000000000000001;
    assign weights1[20][485] = 16'b1111111111111010;
    assign weights1[20][486] = 16'b1111111111111101;
    assign weights1[20][487] = 16'b1111111111100101;
    assign weights1[20][488] = 16'b0000000000000010;
    assign weights1[20][489] = 16'b1111111111110111;
    assign weights1[20][490] = 16'b1111111111101010;
    assign weights1[20][491] = 16'b1111111111100101;
    assign weights1[20][492] = 16'b1111111111101010;
    assign weights1[20][493] = 16'b1111111111101110;
    assign weights1[20][494] = 16'b0000000000000100;
    assign weights1[20][495] = 16'b1111111111110010;
    assign weights1[20][496] = 16'b0000000000001001;
    assign weights1[20][497] = 16'b0000000000011001;
    assign weights1[20][498] = 16'b0000000000010111;
    assign weights1[20][499] = 16'b0000000000000011;
    assign weights1[20][500] = 16'b0000000000011011;
    assign weights1[20][501] = 16'b0000000000010000;
    assign weights1[20][502] = 16'b0000000000100010;
    assign weights1[20][503] = 16'b0000000000000010;
    assign weights1[20][504] = 16'b1111111111110101;
    assign weights1[20][505] = 16'b0000000000001110;
    assign weights1[20][506] = 16'b0000000000011001;
    assign weights1[20][507] = 16'b0000000000001000;
    assign weights1[20][508] = 16'b0000000000011001;
    assign weights1[20][509] = 16'b0000000000000110;
    assign weights1[20][510] = 16'b1111111111110101;
    assign weights1[20][511] = 16'b0000000000001100;
    assign weights1[20][512] = 16'b0000000000000001;
    assign weights1[20][513] = 16'b1111111111111111;
    assign weights1[20][514] = 16'b1111111111110100;
    assign weights1[20][515] = 16'b1111111111100100;
    assign weights1[20][516] = 16'b0000000000001001;
    assign weights1[20][517] = 16'b1111111111110001;
    assign weights1[20][518] = 16'b1111111111100100;
    assign weights1[20][519] = 16'b1111111111111110;
    assign weights1[20][520] = 16'b1111111111110111;
    assign weights1[20][521] = 16'b1111111111111001;
    assign weights1[20][522] = 16'b0000000000000101;
    assign weights1[20][523] = 16'b0000000000000111;
    assign weights1[20][524] = 16'b0000000000000101;
    assign weights1[20][525] = 16'b0000000000001100;
    assign weights1[20][526] = 16'b0000000000010100;
    assign weights1[20][527] = 16'b0000000000010011;
    assign weights1[20][528] = 16'b0000000000001010;
    assign weights1[20][529] = 16'b0000000000010111;
    assign weights1[20][530] = 16'b0000000000010101;
    assign weights1[20][531] = 16'b0000000000000000;
    assign weights1[20][532] = 16'b1111111111110010;
    assign weights1[20][533] = 16'b0000000000000111;
    assign weights1[20][534] = 16'b0000000000001110;
    assign weights1[20][535] = 16'b0000000000001010;
    assign weights1[20][536] = 16'b0000000000001100;
    assign weights1[20][537] = 16'b0000000000000100;
    assign weights1[20][538] = 16'b0000000000000011;
    assign weights1[20][539] = 16'b1111111111111111;
    assign weights1[20][540] = 16'b1111111111110111;
    assign weights1[20][541] = 16'b1111111111111111;
    assign weights1[20][542] = 16'b0000000000000111;
    assign weights1[20][543] = 16'b0000000000010001;
    assign weights1[20][544] = 16'b0000000000001001;
    assign weights1[20][545] = 16'b0000000000001100;
    assign weights1[20][546] = 16'b1111111111111111;
    assign weights1[20][547] = 16'b0000000000000110;
    assign weights1[20][548] = 16'b1111111111111111;
    assign weights1[20][549] = 16'b0000000000000000;
    assign weights1[20][550] = 16'b0000000000010001;
    assign weights1[20][551] = 16'b0000000000000111;
    assign weights1[20][552] = 16'b0000000000000111;
    assign weights1[20][553] = 16'b0000000000000011;
    assign weights1[20][554] = 16'b0000000000001001;
    assign weights1[20][555] = 16'b1111111111111000;
    assign weights1[20][556] = 16'b0000000000000110;
    assign weights1[20][557] = 16'b0000000000000001;
    assign weights1[20][558] = 16'b0000000000000111;
    assign weights1[20][559] = 16'b0000000000000101;
    assign weights1[20][560] = 16'b1111111111101111;
    assign weights1[20][561] = 16'b0000000000000000;
    assign weights1[20][562] = 16'b0000000000000110;
    assign weights1[20][563] = 16'b1111111111111010;
    assign weights1[20][564] = 16'b1111111111111100;
    assign weights1[20][565] = 16'b0000000000001010;
    assign weights1[20][566] = 16'b1111111111111011;
    assign weights1[20][567] = 16'b0000000000000100;
    assign weights1[20][568] = 16'b0000000000001111;
    assign weights1[20][569] = 16'b0000000000000110;
    assign weights1[20][570] = 16'b0000000000000011;
    assign weights1[20][571] = 16'b0000000000000110;
    assign weights1[20][572] = 16'b0000000000010101;
    assign weights1[20][573] = 16'b0000000000010001;
    assign weights1[20][574] = 16'b0000000000000101;
    assign weights1[20][575] = 16'b0000000000001000;
    assign weights1[20][576] = 16'b0000000000010001;
    assign weights1[20][577] = 16'b0000000000000011;
    assign weights1[20][578] = 16'b0000000000010001;
    assign weights1[20][579] = 16'b1111111111111011;
    assign weights1[20][580] = 16'b0000000000010010;
    assign weights1[20][581] = 16'b0000000000011000;
    assign weights1[20][582] = 16'b0000000000001000;
    assign weights1[20][583] = 16'b0000000000001010;
    assign weights1[20][584] = 16'b1111111111110111;
    assign weights1[20][585] = 16'b1111111111110101;
    assign weights1[20][586] = 16'b1111111111111100;
    assign weights1[20][587] = 16'b0000000000000101;
    assign weights1[20][588] = 16'b1111111111110001;
    assign weights1[20][589] = 16'b1111111111101111;
    assign weights1[20][590] = 16'b1111111111101100;
    assign weights1[20][591] = 16'b1111111111111001;
    assign weights1[20][592] = 16'b1111111111101011;
    assign weights1[20][593] = 16'b0000000000001111;
    assign weights1[20][594] = 16'b0000000000000011;
    assign weights1[20][595] = 16'b0000000000000011;
    assign weights1[20][596] = 16'b0000000000000110;
    assign weights1[20][597] = 16'b0000000000000101;
    assign weights1[20][598] = 16'b0000000000010110;
    assign weights1[20][599] = 16'b0000000000000010;
    assign weights1[20][600] = 16'b1111111111111101;
    assign weights1[20][601] = 16'b0000000000001010;
    assign weights1[20][602] = 16'b0000000000001100;
    assign weights1[20][603] = 16'b0000000000010110;
    assign weights1[20][604] = 16'b0000000000001000;
    assign weights1[20][605] = 16'b0000000000000011;
    assign weights1[20][606] = 16'b0000000000010110;
    assign weights1[20][607] = 16'b1111111111111000;
    assign weights1[20][608] = 16'b0000000000000001;
    assign weights1[20][609] = 16'b0000000000000000;
    assign weights1[20][610] = 16'b1111111111110111;
    assign weights1[20][611] = 16'b0000000000000001;
    assign weights1[20][612] = 16'b1111111111111110;
    assign weights1[20][613] = 16'b1111111111111010;
    assign weights1[20][614] = 16'b1111111111110111;
    assign weights1[20][615] = 16'b0000000000000001;
    assign weights1[20][616] = 16'b1111111111111000;
    assign weights1[20][617] = 16'b1111111111110000;
    assign weights1[20][618] = 16'b1111111111101001;
    assign weights1[20][619] = 16'b1111111111110110;
    assign weights1[20][620] = 16'b1111111111110001;
    assign weights1[20][621] = 16'b1111111111101111;
    assign weights1[20][622] = 16'b1111111111110101;
    assign weights1[20][623] = 16'b1111111111110101;
    assign weights1[20][624] = 16'b1111111111111001;
    assign weights1[20][625] = 16'b1111111111110110;
    assign weights1[20][626] = 16'b1111111111101111;
    assign weights1[20][627] = 16'b1111111111101001;
    assign weights1[20][628] = 16'b0000000000000110;
    assign weights1[20][629] = 16'b0000000000001100;
    assign weights1[20][630] = 16'b1111111111110111;
    assign weights1[20][631] = 16'b1111111111111101;
    assign weights1[20][632] = 16'b1111111111111000;
    assign weights1[20][633] = 16'b0000000000000111;
    assign weights1[20][634] = 16'b0000000000001001;
    assign weights1[20][635] = 16'b1111111111111111;
    assign weights1[20][636] = 16'b0000000000000001;
    assign weights1[20][637] = 16'b0000000000001001;
    assign weights1[20][638] = 16'b0000000000000100;
    assign weights1[20][639] = 16'b1111111111110000;
    assign weights1[20][640] = 16'b1111111111111000;
    assign weights1[20][641] = 16'b1111111111110111;
    assign weights1[20][642] = 16'b1111111111110011;
    assign weights1[20][643] = 16'b1111111111111000;
    assign weights1[20][644] = 16'b1111111111110101;
    assign weights1[20][645] = 16'b1111111111100111;
    assign weights1[20][646] = 16'b1111111111100100;
    assign weights1[20][647] = 16'b1111111111100111;
    assign weights1[20][648] = 16'b1111111111110001;
    assign weights1[20][649] = 16'b1111111111110010;
    assign weights1[20][650] = 16'b1111111111100000;
    assign weights1[20][651] = 16'b1111111111101010;
    assign weights1[20][652] = 16'b1111111111110101;
    assign weights1[20][653] = 16'b1111111111110100;
    assign weights1[20][654] = 16'b1111111111111011;
    assign weights1[20][655] = 16'b1111111111110000;
    assign weights1[20][656] = 16'b1111111111101111;
    assign weights1[20][657] = 16'b1111111111111100;
    assign weights1[20][658] = 16'b1111111111111101;
    assign weights1[20][659] = 16'b1111111111111001;
    assign weights1[20][660] = 16'b0000000000000001;
    assign weights1[20][661] = 16'b1111111111111010;
    assign weights1[20][662] = 16'b0000000000000000;
    assign weights1[20][663] = 16'b1111111111101111;
    assign weights1[20][664] = 16'b1111111111111001;
    assign weights1[20][665] = 16'b1111111111101101;
    assign weights1[20][666] = 16'b1111111111101010;
    assign weights1[20][667] = 16'b1111111111101011;
    assign weights1[20][668] = 16'b1111111111111110;
    assign weights1[20][669] = 16'b0000000000000001;
    assign weights1[20][670] = 16'b1111111111110111;
    assign weights1[20][671] = 16'b0000000000000011;
    assign weights1[20][672] = 16'b1111111111110110;
    assign weights1[20][673] = 16'b1111111111100111;
    assign weights1[20][674] = 16'b1111111111110001;
    assign weights1[20][675] = 16'b1111111111111000;
    assign weights1[20][676] = 16'b1111111111011110;
    assign weights1[20][677] = 16'b1111111111100001;
    assign weights1[20][678] = 16'b1111111111101101;
    assign weights1[20][679] = 16'b1111111111100101;
    assign weights1[20][680] = 16'b1111111111110001;
    assign weights1[20][681] = 16'b0000000000001010;
    assign weights1[20][682] = 16'b1111111111110110;
    assign weights1[20][683] = 16'b1111111111111001;
    assign weights1[20][684] = 16'b0000000000000001;
    assign weights1[20][685] = 16'b1111111111111110;
    assign weights1[20][686] = 16'b1111111111110101;
    assign weights1[20][687] = 16'b1111111111101011;
    assign weights1[20][688] = 16'b1111111111111100;
    assign weights1[20][689] = 16'b1111111111111111;
    assign weights1[20][690] = 16'b1111111111111000;
    assign weights1[20][691] = 16'b1111111111111001;
    assign weights1[20][692] = 16'b1111111111110010;
    assign weights1[20][693] = 16'b1111111111110010;
    assign weights1[20][694] = 16'b1111111111111000;
    assign weights1[20][695] = 16'b1111111111101110;
    assign weights1[20][696] = 16'b0000000000001001;
    assign weights1[20][697] = 16'b0000000000001010;
    assign weights1[20][698] = 16'b1111111111111111;
    assign weights1[20][699] = 16'b0000000000000110;
    assign weights1[20][700] = 16'b0000000000000011;
    assign weights1[20][701] = 16'b1111111111110011;
    assign weights1[20][702] = 16'b1111111111110110;
    assign weights1[20][703] = 16'b1111111111111001;
    assign weights1[20][704] = 16'b1111111111110111;
    assign weights1[20][705] = 16'b1111111111100010;
    assign weights1[20][706] = 16'b1111111111100111;
    assign weights1[20][707] = 16'b1111111111101001;
    assign weights1[20][708] = 16'b1111111111011011;
    assign weights1[20][709] = 16'b1111111111100000;
    assign weights1[20][710] = 16'b1111111111101101;
    assign weights1[20][711] = 16'b1111111111101000;
    assign weights1[20][712] = 16'b1111111111100001;
    assign weights1[20][713] = 16'b1111111111101100;
    assign weights1[20][714] = 16'b1111111111110101;
    assign weights1[20][715] = 16'b1111111111101011;
    assign weights1[20][716] = 16'b1111111111101010;
    assign weights1[20][717] = 16'b1111111111111000;
    assign weights1[20][718] = 16'b1111111111011101;
    assign weights1[20][719] = 16'b1111111111011011;
    assign weights1[20][720] = 16'b1111111111110010;
    assign weights1[20][721] = 16'b1111111111111000;
    assign weights1[20][722] = 16'b1111111111111001;
    assign weights1[20][723] = 16'b1111111111110000;
    assign weights1[20][724] = 16'b0000000000010010;
    assign weights1[20][725] = 16'b0000000000010000;
    assign weights1[20][726] = 16'b0000000000000000;
    assign weights1[20][727] = 16'b0000000000001010;
    assign weights1[20][728] = 16'b0000000000000100;
    assign weights1[20][729] = 16'b0000000000000001;
    assign weights1[20][730] = 16'b0000000000000111;
    assign weights1[20][731] = 16'b0000000000001011;
    assign weights1[20][732] = 16'b1111111111111110;
    assign weights1[20][733] = 16'b1111111111111110;
    assign weights1[20][734] = 16'b1111111111111011;
    assign weights1[20][735] = 16'b1111111111111111;
    assign weights1[20][736] = 16'b1111111111110011;
    assign weights1[20][737] = 16'b1111111111110100;
    assign weights1[20][738] = 16'b1111111111101100;
    assign weights1[20][739] = 16'b1111111111101100;
    assign weights1[20][740] = 16'b1111111111101100;
    assign weights1[20][741] = 16'b1111111111010101;
    assign weights1[20][742] = 16'b1111111111100111;
    assign weights1[20][743] = 16'b1111111111101010;
    assign weights1[20][744] = 16'b1111111111010110;
    assign weights1[20][745] = 16'b1111111111101110;
    assign weights1[20][746] = 16'b1111111111110110;
    assign weights1[20][747] = 16'b1111111111100110;
    assign weights1[20][748] = 16'b1111111111101101;
    assign weights1[20][749] = 16'b0000000000000100;
    assign weights1[20][750] = 16'b0000000000001001;
    assign weights1[20][751] = 16'b0000000000010011;
    assign weights1[20][752] = 16'b0000000000010110;
    assign weights1[20][753] = 16'b0000000000011000;
    assign weights1[20][754] = 16'b0000000000001110;
    assign weights1[20][755] = 16'b0000000000001010;
    assign weights1[20][756] = 16'b0000000000000100;
    assign weights1[20][757] = 16'b0000000000000100;
    assign weights1[20][758] = 16'b0000000000000110;
    assign weights1[20][759] = 16'b0000000000000100;
    assign weights1[20][760] = 16'b0000000000001000;
    assign weights1[20][761] = 16'b0000000000010010;
    assign weights1[20][762] = 16'b0000000000011100;
    assign weights1[20][763] = 16'b0000000000010010;
    assign weights1[20][764] = 16'b0000000000010101;
    assign weights1[20][765] = 16'b0000000000001110;
    assign weights1[20][766] = 16'b0000000000001100;
    assign weights1[20][767] = 16'b0000000000001111;
    assign weights1[20][768] = 16'b0000000000010010;
    assign weights1[20][769] = 16'b0000000000011011;
    assign weights1[20][770] = 16'b0000000000010001;
    assign weights1[20][771] = 16'b0000000000001101;
    assign weights1[20][772] = 16'b0000000000011101;
    assign weights1[20][773] = 16'b0000000000011001;
    assign weights1[20][774] = 16'b0000000000011011;
    assign weights1[20][775] = 16'b0000000000010101;
    assign weights1[20][776] = 16'b0000000000100010;
    assign weights1[20][777] = 16'b0000000000100001;
    assign weights1[20][778] = 16'b0000000000010101;
    assign weights1[20][779] = 16'b0000000000011000;
    assign weights1[20][780] = 16'b0000000000011110;
    assign weights1[20][781] = 16'b0000000000011011;
    assign weights1[20][782] = 16'b0000000000010111;
    assign weights1[20][783] = 16'b0000000000000110;
    assign weights1[21][0] = 16'b0000000000000000;
    assign weights1[21][1] = 16'b1111111111111111;
    assign weights1[21][2] = 16'b1111111111111111;
    assign weights1[21][3] = 16'b1111111111111111;
    assign weights1[21][4] = 16'b1111111111111111;
    assign weights1[21][5] = 16'b1111111111111111;
    assign weights1[21][6] = 16'b1111111111110111;
    assign weights1[21][7] = 16'b1111111111111000;
    assign weights1[21][8] = 16'b1111111111101100;
    assign weights1[21][9] = 16'b1111111111101010;
    assign weights1[21][10] = 16'b1111111111100101;
    assign weights1[21][11] = 16'b1111111111100000;
    assign weights1[21][12] = 16'b1111111111100011;
    assign weights1[21][13] = 16'b1111111111101100;
    assign weights1[21][14] = 16'b1111111111111010;
    assign weights1[21][15] = 16'b1111111111111110;
    assign weights1[21][16] = 16'b0000000000001001;
    assign weights1[21][17] = 16'b0000000000001010;
    assign weights1[21][18] = 16'b0000000000000100;
    assign weights1[21][19] = 16'b1111111111111110;
    assign weights1[21][20] = 16'b0000000000000110;
    assign weights1[21][21] = 16'b0000000000000100;
    assign weights1[21][22] = 16'b0000000000001100;
    assign weights1[21][23] = 16'b0000000000001010;
    assign weights1[21][24] = 16'b0000000000000100;
    assign weights1[21][25] = 16'b0000000000000010;
    assign weights1[21][26] = 16'b1111111111111110;
    assign weights1[21][27] = 16'b0000000000000011;
    assign weights1[21][28] = 16'b0000000000000000;
    assign weights1[21][29] = 16'b1111111111111111;
    assign weights1[21][30] = 16'b0000000000000000;
    assign weights1[21][31] = 16'b0000000000000000;
    assign weights1[21][32] = 16'b1111111111111110;
    assign weights1[21][33] = 16'b1111111111111010;
    assign weights1[21][34] = 16'b1111111111110000;
    assign weights1[21][35] = 16'b1111111111110011;
    assign weights1[21][36] = 16'b1111111111110000;
    assign weights1[21][37] = 16'b1111111111101001;
    assign weights1[21][38] = 16'b1111111111100010;
    assign weights1[21][39] = 16'b1111111111011011;
    assign weights1[21][40] = 16'b1111111111010100;
    assign weights1[21][41] = 16'b1111111111010101;
    assign weights1[21][42] = 16'b1111111111111001;
    assign weights1[21][43] = 16'b0000000000001011;
    assign weights1[21][44] = 16'b0000000000000011;
    assign weights1[21][45] = 16'b0000000000000011;
    assign weights1[21][46] = 16'b1111111111111001;
    assign weights1[21][47] = 16'b1111111111111101;
    assign weights1[21][48] = 16'b0000000000000111;
    assign weights1[21][49] = 16'b0000000000001100;
    assign weights1[21][50] = 16'b0000000000010011;
    assign weights1[21][51] = 16'b1111111111111111;
    assign weights1[21][52] = 16'b0000000000000010;
    assign weights1[21][53] = 16'b1111111111111101;
    assign weights1[21][54] = 16'b1111111111111111;
    assign weights1[21][55] = 16'b1111111111111110;
    assign weights1[21][56] = 16'b1111111111111111;
    assign weights1[21][57] = 16'b0000000000000001;
    assign weights1[21][58] = 16'b1111111111111111;
    assign weights1[21][59] = 16'b1111111111111101;
    assign weights1[21][60] = 16'b1111111111110011;
    assign weights1[21][61] = 16'b1111111111110010;
    assign weights1[21][62] = 16'b1111111111101101;
    assign weights1[21][63] = 16'b1111111111111000;
    assign weights1[21][64] = 16'b1111111111110001;
    assign weights1[21][65] = 16'b1111111111101010;
    assign weights1[21][66] = 16'b1111111111010101;
    assign weights1[21][67] = 16'b1111111111001110;
    assign weights1[21][68] = 16'b1111111111011011;
    assign weights1[21][69] = 16'b1111111111101101;
    assign weights1[21][70] = 16'b1111111111111010;
    assign weights1[21][71] = 16'b0000000000001110;
    assign weights1[21][72] = 16'b0000000000001111;
    assign weights1[21][73] = 16'b1111111111110000;
    assign weights1[21][74] = 16'b0000000000000110;
    assign weights1[21][75] = 16'b1111111111111101;
    assign weights1[21][76] = 16'b1111111111111110;
    assign weights1[21][77] = 16'b0000000000000100;
    assign weights1[21][78] = 16'b0000000000000000;
    assign weights1[21][79] = 16'b1111111111111101;
    assign weights1[21][80] = 16'b1111111111111111;
    assign weights1[21][81] = 16'b1111111111111110;
    assign weights1[21][82] = 16'b1111111111111011;
    assign weights1[21][83] = 16'b1111111111111101;
    assign weights1[21][84] = 16'b1111111111111111;
    assign weights1[21][85] = 16'b1111111111111111;
    assign weights1[21][86] = 16'b1111111111111011;
    assign weights1[21][87] = 16'b1111111111110001;
    assign weights1[21][88] = 16'b1111111111101110;
    assign weights1[21][89] = 16'b1111111111101111;
    assign weights1[21][90] = 16'b1111111111111001;
    assign weights1[21][91] = 16'b1111111111110101;
    assign weights1[21][92] = 16'b1111111111101011;
    assign weights1[21][93] = 16'b1111111111111011;
    assign weights1[21][94] = 16'b1111111111110001;
    assign weights1[21][95] = 16'b1111111111110101;
    assign weights1[21][96] = 16'b1111111111100000;
    assign weights1[21][97] = 16'b1111111111110100;
    assign weights1[21][98] = 16'b1111111111100011;
    assign weights1[21][99] = 16'b1111111111110010;
    assign weights1[21][100] = 16'b0000000000000010;
    assign weights1[21][101] = 16'b1111111111101011;
    assign weights1[21][102] = 16'b1111111111110011;
    assign weights1[21][103] = 16'b1111111111111001;
    assign weights1[21][104] = 16'b1111111111101111;
    assign weights1[21][105] = 16'b1111111111110000;
    assign weights1[21][106] = 16'b1111111111110010;
    assign weights1[21][107] = 16'b0000000000000011;
    assign weights1[21][108] = 16'b1111111111111010;
    assign weights1[21][109] = 16'b1111111111110000;
    assign weights1[21][110] = 16'b1111111111110000;
    assign weights1[21][111] = 16'b0000000000000000;
    assign weights1[21][112] = 16'b0000000000000000;
    assign weights1[21][113] = 16'b0000000000000010;
    assign weights1[21][114] = 16'b1111111111111100;
    assign weights1[21][115] = 16'b1111111111110000;
    assign weights1[21][116] = 16'b1111111111101101;
    assign weights1[21][117] = 16'b1111111111111000;
    assign weights1[21][118] = 16'b0000000000001011;
    assign weights1[21][119] = 16'b0000000000000111;
    assign weights1[21][120] = 16'b0000000000010100;
    assign weights1[21][121] = 16'b0000000000000000;
    assign weights1[21][122] = 16'b1111111111101000;
    assign weights1[21][123] = 16'b1111111111110100;
    assign weights1[21][124] = 16'b1111111111111111;
    assign weights1[21][125] = 16'b1111111111110101;
    assign weights1[21][126] = 16'b0000000000011000;
    assign weights1[21][127] = 16'b0000000000000111;
    assign weights1[21][128] = 16'b0000000000001110;
    assign weights1[21][129] = 16'b0000000000001100;
    assign weights1[21][130] = 16'b0000000000001111;
    assign weights1[21][131] = 16'b0000000000000010;
    assign weights1[21][132] = 16'b0000000000000110;
    assign weights1[21][133] = 16'b0000000000000000;
    assign weights1[21][134] = 16'b1111111111101110;
    assign weights1[21][135] = 16'b0000000000000101;
    assign weights1[21][136] = 16'b1111111111111101;
    assign weights1[21][137] = 16'b1111111111100001;
    assign weights1[21][138] = 16'b1111111111111001;
    assign weights1[21][139] = 16'b1111111111110111;
    assign weights1[21][140] = 16'b0000000000000001;
    assign weights1[21][141] = 16'b1111111111111011;
    assign weights1[21][142] = 16'b1111111111110110;
    assign weights1[21][143] = 16'b1111111111101100;
    assign weights1[21][144] = 16'b1111111111110111;
    assign weights1[21][145] = 16'b1111111111110101;
    assign weights1[21][146] = 16'b0000000000010110;
    assign weights1[21][147] = 16'b0000000000001011;
    assign weights1[21][148] = 16'b0000000000100100;
    assign weights1[21][149] = 16'b0000000000011111;
    assign weights1[21][150] = 16'b1111111111111100;
    assign weights1[21][151] = 16'b0000000000010001;
    assign weights1[21][152] = 16'b1111111111111100;
    assign weights1[21][153] = 16'b1111111111110011;
    assign weights1[21][154] = 16'b0000000000010001;
    assign weights1[21][155] = 16'b1111111111110100;
    assign weights1[21][156] = 16'b1111111111111010;
    assign weights1[21][157] = 16'b0000000000000011;
    assign weights1[21][158] = 16'b0000000000000111;
    assign weights1[21][159] = 16'b1111111111110001;
    assign weights1[21][160] = 16'b1111111111111011;
    assign weights1[21][161] = 16'b0000000000001111;
    assign weights1[21][162] = 16'b0000000000000001;
    assign weights1[21][163] = 16'b0000000000010001;
    assign weights1[21][164] = 16'b0000000000001000;
    assign weights1[21][165] = 16'b1111111111110011;
    assign weights1[21][166] = 16'b1111111111111000;
    assign weights1[21][167] = 16'b1111111111101111;
    assign weights1[21][168] = 16'b0000000000000010;
    assign weights1[21][169] = 16'b0000000000000010;
    assign weights1[21][170] = 16'b0000000000000001;
    assign weights1[21][171] = 16'b1111111111110000;
    assign weights1[21][172] = 16'b1111111111111101;
    assign weights1[21][173] = 16'b0000000000001010;
    assign weights1[21][174] = 16'b1111111111111001;
    assign weights1[21][175] = 16'b0000000000010000;
    assign weights1[21][176] = 16'b0000000000010100;
    assign weights1[21][177] = 16'b0000000000101111;
    assign weights1[21][178] = 16'b0000000000000100;
    assign weights1[21][179] = 16'b1111111111110001;
    assign weights1[21][180] = 16'b0000000000001001;
    assign weights1[21][181] = 16'b1111111111111001;
    assign weights1[21][182] = 16'b1111111111111000;
    assign weights1[21][183] = 16'b0000000000001101;
    assign weights1[21][184] = 16'b0000000000001110;
    assign weights1[21][185] = 16'b0000000000010001;
    assign weights1[21][186] = 16'b1111111111111101;
    assign weights1[21][187] = 16'b0000000000000011;
    assign weights1[21][188] = 16'b1111111111111110;
    assign weights1[21][189] = 16'b1111111111111100;
    assign weights1[21][190] = 16'b0000000000010010;
    assign weights1[21][191] = 16'b1111111111111000;
    assign weights1[21][192] = 16'b1111111111111100;
    assign weights1[21][193] = 16'b0000000000000001;
    assign weights1[21][194] = 16'b0000000000001001;
    assign weights1[21][195] = 16'b0000000000000100;
    assign weights1[21][196] = 16'b0000000000000001;
    assign weights1[21][197] = 16'b0000000000000011;
    assign weights1[21][198] = 16'b0000000000000101;
    assign weights1[21][199] = 16'b1111111111111111;
    assign weights1[21][200] = 16'b1111111111111010;
    assign weights1[21][201] = 16'b1111111111111110;
    assign weights1[21][202] = 16'b0000000000000111;
    assign weights1[21][203] = 16'b0000000000000010;
    assign weights1[21][204] = 16'b1111111111111010;
    assign weights1[21][205] = 16'b0000000000011010;
    assign weights1[21][206] = 16'b0000000000011101;
    assign weights1[21][207] = 16'b0000000000010100;
    assign weights1[21][208] = 16'b1111111111111100;
    assign weights1[21][209] = 16'b0000000000010001;
    assign weights1[21][210] = 16'b1111111111100100;
    assign weights1[21][211] = 16'b0000000000001000;
    assign weights1[21][212] = 16'b1111111111111111;
    assign weights1[21][213] = 16'b1111111111111000;
    assign weights1[21][214] = 16'b0000000000010100;
    assign weights1[21][215] = 16'b0000000000100010;
    assign weights1[21][216] = 16'b0000000000000001;
    assign weights1[21][217] = 16'b1111111111101110;
    assign weights1[21][218] = 16'b0000000000001101;
    assign weights1[21][219] = 16'b1111111111111000;
    assign weights1[21][220] = 16'b0000000000010011;
    assign weights1[21][221] = 16'b0000000000001110;
    assign weights1[21][222] = 16'b0000000000000001;
    assign weights1[21][223] = 16'b0000000000000100;
    assign weights1[21][224] = 16'b0000000000000010;
    assign weights1[21][225] = 16'b0000000000000011;
    assign weights1[21][226] = 16'b1111111111111110;
    assign weights1[21][227] = 16'b1111111111111111;
    assign weights1[21][228] = 16'b1111111111111010;
    assign weights1[21][229] = 16'b0000000000011010;
    assign weights1[21][230] = 16'b1111111111110100;
    assign weights1[21][231] = 16'b1111111111101100;
    assign weights1[21][232] = 16'b0000000000001000;
    assign weights1[21][233] = 16'b0000000000011110;
    assign weights1[21][234] = 16'b0000000000011010;
    assign weights1[21][235] = 16'b0000000000010000;
    assign weights1[21][236] = 16'b0000000000010000;
    assign weights1[21][237] = 16'b0000000000000011;
    assign weights1[21][238] = 16'b0000000000000011;
    assign weights1[21][239] = 16'b1111111111111111;
    assign weights1[21][240] = 16'b0000000000000001;
    assign weights1[21][241] = 16'b0000000000001101;
    assign weights1[21][242] = 16'b0000000000000101;
    assign weights1[21][243] = 16'b0000000000000100;
    assign weights1[21][244] = 16'b0000000000001001;
    assign weights1[21][245] = 16'b1111111111111110;
    assign weights1[21][246] = 16'b0000000000000110;
    assign weights1[21][247] = 16'b0000000000000010;
    assign weights1[21][248] = 16'b1111111111110000;
    assign weights1[21][249] = 16'b1111111111111001;
    assign weights1[21][250] = 16'b0000000000001000;
    assign weights1[21][251] = 16'b0000000000000101;
    assign weights1[21][252] = 16'b1111111111111111;
    assign weights1[21][253] = 16'b0000000000000010;
    assign weights1[21][254] = 16'b0000000000001110;
    assign weights1[21][255] = 16'b1111111111111101;
    assign weights1[21][256] = 16'b0000000000000110;
    assign weights1[21][257] = 16'b0000000000010011;
    assign weights1[21][258] = 16'b0000000000011011;
    assign weights1[21][259] = 16'b0000000000100010;
    assign weights1[21][260] = 16'b0000000000011001;
    assign weights1[21][261] = 16'b0000000000000111;
    assign weights1[21][262] = 16'b0000000000000000;
    assign weights1[21][263] = 16'b0000000000101000;
    assign weights1[21][264] = 16'b0000000000010101;
    assign weights1[21][265] = 16'b0000000000000011;
    assign weights1[21][266] = 16'b1111111110011011;
    assign weights1[21][267] = 16'b1111111111101000;
    assign weights1[21][268] = 16'b1111111111111010;
    assign weights1[21][269] = 16'b1111111111111101;
    assign weights1[21][270] = 16'b0000000000001001;
    assign weights1[21][271] = 16'b0000000000000101;
    assign weights1[21][272] = 16'b1111111111111101;
    assign weights1[21][273] = 16'b1111111111111111;
    assign weights1[21][274] = 16'b1111111111111001;
    assign weights1[21][275] = 16'b1111111111110011;
    assign weights1[21][276] = 16'b1111111111111110;
    assign weights1[21][277] = 16'b1111111111111110;
    assign weights1[21][278] = 16'b1111111111110110;
    assign weights1[21][279] = 16'b1111111111110101;
    assign weights1[21][280] = 16'b0000000000000000;
    assign weights1[21][281] = 16'b0000000000000100;
    assign weights1[21][282] = 16'b0000000000001001;
    assign weights1[21][283] = 16'b0000000000001000;
    assign weights1[21][284] = 16'b1111111111110000;
    assign weights1[21][285] = 16'b0000000000000010;
    assign weights1[21][286] = 16'b0000000000000011;
    assign weights1[21][287] = 16'b1111111111101111;
    assign weights1[21][288] = 16'b0000000000100011;
    assign weights1[21][289] = 16'b0000000000010010;
    assign weights1[21][290] = 16'b0000000000011100;
    assign weights1[21][291] = 16'b1111111111101001;
    assign weights1[21][292] = 16'b0000000000001001;
    assign weights1[21][293] = 16'b1111111110001100;
    assign weights1[21][294] = 16'b1111111101100111;
    assign weights1[21][295] = 16'b1111111111010000;
    assign weights1[21][296] = 16'b1111111111111001;
    assign weights1[21][297] = 16'b0000000000001101;
    assign weights1[21][298] = 16'b1111111111111111;
    assign weights1[21][299] = 16'b1111111111110000;
    assign weights1[21][300] = 16'b1111111111110110;
    assign weights1[21][301] = 16'b1111111111111010;
    assign weights1[21][302] = 16'b0000000000000001;
    assign weights1[21][303] = 16'b1111111111110011;
    assign weights1[21][304] = 16'b1111111111111100;
    assign weights1[21][305] = 16'b1111111111110111;
    assign weights1[21][306] = 16'b1111111111101111;
    assign weights1[21][307] = 16'b1111111111101110;
    assign weights1[21][308] = 16'b0000000000000000;
    assign weights1[21][309] = 16'b0000000000001001;
    assign weights1[21][310] = 16'b0000000000001001;
    assign weights1[21][311] = 16'b1111111111110110;
    assign weights1[21][312] = 16'b1111111111110111;
    assign weights1[21][313] = 16'b1111111111110110;
    assign weights1[21][314] = 16'b0000000000101100;
    assign weights1[21][315] = 16'b0000000000000111;
    assign weights1[21][316] = 16'b0000000000001000;
    assign weights1[21][317] = 16'b0000000000001111;
    assign weights1[21][318] = 16'b0000000000010001;
    assign weights1[21][319] = 16'b0000000000001110;
    assign weights1[21][320] = 16'b1111111110011110;
    assign weights1[21][321] = 16'b1111111101000110;
    assign weights1[21][322] = 16'b1111111111001011;
    assign weights1[21][323] = 16'b1111111111101010;
    assign weights1[21][324] = 16'b1111111111110110;
    assign weights1[21][325] = 16'b0000000000000011;
    assign weights1[21][326] = 16'b1111111111111110;
    assign weights1[21][327] = 16'b0000000000001011;
    assign weights1[21][328] = 16'b1111111111110111;
    assign weights1[21][329] = 16'b1111111111111001;
    assign weights1[21][330] = 16'b1111111111111100;
    assign weights1[21][331] = 16'b0000000000000101;
    assign weights1[21][332] = 16'b0000000000001000;
    assign weights1[21][333] = 16'b1111111111110000;
    assign weights1[21][334] = 16'b1111111111110010;
    assign weights1[21][335] = 16'b1111111111101010;
    assign weights1[21][336] = 16'b0000000000000010;
    assign weights1[21][337] = 16'b0000000000000000;
    assign weights1[21][338] = 16'b1111111111110111;
    assign weights1[21][339] = 16'b0000000000000011;
    assign weights1[21][340] = 16'b1111111111111100;
    assign weights1[21][341] = 16'b1111111111111110;
    assign weights1[21][342] = 16'b0000000000000011;
    assign weights1[21][343] = 16'b0000000000001011;
    assign weights1[21][344] = 16'b0000000000011010;
    assign weights1[21][345] = 16'b0000000000001100;
    assign weights1[21][346] = 16'b1111111111100111;
    assign weights1[21][347] = 16'b1111111111001111;
    assign weights1[21][348] = 16'b1111111100110101;
    assign weights1[21][349] = 16'b1111111110000100;
    assign weights1[21][350] = 16'b0000000000010000;
    assign weights1[21][351] = 16'b1111111111111001;
    assign weights1[21][352] = 16'b0000000000001001;
    assign weights1[21][353] = 16'b0000000000001010;
    assign weights1[21][354] = 16'b1111111111110110;
    assign weights1[21][355] = 16'b0000000000000000;
    assign weights1[21][356] = 16'b1111111111110111;
    assign weights1[21][357] = 16'b1111111111110011;
    assign weights1[21][358] = 16'b1111111111110011;
    assign weights1[21][359] = 16'b0000000000000011;
    assign weights1[21][360] = 16'b1111111111101110;
    assign weights1[21][361] = 16'b1111111111100110;
    assign weights1[21][362] = 16'b1111111111101110;
    assign weights1[21][363] = 16'b1111111111101010;
    assign weights1[21][364] = 16'b1111111111111110;
    assign weights1[21][365] = 16'b1111111111110110;
    assign weights1[21][366] = 16'b1111111111111100;
    assign weights1[21][367] = 16'b1111111111110100;
    assign weights1[21][368] = 16'b1111111111110011;
    assign weights1[21][369] = 16'b1111111111110101;
    assign weights1[21][370] = 16'b0000000000000011;
    assign weights1[21][371] = 16'b1111111111101001;
    assign weights1[21][372] = 16'b1111111111110010;
    assign weights1[21][373] = 16'b1111111111001100;
    assign weights1[21][374] = 16'b1111111110100001;
    assign weights1[21][375] = 16'b1111111100101011;
    assign weights1[21][376] = 16'b1111111101111100;
    assign weights1[21][377] = 16'b0000000000000010;
    assign weights1[21][378] = 16'b1111111111011101;
    assign weights1[21][379] = 16'b1111111111111111;
    assign weights1[21][380] = 16'b0000000000000011;
    assign weights1[21][381] = 16'b0000000000001010;
    assign weights1[21][382] = 16'b1111111111110001;
    assign weights1[21][383] = 16'b1111111111101000;
    assign weights1[21][384] = 16'b1111111111110010;
    assign weights1[21][385] = 16'b1111111111110000;
    assign weights1[21][386] = 16'b1111111111010110;
    assign weights1[21][387] = 16'b1111111111011100;
    assign weights1[21][388] = 16'b1111111111100100;
    assign weights1[21][389] = 16'b1111111111101101;
    assign weights1[21][390] = 16'b1111111111101100;
    assign weights1[21][391] = 16'b1111111111101111;
    assign weights1[21][392] = 16'b1111111111110101;
    assign weights1[21][393] = 16'b1111111111110100;
    assign weights1[21][394] = 16'b1111111111100110;
    assign weights1[21][395] = 16'b1111111111101100;
    assign weights1[21][396] = 16'b1111111111010110;
    assign weights1[21][397] = 16'b1111111111011111;
    assign weights1[21][398] = 16'b1111111111001101;
    assign weights1[21][399] = 16'b1111111111001001;
    assign weights1[21][400] = 16'b1111111101111101;
    assign weights1[21][401] = 16'b1111111101110000;
    assign weights1[21][402] = 16'b1111111100110001;
    assign weights1[21][403] = 16'b1111111110110110;
    assign weights1[21][404] = 16'b1111111111101000;
    assign weights1[21][405] = 16'b1111111111110011;
    assign weights1[21][406] = 16'b1111111111111000;
    assign weights1[21][407] = 16'b1111111111110110;
    assign weights1[21][408] = 16'b0000000000000100;
    assign weights1[21][409] = 16'b0000000000010001;
    assign weights1[21][410] = 16'b0000000000001101;
    assign weights1[21][411] = 16'b0000000000000011;
    assign weights1[21][412] = 16'b1111111111101100;
    assign weights1[21][413] = 16'b1111111111100110;
    assign weights1[21][414] = 16'b1111111111101000;
    assign weights1[21][415] = 16'b1111111111010110;
    assign weights1[21][416] = 16'b1111111111100100;
    assign weights1[21][417] = 16'b1111111111100001;
    assign weights1[21][418] = 16'b1111111111100011;
    assign weights1[21][419] = 16'b1111111111101100;
    assign weights1[21][420] = 16'b1111111111101010;
    assign weights1[21][421] = 16'b1111111111100110;
    assign weights1[21][422] = 16'b1111111111100010;
    assign weights1[21][423] = 16'b1111111111001111;
    assign weights1[21][424] = 16'b1111111110111110;
    assign weights1[21][425] = 16'b1111111110110011;
    assign weights1[21][426] = 16'b1111111110010001;
    assign weights1[21][427] = 16'b1111111101101001;
    assign weights1[21][428] = 16'b1111111101001110;
    assign weights1[21][429] = 16'b1111111101010011;
    assign weights1[21][430] = 16'b1111111111000101;
    assign weights1[21][431] = 16'b1111111111100101;
    assign weights1[21][432] = 16'b1111111111110111;
    assign weights1[21][433] = 16'b1111111111111100;
    assign weights1[21][434] = 16'b0000000000000001;
    assign weights1[21][435] = 16'b0000000000000001;
    assign weights1[21][436] = 16'b0000000000000010;
    assign weights1[21][437] = 16'b0000000000000100;
    assign weights1[21][438] = 16'b0000000000010010;
    assign weights1[21][439] = 16'b0000000000010111;
    assign weights1[21][440] = 16'b1111111111110001;
    assign weights1[21][441] = 16'b1111111111101110;
    assign weights1[21][442] = 16'b1111111111100001;
    assign weights1[21][443] = 16'b1111111111110100;
    assign weights1[21][444] = 16'b1111111111101100;
    assign weights1[21][445] = 16'b1111111111011111;
    assign weights1[21][446] = 16'b1111111111101010;
    assign weights1[21][447] = 16'b1111111111101010;
    assign weights1[21][448] = 16'b1111111111101101;
    assign weights1[21][449] = 16'b1111111111011101;
    assign weights1[21][450] = 16'b1111111111010101;
    assign weights1[21][451] = 16'b1111111111001101;
    assign weights1[21][452] = 16'b1111111110110001;
    assign weights1[21][453] = 16'b1111111110100010;
    assign weights1[21][454] = 16'b1111111101111110;
    assign weights1[21][455] = 16'b1111111101111000;
    assign weights1[21][456] = 16'b1111111110010010;
    assign weights1[21][457] = 16'b1111111111111000;
    assign weights1[21][458] = 16'b0000000000000001;
    assign weights1[21][459] = 16'b0000000000001010;
    assign weights1[21][460] = 16'b0000000000000001;
    assign weights1[21][461] = 16'b0000000000001001;
    assign weights1[21][462] = 16'b1111111111111100;
    assign weights1[21][463] = 16'b0000000000000111;
    assign weights1[21][464] = 16'b0000000000001111;
    assign weights1[21][465] = 16'b0000000000011010;
    assign weights1[21][466] = 16'b0000000000000101;
    assign weights1[21][467] = 16'b1111111111100111;
    assign weights1[21][468] = 16'b1111111111011100;
    assign weights1[21][469] = 16'b1111111111100100;
    assign weights1[21][470] = 16'b1111111111110010;
    assign weights1[21][471] = 16'b0000000000000111;
    assign weights1[21][472] = 16'b0000000000000101;
    assign weights1[21][473] = 16'b1111111111111100;
    assign weights1[21][474] = 16'b1111111111110111;
    assign weights1[21][475] = 16'b1111111111111111;
    assign weights1[21][476] = 16'b1111111111101001;
    assign weights1[21][477] = 16'b1111111111011000;
    assign weights1[21][478] = 16'b1111111111001110;
    assign weights1[21][479] = 16'b1111111111001010;
    assign weights1[21][480] = 16'b1111111110110000;
    assign weights1[21][481] = 16'b1111111110110101;
    assign weights1[21][482] = 16'b1111111110111011;
    assign weights1[21][483] = 16'b1111111111010111;
    assign weights1[21][484] = 16'b0000000000010111;
    assign weights1[21][485] = 16'b0000000000101010;
    assign weights1[21][486] = 16'b0000000000000001;
    assign weights1[21][487] = 16'b0000000000100001;
    assign weights1[21][488] = 16'b1111111111111100;
    assign weights1[21][489] = 16'b0000000000000111;
    assign weights1[21][490] = 16'b1111111111111100;
    assign weights1[21][491] = 16'b0000000000010101;
    assign weights1[21][492] = 16'b1111111111111101;
    assign weights1[21][493] = 16'b1111111111110110;
    assign weights1[21][494] = 16'b0000000000000011;
    assign weights1[21][495] = 16'b1111111111101001;
    assign weights1[21][496] = 16'b1111111111101101;
    assign weights1[21][497] = 16'b1111111111101100;
    assign weights1[21][498] = 16'b0000000000000110;
    assign weights1[21][499] = 16'b0000000000011100;
    assign weights1[21][500] = 16'b0000000000011110;
    assign weights1[21][501] = 16'b0000000000000110;
    assign weights1[21][502] = 16'b0000000000010100;
    assign weights1[21][503] = 16'b0000000000000110;
    assign weights1[21][504] = 16'b1111111111100110;
    assign weights1[21][505] = 16'b1111111111011001;
    assign weights1[21][506] = 16'b1111111111001110;
    assign weights1[21][507] = 16'b1111111111001101;
    assign weights1[21][508] = 16'b1111111111010010;
    assign weights1[21][509] = 16'b1111111111000100;
    assign weights1[21][510] = 16'b1111111111101111;
    assign weights1[21][511] = 16'b0000000000100011;
    assign weights1[21][512] = 16'b0000000000010101;
    assign weights1[21][513] = 16'b0000000000000010;
    assign weights1[21][514] = 16'b0000000000000010;
    assign weights1[21][515] = 16'b1111111111111011;
    assign weights1[21][516] = 16'b0000000000000000;
    assign weights1[21][517] = 16'b0000000000000000;
    assign weights1[21][518] = 16'b0000000000001101;
    assign weights1[21][519] = 16'b0000000000000100;
    assign weights1[21][520] = 16'b0000000000000011;
    assign weights1[21][521] = 16'b0000000000000011;
    assign weights1[21][522] = 16'b1111111111111011;
    assign weights1[21][523] = 16'b1111111111110000;
    assign weights1[21][524] = 16'b0000000000000001;
    assign weights1[21][525] = 16'b0000000000011111;
    assign weights1[21][526] = 16'b1111111111111110;
    assign weights1[21][527] = 16'b1111111111110001;
    assign weights1[21][528] = 16'b0000000000001111;
    assign weights1[21][529] = 16'b0000000000010110;
    assign weights1[21][530] = 16'b0000000000001111;
    assign weights1[21][531] = 16'b0000000000001011;
    assign weights1[21][532] = 16'b1111111111101010;
    assign weights1[21][533] = 16'b1111111111011010;
    assign weights1[21][534] = 16'b1111111111010100;
    assign weights1[21][535] = 16'b1111111111010111;
    assign weights1[21][536] = 16'b1111111111011011;
    assign weights1[21][537] = 16'b1111111111101110;
    assign weights1[21][538] = 16'b1111111111110011;
    assign weights1[21][539] = 16'b0000000000001100;
    assign weights1[21][540] = 16'b1111111111110110;
    assign weights1[21][541] = 16'b0000000000011001;
    assign weights1[21][542] = 16'b1111111111111000;
    assign weights1[21][543] = 16'b0000000000011011;
    assign weights1[21][544] = 16'b0000000000001000;
    assign weights1[21][545] = 16'b0000000000000001;
    assign weights1[21][546] = 16'b0000000000000100;
    assign weights1[21][547] = 16'b1111111111110010;
    assign weights1[21][548] = 16'b0000000000000111;
    assign weights1[21][549] = 16'b1111111111101111;
    assign weights1[21][550] = 16'b1111111111101001;
    assign weights1[21][551] = 16'b0000000000001010;
    assign weights1[21][552] = 16'b0000000000001000;
    assign weights1[21][553] = 16'b1111111111110100;
    assign weights1[21][554] = 16'b0000000000010101;
    assign weights1[21][555] = 16'b0000000000001010;
    assign weights1[21][556] = 16'b0000000000010111;
    assign weights1[21][557] = 16'b0000000000010100;
    assign weights1[21][558] = 16'b0000000000010011;
    assign weights1[21][559] = 16'b0000000000000000;
    assign weights1[21][560] = 16'b1111111111110010;
    assign weights1[21][561] = 16'b1111111111100100;
    assign weights1[21][562] = 16'b1111111111100000;
    assign weights1[21][563] = 16'b1111111111010100;
    assign weights1[21][564] = 16'b1111111111011010;
    assign weights1[21][565] = 16'b1111111111101101;
    assign weights1[21][566] = 16'b0000000000000010;
    assign weights1[21][567] = 16'b1111111111111110;
    assign weights1[21][568] = 16'b0000000000011100;
    assign weights1[21][569] = 16'b0000000000001011;
    assign weights1[21][570] = 16'b0000000000010010;
    assign weights1[21][571] = 16'b0000000000010110;
    assign weights1[21][572] = 16'b0000000000010110;
    assign weights1[21][573] = 16'b0000000000000000;
    assign weights1[21][574] = 16'b1111111111110101;
    assign weights1[21][575] = 16'b1111111111111101;
    assign weights1[21][576] = 16'b1111111111101111;
    assign weights1[21][577] = 16'b1111111111101001;
    assign weights1[21][578] = 16'b1111111111111010;
    assign weights1[21][579] = 16'b1111111111110111;
    assign weights1[21][580] = 16'b1111111111111011;
    assign weights1[21][581] = 16'b0000000000001101;
    assign weights1[21][582] = 16'b1111111111111111;
    assign weights1[21][583] = 16'b0000000000000101;
    assign weights1[21][584] = 16'b0000000000010001;
    assign weights1[21][585] = 16'b0000000000001001;
    assign weights1[21][586] = 16'b0000000000000101;
    assign weights1[21][587] = 16'b0000000000000100;
    assign weights1[21][588] = 16'b1111111111110110;
    assign weights1[21][589] = 16'b1111111111101010;
    assign weights1[21][590] = 16'b1111111111110010;
    assign weights1[21][591] = 16'b1111111111110101;
    assign weights1[21][592] = 16'b1111111111111111;
    assign weights1[21][593] = 16'b0000000000011001;
    assign weights1[21][594] = 16'b1111111111101111;
    assign weights1[21][595] = 16'b0000000000001011;
    assign weights1[21][596] = 16'b0000000000010001;
    assign weights1[21][597] = 16'b0000000000010101;
    assign weights1[21][598] = 16'b0000000000010011;
    assign weights1[21][599] = 16'b0000000000010001;
    assign weights1[21][600] = 16'b1111111111111111;
    assign weights1[21][601] = 16'b0000000000000000;
    assign weights1[21][602] = 16'b1111111111011101;
    assign weights1[21][603] = 16'b1111111111101110;
    assign weights1[21][604] = 16'b1111111111100110;
    assign weights1[21][605] = 16'b1111111111110010;
    assign weights1[21][606] = 16'b1111111111110010;
    assign weights1[21][607] = 16'b1111111111111110;
    assign weights1[21][608] = 16'b1111111111101111;
    assign weights1[21][609] = 16'b0000000000010110;
    assign weights1[21][610] = 16'b0000000000001100;
    assign weights1[21][611] = 16'b0000000000001110;
    assign weights1[21][612] = 16'b0000000000000100;
    assign weights1[21][613] = 16'b0000000000001100;
    assign weights1[21][614] = 16'b0000000000000001;
    assign weights1[21][615] = 16'b0000000000000101;
    assign weights1[21][616] = 16'b1111111111111011;
    assign weights1[21][617] = 16'b1111111111111110;
    assign weights1[21][618] = 16'b0000000000000111;
    assign weights1[21][619] = 16'b0000000000011011;
    assign weights1[21][620] = 16'b0000000000000010;
    assign weights1[21][621] = 16'b0000000000010101;
    assign weights1[21][622] = 16'b1111111111111010;
    assign weights1[21][623] = 16'b0000000000001111;
    assign weights1[21][624] = 16'b0000000000001000;
    assign weights1[21][625] = 16'b0000000000000111;
    assign weights1[21][626] = 16'b1111111111110110;
    assign weights1[21][627] = 16'b1111111111111110;
    assign weights1[21][628] = 16'b1111111111111110;
    assign weights1[21][629] = 16'b1111111111110010;
    assign weights1[21][630] = 16'b0000000000010010;
    assign weights1[21][631] = 16'b1111111111100000;
    assign weights1[21][632] = 16'b1111111111110101;
    assign weights1[21][633] = 16'b0000000000001000;
    assign weights1[21][634] = 16'b1111111111110001;
    assign weights1[21][635] = 16'b0000000000000000;
    assign weights1[21][636] = 16'b1111111111110011;
    assign weights1[21][637] = 16'b0000000000000000;
    assign weights1[21][638] = 16'b0000000000000010;
    assign weights1[21][639] = 16'b0000000000000100;
    assign weights1[21][640] = 16'b1111111111111011;
    assign weights1[21][641] = 16'b1111111111110111;
    assign weights1[21][642] = 16'b0000000000000100;
    assign weights1[21][643] = 16'b0000000000000011;
    assign weights1[21][644] = 16'b0000000000000101;
    assign weights1[21][645] = 16'b0000000000000110;
    assign weights1[21][646] = 16'b0000000000100101;
    assign weights1[21][647] = 16'b0000000000000101;
    assign weights1[21][648] = 16'b1111111111111000;
    assign weights1[21][649] = 16'b0000000000001101;
    assign weights1[21][650] = 16'b0000000000010000;
    assign weights1[21][651] = 16'b0000000000011000;
    assign weights1[21][652] = 16'b0000000000001011;
    assign weights1[21][653] = 16'b1111111111110000;
    assign weights1[21][654] = 16'b0000000000011011;
    assign weights1[21][655] = 16'b1111111111101010;
    assign weights1[21][656] = 16'b1111111111110110;
    assign weights1[21][657] = 16'b0000000000001100;
    assign weights1[21][658] = 16'b1111111111011101;
    assign weights1[21][659] = 16'b1111111111110000;
    assign weights1[21][660] = 16'b1111111111101011;
    assign weights1[21][661] = 16'b1111111111011111;
    assign weights1[21][662] = 16'b1111111111110101;
    assign weights1[21][663] = 16'b1111111111110001;
    assign weights1[21][664] = 16'b1111111111111100;
    assign weights1[21][665] = 16'b1111111111111111;
    assign weights1[21][666] = 16'b1111111111111111;
    assign weights1[21][667] = 16'b1111111111111100;
    assign weights1[21][668] = 16'b0000000000000001;
    assign weights1[21][669] = 16'b1111111111111001;
    assign weights1[21][670] = 16'b1111111111111011;
    assign weights1[21][671] = 16'b0000000000000000;
    assign weights1[21][672] = 16'b0000000000000111;
    assign weights1[21][673] = 16'b0000000000001000;
    assign weights1[21][674] = 16'b0000000000011000;
    assign weights1[21][675] = 16'b0000000000001110;
    assign weights1[21][676] = 16'b0000000000011001;
    assign weights1[21][677] = 16'b0000000000011110;
    assign weights1[21][678] = 16'b1111111111111111;
    assign weights1[21][679] = 16'b1111111111111111;
    assign weights1[21][680] = 16'b1111111111111010;
    assign weights1[21][681] = 16'b0000000000001101;
    assign weights1[21][682] = 16'b1111111111101011;
    assign weights1[21][683] = 16'b1111111111011111;
    assign weights1[21][684] = 16'b0000000000010001;
    assign weights1[21][685] = 16'b0000000000001010;
    assign weights1[21][686] = 16'b1111111111110111;
    assign weights1[21][687] = 16'b0000000000001101;
    assign weights1[21][688] = 16'b1111111111101110;
    assign weights1[21][689] = 16'b1111111111101111;
    assign weights1[21][690] = 16'b1111111111010111;
    assign weights1[21][691] = 16'b1111111111100100;
    assign weights1[21][692] = 16'b1111111111110001;
    assign weights1[21][693] = 16'b1111111111110111;
    assign weights1[21][694] = 16'b1111111111111001;
    assign weights1[21][695] = 16'b1111111111101111;
    assign weights1[21][696] = 16'b1111111111111011;
    assign weights1[21][697] = 16'b1111111111111010;
    assign weights1[21][698] = 16'b1111111111111000;
    assign weights1[21][699] = 16'b1111111111111111;
    assign weights1[21][700] = 16'b0000000000000111;
    assign weights1[21][701] = 16'b0000000000010001;
    assign weights1[21][702] = 16'b0000000000001110;
    assign weights1[21][703] = 16'b0000000000010001;
    assign weights1[21][704] = 16'b0000000000100100;
    assign weights1[21][705] = 16'b0000000000010010;
    assign weights1[21][706] = 16'b0000000000000010;
    assign weights1[21][707] = 16'b0000000000001010;
    assign weights1[21][708] = 16'b0000000000000111;
    assign weights1[21][709] = 16'b0000000000001101;
    assign weights1[21][710] = 16'b1111111111101111;
    assign weights1[21][711] = 16'b0000000000010010;
    assign weights1[21][712] = 16'b1111111111111110;
    assign weights1[21][713] = 16'b0000000000001100;
    assign weights1[21][714] = 16'b1111111111101000;
    assign weights1[21][715] = 16'b0000000000001110;
    assign weights1[21][716] = 16'b1111111111100101;
    assign weights1[21][717] = 16'b1111111111110111;
    assign weights1[21][718] = 16'b1111111111110011;
    assign weights1[21][719] = 16'b1111111111010110;
    assign weights1[21][720] = 16'b1111111111100000;
    assign weights1[21][721] = 16'b1111111111110010;
    assign weights1[21][722] = 16'b1111111111101101;
    assign weights1[21][723] = 16'b1111111111101110;
    assign weights1[21][724] = 16'b1111111111101011;
    assign weights1[21][725] = 16'b1111111111110101;
    assign weights1[21][726] = 16'b1111111111111000;
    assign weights1[21][727] = 16'b1111111111111111;
    assign weights1[21][728] = 16'b0000000000000101;
    assign weights1[21][729] = 16'b0000000000001110;
    assign weights1[21][730] = 16'b0000000000000110;
    assign weights1[21][731] = 16'b0000000000001001;
    assign weights1[21][732] = 16'b0000000000010101;
    assign weights1[21][733] = 16'b0000000000000011;
    assign weights1[21][734] = 16'b1111111111110101;
    assign weights1[21][735] = 16'b0000000000000111;
    assign weights1[21][736] = 16'b1111111111110011;
    assign weights1[21][737] = 16'b1111111111111001;
    assign weights1[21][738] = 16'b1111111111111100;
    assign weights1[21][739] = 16'b1111111111111001;
    assign weights1[21][740] = 16'b1111111111111100;
    assign weights1[21][741] = 16'b0000000000001111;
    assign weights1[21][742] = 16'b1111111111111001;
    assign weights1[21][743] = 16'b1111111111110111;
    assign weights1[21][744] = 16'b0000000000001110;
    assign weights1[21][745] = 16'b1111111111111111;
    assign weights1[21][746] = 16'b1111111111111000;
    assign weights1[21][747] = 16'b1111111111111100;
    assign weights1[21][748] = 16'b1111111111101111;
    assign weights1[21][749] = 16'b1111111111101110;
    assign weights1[21][750] = 16'b1111111111110100;
    assign weights1[21][751] = 16'b1111111111101101;
    assign weights1[21][752] = 16'b1111111111110100;
    assign weights1[21][753] = 16'b1111111111111110;
    assign weights1[21][754] = 16'b1111111111111111;
    assign weights1[21][755] = 16'b0000000000000000;
    assign weights1[21][756] = 16'b0000000000000011;
    assign weights1[21][757] = 16'b0000000000001001;
    assign weights1[21][758] = 16'b0000000000001110;
    assign weights1[21][759] = 16'b0000000000010001;
    assign weights1[21][760] = 16'b0000000000010001;
    assign weights1[21][761] = 16'b0000000000001100;
    assign weights1[21][762] = 16'b0000000000000000;
    assign weights1[21][763] = 16'b1111111111100100;
    assign weights1[21][764] = 16'b1111111111100011;
    assign weights1[21][765] = 16'b1111111111110100;
    assign weights1[21][766] = 16'b1111111111100101;
    assign weights1[21][767] = 16'b1111111111011100;
    assign weights1[21][768] = 16'b1111111111101011;
    assign weights1[21][769] = 16'b1111111111111101;
    assign weights1[21][770] = 16'b1111111111110100;
    assign weights1[21][771] = 16'b1111111111101010;
    assign weights1[21][772] = 16'b1111111111110010;
    assign weights1[21][773] = 16'b1111111111101111;
    assign weights1[21][774] = 16'b0000000000000011;
    assign weights1[21][775] = 16'b1111111111111101;
    assign weights1[21][776] = 16'b0000000000000011;
    assign weights1[21][777] = 16'b1111111111111101;
    assign weights1[21][778] = 16'b1111111111110100;
    assign weights1[21][779] = 16'b1111111111110111;
    assign weights1[21][780] = 16'b1111111111111011;
    assign weights1[21][781] = 16'b0000000000000010;
    assign weights1[21][782] = 16'b0000000000000000;
    assign weights1[21][783] = 16'b0000000000000001;
    assign weights1[22][0] = 16'b0000000000000000;
    assign weights1[22][1] = 16'b0000000000000001;
    assign weights1[22][2] = 16'b0000000000000000;
    assign weights1[22][3] = 16'b0000000000000001;
    assign weights1[22][4] = 16'b0000000000001101;
    assign weights1[22][5] = 16'b0000000000011101;
    assign weights1[22][6] = 16'b0000000000100011;
    assign weights1[22][7] = 16'b0000000000101110;
    assign weights1[22][8] = 16'b0000000000101011;
    assign weights1[22][9] = 16'b0000000000011101;
    assign weights1[22][10] = 16'b0000000000011110;
    assign weights1[22][11] = 16'b0000000000010111;
    assign weights1[22][12] = 16'b0000000000011100;
    assign weights1[22][13] = 16'b0000000000100111;
    assign weights1[22][14] = 16'b0000000000100001;
    assign weights1[22][15] = 16'b0000000000100000;
    assign weights1[22][16] = 16'b0000000000000111;
    assign weights1[22][17] = 16'b0000000000001110;
    assign weights1[22][18] = 16'b0000000000010010;
    assign weights1[22][19] = 16'b1111111111111111;
    assign weights1[22][20] = 16'b0000000000000101;
    assign weights1[22][21] = 16'b0000000000000110;
    assign weights1[22][22] = 16'b0000000000001001;
    assign weights1[22][23] = 16'b0000000000001000;
    assign weights1[22][24] = 16'b0000000000000100;
    assign weights1[22][25] = 16'b1111111111111011;
    assign weights1[22][26] = 16'b1111111111111011;
    assign weights1[22][27] = 16'b1111111111111011;
    assign weights1[22][28] = 16'b1111111111111111;
    assign weights1[22][29] = 16'b0000000000000001;
    assign weights1[22][30] = 16'b0000000000000011;
    assign weights1[22][31] = 16'b0000000000001110;
    assign weights1[22][32] = 16'b0000000000011111;
    assign weights1[22][33] = 16'b0000000000010100;
    assign weights1[22][34] = 16'b0000000000100011;
    assign weights1[22][35] = 16'b0000000000011111;
    assign weights1[22][36] = 16'b0000000000011101;
    assign weights1[22][37] = 16'b0000000000001001;
    assign weights1[22][38] = 16'b0000000000000000;
    assign weights1[22][39] = 16'b0000000000001000;
    assign weights1[22][40] = 16'b1111111111101100;
    assign weights1[22][41] = 16'b1111111111111000;
    assign weights1[22][42] = 16'b1111111111111101;
    assign weights1[22][43] = 16'b1111111111111100;
    assign weights1[22][44] = 16'b1111111111111010;
    assign weights1[22][45] = 16'b1111111111111001;
    assign weights1[22][46] = 16'b1111111111111111;
    assign weights1[22][47] = 16'b0000000000000100;
    assign weights1[22][48] = 16'b0000000000001001;
    assign weights1[22][49] = 16'b0000000000001000;
    assign weights1[22][50] = 16'b1111111111110010;
    assign weights1[22][51] = 16'b0000000000000000;
    assign weights1[22][52] = 16'b0000000000000100;
    assign weights1[22][53] = 16'b0000000000000101;
    assign weights1[22][54] = 16'b1111111111111110;
    assign weights1[22][55] = 16'b0000000000000011;
    assign weights1[22][56] = 16'b0000000000000001;
    assign weights1[22][57] = 16'b0000000000000111;
    assign weights1[22][58] = 16'b0000000000001011;
    assign weights1[22][59] = 16'b0000000000011011;
    assign weights1[22][60] = 16'b0000000000011101;
    assign weights1[22][61] = 16'b0000000000011001;
    assign weights1[22][62] = 16'b0000000000100010;
    assign weights1[22][63] = 16'b0000000000100111;
    assign weights1[22][64] = 16'b0000000000100101;
    assign weights1[22][65] = 16'b0000000000100110;
    assign weights1[22][66] = 16'b0000000000010011;
    assign weights1[22][67] = 16'b0000000000001001;
    assign weights1[22][68] = 16'b0000000000010001;
    assign weights1[22][69] = 16'b1111111111111110;
    assign weights1[22][70] = 16'b1111111111101110;
    assign weights1[22][71] = 16'b1111111111110110;
    assign weights1[22][72] = 16'b0000000000000111;
    assign weights1[22][73] = 16'b1111111111111110;
    assign weights1[22][74] = 16'b1111111111110011;
    assign weights1[22][75] = 16'b0000000000000110;
    assign weights1[22][76] = 16'b1111111111111110;
    assign weights1[22][77] = 16'b0000000000000011;
    assign weights1[22][78] = 16'b0000000000000100;
    assign weights1[22][79] = 16'b0000000000000111;
    assign weights1[22][80] = 16'b0000000000010010;
    assign weights1[22][81] = 16'b1111111111111100;
    assign weights1[22][82] = 16'b1111111111101110;
    assign weights1[22][83] = 16'b1111111111111000;
    assign weights1[22][84] = 16'b0000000000000010;
    assign weights1[22][85] = 16'b0000000000001100;
    assign weights1[22][86] = 16'b0000000000001000;
    assign weights1[22][87] = 16'b0000000000011100;
    assign weights1[22][88] = 16'b0000000000011100;
    assign weights1[22][89] = 16'b0000000000100011;
    assign weights1[22][90] = 16'b0000000000100101;
    assign weights1[22][91] = 16'b0000000000111101;
    assign weights1[22][92] = 16'b0000000001000101;
    assign weights1[22][93] = 16'b0000000000101011;
    assign weights1[22][94] = 16'b0000000000110000;
    assign weights1[22][95] = 16'b0000000000011010;
    assign weights1[22][96] = 16'b0000000000000110;
    assign weights1[22][97] = 16'b0000000000101100;
    assign weights1[22][98] = 16'b0000000000011001;
    assign weights1[22][99] = 16'b1111111111111111;
    assign weights1[22][100] = 16'b0000000000010011;
    assign weights1[22][101] = 16'b0000000000010000;
    assign weights1[22][102] = 16'b0000000000000100;
    assign weights1[22][103] = 16'b1111111111111100;
    assign weights1[22][104] = 16'b1111111111110111;
    assign weights1[22][105] = 16'b0000000000000000;
    assign weights1[22][106] = 16'b1111111111110001;
    assign weights1[22][107] = 16'b0000000000001001;
    assign weights1[22][108] = 16'b0000000000010000;
    assign weights1[22][109] = 16'b1111111111110101;
    assign weights1[22][110] = 16'b0000000000000000;
    assign weights1[22][111] = 16'b1111111111111000;
    assign weights1[22][112] = 16'b0000000000000110;
    assign weights1[22][113] = 16'b0000000000001100;
    assign weights1[22][114] = 16'b0000000000000110;
    assign weights1[22][115] = 16'b0000000000011000;
    assign weights1[22][116] = 16'b0000000000100110;
    assign weights1[22][117] = 16'b0000000000110001;
    assign weights1[22][118] = 16'b0000000001000101;
    assign weights1[22][119] = 16'b0000000000111100;
    assign weights1[22][120] = 16'b0000000000101101;
    assign weights1[22][121] = 16'b0000000000110010;
    assign weights1[22][122] = 16'b0000000001000001;
    assign weights1[22][123] = 16'b0000000000011110;
    assign weights1[22][124] = 16'b0000000000011010;
    assign weights1[22][125] = 16'b0000000000000110;
    assign weights1[22][126] = 16'b0000000000001010;
    assign weights1[22][127] = 16'b0000000000010001;
    assign weights1[22][128] = 16'b0000000000010001;
    assign weights1[22][129] = 16'b0000000000000101;
    assign weights1[22][130] = 16'b0000000000000101;
    assign weights1[22][131] = 16'b0000000000001111;
    assign weights1[22][132] = 16'b0000000000010011;
    assign weights1[22][133] = 16'b0000000000000001;
    assign weights1[22][134] = 16'b0000000000000000;
    assign weights1[22][135] = 16'b1111111111110101;
    assign weights1[22][136] = 16'b0000000000000100;
    assign weights1[22][137] = 16'b0000000000000001;
    assign weights1[22][138] = 16'b0000000000000000;
    assign weights1[22][139] = 16'b0000000000000001;
    assign weights1[22][140] = 16'b0000000000000010;
    assign weights1[22][141] = 16'b0000000000000001;
    assign weights1[22][142] = 16'b0000000000000010;
    assign weights1[22][143] = 16'b0000000000011110;
    assign weights1[22][144] = 16'b0000000000110010;
    assign weights1[22][145] = 16'b0000000000100111;
    assign weights1[22][146] = 16'b0000000000111101;
    assign weights1[22][147] = 16'b0000000001000111;
    assign weights1[22][148] = 16'b0000000000110100;
    assign weights1[22][149] = 16'b0000000000100110;
    assign weights1[22][150] = 16'b0000000000101110;
    assign weights1[22][151] = 16'b0000000001001101;
    assign weights1[22][152] = 16'b0000000000110011;
    assign weights1[22][153] = 16'b0000000000011001;
    assign weights1[22][154] = 16'b0000000000010101;
    assign weights1[22][155] = 16'b0000000000010001;
    assign weights1[22][156] = 16'b0000000000000111;
    assign weights1[22][157] = 16'b0000000000000101;
    assign weights1[22][158] = 16'b0000000000010100;
    assign weights1[22][159] = 16'b0000000000001010;
    assign weights1[22][160] = 16'b0000000000001000;
    assign weights1[22][161] = 16'b1111111111111111;
    assign weights1[22][162] = 16'b0000000000001010;
    assign weights1[22][163] = 16'b0000000000000101;
    assign weights1[22][164] = 16'b0000000000001010;
    assign weights1[22][165] = 16'b0000000000000111;
    assign weights1[22][166] = 16'b1111111111111001;
    assign weights1[22][167] = 16'b1111111111111110;
    assign weights1[22][168] = 16'b1111111111111100;
    assign weights1[22][169] = 16'b1111111111111101;
    assign weights1[22][170] = 16'b1111111111110111;
    assign weights1[22][171] = 16'b0000000000010000;
    assign weights1[22][172] = 16'b0000000000101100;
    assign weights1[22][173] = 16'b0000000000101000;
    assign weights1[22][174] = 16'b0000000000011100;
    assign weights1[22][175] = 16'b0000000001010101;
    assign weights1[22][176] = 16'b0000000001010011;
    assign weights1[22][177] = 16'b0000000001011101;
    assign weights1[22][178] = 16'b0000000000111011;
    assign weights1[22][179] = 16'b0000000001010001;
    assign weights1[22][180] = 16'b0000000001001001;
    assign weights1[22][181] = 16'b0000000000110110;
    assign weights1[22][182] = 16'b0000000000100101;
    assign weights1[22][183] = 16'b0000000000100011;
    assign weights1[22][184] = 16'b0000000000011101;
    assign weights1[22][185] = 16'b0000000000000100;
    assign weights1[22][186] = 16'b0000000000000101;
    assign weights1[22][187] = 16'b0000000000001100;
    assign weights1[22][188] = 16'b0000000000000111;
    assign weights1[22][189] = 16'b0000000000001001;
    assign weights1[22][190] = 16'b0000000000000110;
    assign weights1[22][191] = 16'b0000000000001100;
    assign weights1[22][192] = 16'b0000000000000011;
    assign weights1[22][193] = 16'b0000000000000101;
    assign weights1[22][194] = 16'b1111111111111101;
    assign weights1[22][195] = 16'b0000000000000010;
    assign weights1[22][196] = 16'b1111111111100111;
    assign weights1[22][197] = 16'b1111111111100001;
    assign weights1[22][198] = 16'b1111111111011100;
    assign weights1[22][199] = 16'b1111111111101000;
    assign weights1[22][200] = 16'b1111111111111111;
    assign weights1[22][201] = 16'b0000000000010001;
    assign weights1[22][202] = 16'b0000000000011110;
    assign weights1[22][203] = 16'b0000000000011011;
    assign weights1[22][204] = 16'b0000000000100101;
    assign weights1[22][205] = 16'b0000000000000110;
    assign weights1[22][206] = 16'b0000000000010101;
    assign weights1[22][207] = 16'b0000000000000011;
    assign weights1[22][208] = 16'b0000000000001011;
    assign weights1[22][209] = 16'b0000000000010111;
    assign weights1[22][210] = 16'b0000000000100010;
    assign weights1[22][211] = 16'b0000000000001010;
    assign weights1[22][212] = 16'b0000000000100011;
    assign weights1[22][213] = 16'b1111111111111111;
    assign weights1[22][214] = 16'b0000000000001111;
    assign weights1[22][215] = 16'b1111111111111100;
    assign weights1[22][216] = 16'b0000000000000100;
    assign weights1[22][217] = 16'b0000000000001001;
    assign weights1[22][218] = 16'b0000000000001101;
    assign weights1[22][219] = 16'b1111111111110101;
    assign weights1[22][220] = 16'b0000000000001110;
    assign weights1[22][221] = 16'b0000000000000111;
    assign weights1[22][222] = 16'b1111111111111111;
    assign weights1[22][223] = 16'b1111111111110110;
    assign weights1[22][224] = 16'b1111111111011111;
    assign weights1[22][225] = 16'b1111111111000111;
    assign weights1[22][226] = 16'b1111111110011110;
    assign weights1[22][227] = 16'b1111111110011000;
    assign weights1[22][228] = 16'b1111111110001011;
    assign weights1[22][229] = 16'b1111111110010111;
    assign weights1[22][230] = 16'b1111111110111111;
    assign weights1[22][231] = 16'b1111111110011110;
    assign weights1[22][232] = 16'b1111111110101001;
    assign weights1[22][233] = 16'b1111111110010001;
    assign weights1[22][234] = 16'b1111111110110000;
    assign weights1[22][235] = 16'b1111111110111110;
    assign weights1[22][236] = 16'b1111111110111111;
    assign weights1[22][237] = 16'b1111111111001000;
    assign weights1[22][238] = 16'b1111111111000111;
    assign weights1[22][239] = 16'b1111111111010110;
    assign weights1[22][240] = 16'b1111111111101001;
    assign weights1[22][241] = 16'b1111111111111010;
    assign weights1[22][242] = 16'b0000000000001001;
    assign weights1[22][243] = 16'b1111111111110011;
    assign weights1[22][244] = 16'b1111111111111111;
    assign weights1[22][245] = 16'b1111111111111110;
    assign weights1[22][246] = 16'b0000000000001010;
    assign weights1[22][247] = 16'b0000000000000011;
    assign weights1[22][248] = 16'b1111111111111011;
    assign weights1[22][249] = 16'b0000000000000001;
    assign weights1[22][250] = 16'b1111111111111011;
    assign weights1[22][251] = 16'b0000000000000100;
    assign weights1[22][252] = 16'b1111111111001100;
    assign weights1[22][253] = 16'b1111111110011001;
    assign weights1[22][254] = 16'b1111111101111011;
    assign weights1[22][255] = 16'b1111111101100001;
    assign weights1[22][256] = 16'b1111111101010101;
    assign weights1[22][257] = 16'b1111111100110101;
    assign weights1[22][258] = 16'b1111111100001100;
    assign weights1[22][259] = 16'b1111111011101100;
    assign weights1[22][260] = 16'b1111111011101111;
    assign weights1[22][261] = 16'b1111111100000000;
    assign weights1[22][262] = 16'b1111111100011101;
    assign weights1[22][263] = 16'b1111111100111100;
    assign weights1[22][264] = 16'b1111111101110100;
    assign weights1[22][265] = 16'b1111111110011001;
    assign weights1[22][266] = 16'b1111111111000011;
    assign weights1[22][267] = 16'b1111111111001111;
    assign weights1[22][268] = 16'b1111111111011000;
    assign weights1[22][269] = 16'b1111111111100111;
    assign weights1[22][270] = 16'b1111111111111000;
    assign weights1[22][271] = 16'b1111111111110001;
    assign weights1[22][272] = 16'b0000000000001100;
    assign weights1[22][273] = 16'b1111111111100100;
    assign weights1[22][274] = 16'b0000000000000101;
    assign weights1[22][275] = 16'b0000000000000110;
    assign weights1[22][276] = 16'b0000000000000011;
    assign weights1[22][277] = 16'b0000000000000001;
    assign weights1[22][278] = 16'b1111111111111100;
    assign weights1[22][279] = 16'b1111111111101001;
    assign weights1[22][280] = 16'b1111111110111011;
    assign weights1[22][281] = 16'b1111111101111011;
    assign weights1[22][282] = 16'b1111111101100000;
    assign weights1[22][283] = 16'b1111111101001011;
    assign weights1[22][284] = 16'b1111111100101110;
    assign weights1[22][285] = 16'b1111111011111010;
    assign weights1[22][286] = 16'b1111111011110111;
    assign weights1[22][287] = 16'b1111111011111010;
    assign weights1[22][288] = 16'b1111111100011011;
    assign weights1[22][289] = 16'b1111111110000001;
    assign weights1[22][290] = 16'b1111111110111000;
    assign weights1[22][291] = 16'b1111111111010110;
    assign weights1[22][292] = 16'b1111111111101000;
    assign weights1[22][293] = 16'b1111111111101110;
    assign weights1[22][294] = 16'b1111111111101011;
    assign weights1[22][295] = 16'b1111111111101101;
    assign weights1[22][296] = 16'b1111111111110111;
    assign weights1[22][297] = 16'b1111111111101001;
    assign weights1[22][298] = 16'b1111111111110101;
    assign weights1[22][299] = 16'b1111111111111001;
    assign weights1[22][300] = 16'b1111111111111001;
    assign weights1[22][301] = 16'b0000000000001100;
    assign weights1[22][302] = 16'b1111111111111001;
    assign weights1[22][303] = 16'b1111111111111100;
    assign weights1[22][304] = 16'b0000000000010100;
    assign weights1[22][305] = 16'b1111111111110111;
    assign weights1[22][306] = 16'b0000000000000110;
    assign weights1[22][307] = 16'b1111111111110000;
    assign weights1[22][308] = 16'b1111111111000000;
    assign weights1[22][309] = 16'b1111111110010100;
    assign weights1[22][310] = 16'b1111111101110011;
    assign weights1[22][311] = 16'b1111111101110000;
    assign weights1[22][312] = 16'b1111111101110010;
    assign weights1[22][313] = 16'b1111111110000111;
    assign weights1[22][314] = 16'b1111111110100110;
    assign weights1[22][315] = 16'b1111111111010111;
    assign weights1[22][316] = 16'b1111111111111101;
    assign weights1[22][317] = 16'b1111111111111110;
    assign weights1[22][318] = 16'b1111111111110111;
    assign weights1[22][319] = 16'b0000000000000000;
    assign weights1[22][320] = 16'b1111111111111000;
    assign weights1[22][321] = 16'b1111111111111001;
    assign weights1[22][322] = 16'b1111111111111011;
    assign weights1[22][323] = 16'b0000000000000010;
    assign weights1[22][324] = 16'b0000000000000010;
    assign weights1[22][325] = 16'b0000000000010101;
    assign weights1[22][326] = 16'b1111111111111011;
    assign weights1[22][327] = 16'b0000000000000010;
    assign weights1[22][328] = 16'b0000000000001100;
    assign weights1[22][329] = 16'b0000000000000000;
    assign weights1[22][330] = 16'b1111111111110010;
    assign weights1[22][331] = 16'b0000000000001000;
    assign weights1[22][332] = 16'b1111111111111101;
    assign weights1[22][333] = 16'b1111111111111100;
    assign weights1[22][334] = 16'b1111111111100111;
    assign weights1[22][335] = 16'b1111111111110001;
    assign weights1[22][336] = 16'b1111111111010100;
    assign weights1[22][337] = 16'b1111111110110010;
    assign weights1[22][338] = 16'b1111111111001000;
    assign weights1[22][339] = 16'b1111111111001010;
    assign weights1[22][340] = 16'b1111111111101011;
    assign weights1[22][341] = 16'b1111111111110110;
    assign weights1[22][342] = 16'b0000000000011101;
    assign weights1[22][343] = 16'b0000000000100111;
    assign weights1[22][344] = 16'b0000000000111001;
    assign weights1[22][345] = 16'b0000000000100001;
    assign weights1[22][346] = 16'b0000000000011110;
    assign weights1[22][347] = 16'b0000000000010111;
    assign weights1[22][348] = 16'b0000000000010001;
    assign weights1[22][349] = 16'b0000000000000110;
    assign weights1[22][350] = 16'b0000000000001010;
    assign weights1[22][351] = 16'b0000000000000100;
    assign weights1[22][352] = 16'b0000000000001000;
    assign weights1[22][353] = 16'b1111111111110010;
    assign weights1[22][354] = 16'b0000000000001100;
    assign weights1[22][355] = 16'b1111111111110100;
    assign weights1[22][356] = 16'b1111111111111111;
    assign weights1[22][357] = 16'b1111111111110111;
    assign weights1[22][358] = 16'b0000000000010011;
    assign weights1[22][359] = 16'b0000000000000001;
    assign weights1[22][360] = 16'b1111111111101110;
    assign weights1[22][361] = 16'b0000000000010010;
    assign weights1[22][362] = 16'b0000000000000010;
    assign weights1[22][363] = 16'b0000000000000011;
    assign weights1[22][364] = 16'b1111111111101110;
    assign weights1[22][365] = 16'b1111111111111011;
    assign weights1[22][366] = 16'b0000000000000101;
    assign weights1[22][367] = 16'b0000000000010011;
    assign weights1[22][368] = 16'b0000000000111010;
    assign weights1[22][369] = 16'b0000000000100101;
    assign weights1[22][370] = 16'b0000000000100000;
    assign weights1[22][371] = 16'b0000000000011100;
    assign weights1[22][372] = 16'b0000000000100000;
    assign weights1[22][373] = 16'b0000000000001100;
    assign weights1[22][374] = 16'b0000000000001111;
    assign weights1[22][375] = 16'b0000000000010001;
    assign weights1[22][376] = 16'b0000000000011000;
    assign weights1[22][377] = 16'b0000000000011110;
    assign weights1[22][378] = 16'b0000000000001000;
    assign weights1[22][379] = 16'b0000000000010001;
    assign weights1[22][380] = 16'b0000000000001001;
    assign weights1[22][381] = 16'b0000000000000010;
    assign weights1[22][382] = 16'b1111111111111011;
    assign weights1[22][383] = 16'b0000000000001100;
    assign weights1[22][384] = 16'b0000000000000001;
    assign weights1[22][385] = 16'b0000000000000000;
    assign weights1[22][386] = 16'b0000000000001001;
    assign weights1[22][387] = 16'b0000000000000000;
    assign weights1[22][388] = 16'b1111111111111110;
    assign weights1[22][389] = 16'b1111111111111010;
    assign weights1[22][390] = 16'b0000000000001001;
    assign weights1[22][391] = 16'b1111111111111000;
    assign weights1[22][392] = 16'b1111111111111011;
    assign weights1[22][393] = 16'b0000000000100101;
    assign weights1[22][394] = 16'b0000000000011010;
    assign weights1[22][395] = 16'b0000000000111001;
    assign weights1[22][396] = 16'b0000000000111001;
    assign weights1[22][397] = 16'b0000000000110000;
    assign weights1[22][398] = 16'b0000000000101001;
    assign weights1[22][399] = 16'b0000000000011100;
    assign weights1[22][400] = 16'b0000000000011111;
    assign weights1[22][401] = 16'b0000000000010110;
    assign weights1[22][402] = 16'b0000000000000000;
    assign weights1[22][403] = 16'b0000000000010100;
    assign weights1[22][404] = 16'b1111111111111010;
    assign weights1[22][405] = 16'b0000000000000001;
    assign weights1[22][406] = 16'b1111111111111100;
    assign weights1[22][407] = 16'b0000000000001001;
    assign weights1[22][408] = 16'b0000000000001011;
    assign weights1[22][409] = 16'b1111111111111001;
    assign weights1[22][410] = 16'b0000000000010010;
    assign weights1[22][411] = 16'b1111111111111101;
    assign weights1[22][412] = 16'b0000000000001111;
    assign weights1[22][413] = 16'b1111111111111110;
    assign weights1[22][414] = 16'b1111111111101110;
    assign weights1[22][415] = 16'b0000000000000011;
    assign weights1[22][416] = 16'b1111111111111010;
    assign weights1[22][417] = 16'b1111111111111100;
    assign weights1[22][418] = 16'b0000000000000001;
    assign weights1[22][419] = 16'b0000000000000011;
    assign weights1[22][420] = 16'b0000000000001101;
    assign weights1[22][421] = 16'b0000000000100010;
    assign weights1[22][422] = 16'b0000000000100001;
    assign weights1[22][423] = 16'b0000000000001100;
    assign weights1[22][424] = 16'b0000000000000000;
    assign weights1[22][425] = 16'b0000000000010011;
    assign weights1[22][426] = 16'b0000000000000111;
    assign weights1[22][427] = 16'b1111111111110101;
    assign weights1[22][428] = 16'b1111111111111011;
    assign weights1[22][429] = 16'b0000000000000111;
    assign weights1[22][430] = 16'b0000000000001010;
    assign weights1[22][431] = 16'b0000000000000011;
    assign weights1[22][432] = 16'b0000000000010010;
    assign weights1[22][433] = 16'b0000000000000100;
    assign weights1[22][434] = 16'b0000000000001000;
    assign weights1[22][435] = 16'b0000000000000010;
    assign weights1[22][436] = 16'b0000000000001111;
    assign weights1[22][437] = 16'b0000000000000011;
    assign weights1[22][438] = 16'b1111111111110111;
    assign weights1[22][439] = 16'b1111111111110101;
    assign weights1[22][440] = 16'b1111111111111110;
    assign weights1[22][441] = 16'b0000000000000110;
    assign weights1[22][442] = 16'b0000000000000100;
    assign weights1[22][443] = 16'b0000000000000001;
    assign weights1[22][444] = 16'b0000000000000011;
    assign weights1[22][445] = 16'b1111111111111100;
    assign weights1[22][446] = 16'b1111111111111011;
    assign weights1[22][447] = 16'b0000000000000101;
    assign weights1[22][448] = 16'b0000000000011000;
    assign weights1[22][449] = 16'b0000000000010010;
    assign weights1[22][450] = 16'b1111111111111111;
    assign weights1[22][451] = 16'b0000000000000010;
    assign weights1[22][452] = 16'b1111111111110100;
    assign weights1[22][453] = 16'b1111111111111000;
    assign weights1[22][454] = 16'b0000000000001010;
    assign weights1[22][455] = 16'b1111111111111000;
    assign weights1[22][456] = 16'b0000000000000011;
    assign weights1[22][457] = 16'b0000000000001000;
    assign weights1[22][458] = 16'b0000000000000111;
    assign weights1[22][459] = 16'b1111111111110111;
    assign weights1[22][460] = 16'b1111111111110011;
    assign weights1[22][461] = 16'b0000000000000111;
    assign weights1[22][462] = 16'b1111111111111010;
    assign weights1[22][463] = 16'b1111111111110110;
    assign weights1[22][464] = 16'b1111111111110011;
    assign weights1[22][465] = 16'b0000000000000010;
    assign weights1[22][466] = 16'b0000000000000000;
    assign weights1[22][467] = 16'b1111111111111000;
    assign weights1[22][468] = 16'b1111111111111101;
    assign weights1[22][469] = 16'b1111111111110110;
    assign weights1[22][470] = 16'b0000000000001011;
    assign weights1[22][471] = 16'b1111111111110001;
    assign weights1[22][472] = 16'b0000000000000101;
    assign weights1[22][473] = 16'b1111111111111110;
    assign weights1[22][474] = 16'b0000000000000101;
    assign weights1[22][475] = 16'b0000000000010101;
    assign weights1[22][476] = 16'b0000000000001111;
    assign weights1[22][477] = 16'b0000000000001110;
    assign weights1[22][478] = 16'b1111111111110001;
    assign weights1[22][479] = 16'b1111111111110110;
    assign weights1[22][480] = 16'b0000000000001000;
    assign weights1[22][481] = 16'b0000000000001110;
    assign weights1[22][482] = 16'b1111111111111011;
    assign weights1[22][483] = 16'b0000000000000000;
    assign weights1[22][484] = 16'b0000000000001010;
    assign weights1[22][485] = 16'b1111111111101000;
    assign weights1[22][486] = 16'b0000000000000010;
    assign weights1[22][487] = 16'b0000000000000001;
    assign weights1[22][488] = 16'b1111111111111101;
    assign weights1[22][489] = 16'b1111111111110101;
    assign weights1[22][490] = 16'b1111111111111010;
    assign weights1[22][491] = 16'b1111111111111110;
    assign weights1[22][492] = 16'b1111111111111111;
    assign weights1[22][493] = 16'b1111111111111011;
    assign weights1[22][494] = 16'b1111111111110100;
    assign weights1[22][495] = 16'b0000000000000001;
    assign weights1[22][496] = 16'b0000000000000010;
    assign weights1[22][497] = 16'b1111111111111010;
    assign weights1[22][498] = 16'b0000000000000101;
    assign weights1[22][499] = 16'b1111111111110111;
    assign weights1[22][500] = 16'b0000000000000100;
    assign weights1[22][501] = 16'b0000000000000101;
    assign weights1[22][502] = 16'b0000000000000111;
    assign weights1[22][503] = 16'b0000000000000011;
    assign weights1[22][504] = 16'b0000000000001101;
    assign weights1[22][505] = 16'b0000000000000011;
    assign weights1[22][506] = 16'b1111111111101010;
    assign weights1[22][507] = 16'b1111111111101101;
    assign weights1[22][508] = 16'b1111111111101110;
    assign weights1[22][509] = 16'b0000000000000000;
    assign weights1[22][510] = 16'b1111111111110100;
    assign weights1[22][511] = 16'b1111111111110111;
    assign weights1[22][512] = 16'b0000000000010011;
    assign weights1[22][513] = 16'b0000000000000110;
    assign weights1[22][514] = 16'b0000000000000010;
    assign weights1[22][515] = 16'b0000000000000111;
    assign weights1[22][516] = 16'b1111111111111100;
    assign weights1[22][517] = 16'b0000000000000000;
    assign weights1[22][518] = 16'b1111111111111110;
    assign weights1[22][519] = 16'b1111111111100110;
    assign weights1[22][520] = 16'b0000000000010010;
    assign weights1[22][521] = 16'b1111111111110101;
    assign weights1[22][522] = 16'b1111111111111000;
    assign weights1[22][523] = 16'b1111111111111011;
    assign weights1[22][524] = 16'b0000000000000110;
    assign weights1[22][525] = 16'b0000000000010100;
    assign weights1[22][526] = 16'b0000000000000110;
    assign weights1[22][527] = 16'b0000000000010100;
    assign weights1[22][528] = 16'b1111111111110000;
    assign weights1[22][529] = 16'b0000000000001010;
    assign weights1[22][530] = 16'b1111111111111101;
    assign weights1[22][531] = 16'b0000000000000111;
    assign weights1[22][532] = 16'b1111111111111001;
    assign weights1[22][533] = 16'b1111111111111000;
    assign weights1[22][534] = 16'b1111111111011010;
    assign weights1[22][535] = 16'b1111111111101101;
    assign weights1[22][536] = 16'b0000000000001110;
    assign weights1[22][537] = 16'b0000000000001111;
    assign weights1[22][538] = 16'b0000000000000010;
    assign weights1[22][539] = 16'b1111111111110100;
    assign weights1[22][540] = 16'b1111111111110110;
    assign weights1[22][541] = 16'b1111111111111011;
    assign weights1[22][542] = 16'b0000000000000010;
    assign weights1[22][543] = 16'b0000000000000001;
    assign weights1[22][544] = 16'b1111111111110100;
    assign weights1[22][545] = 16'b1111111111111010;
    assign weights1[22][546] = 16'b0000000000000100;
    assign weights1[22][547] = 16'b1111111111110100;
    assign weights1[22][548] = 16'b1111111111111010;
    assign weights1[22][549] = 16'b0000000000000010;
    assign weights1[22][550] = 16'b0000000000000110;
    assign weights1[22][551] = 16'b1111111111111101;
    assign weights1[22][552] = 16'b1111111111111001;
    assign weights1[22][553] = 16'b1111111111101101;
    assign weights1[22][554] = 16'b1111111111100101;
    assign weights1[22][555] = 16'b1111111111110100;
    assign weights1[22][556] = 16'b1111111111111101;
    assign weights1[22][557] = 16'b1111111111111001;
    assign weights1[22][558] = 16'b1111111111111110;
    assign weights1[22][559] = 16'b0000000000001000;
    assign weights1[22][560] = 16'b1111111111110101;
    assign weights1[22][561] = 16'b1111111111111111;
    assign weights1[22][562] = 16'b1111111111100110;
    assign weights1[22][563] = 16'b1111111111111110;
    assign weights1[22][564] = 16'b0000000000000101;
    assign weights1[22][565] = 16'b0000000000010100;
    assign weights1[22][566] = 16'b1111111111111001;
    assign weights1[22][567] = 16'b0000000000001000;
    assign weights1[22][568] = 16'b1111111111111111;
    assign weights1[22][569] = 16'b1111111111110101;
    assign weights1[22][570] = 16'b1111111111111111;
    assign weights1[22][571] = 16'b0000000000000000;
    assign weights1[22][572] = 16'b1111111111111000;
    assign weights1[22][573] = 16'b0000000000001010;
    assign weights1[22][574] = 16'b1111111111110111;
    assign weights1[22][575] = 16'b1111111111111111;
    assign weights1[22][576] = 16'b1111111111110001;
    assign weights1[22][577] = 16'b1111111111111110;
    assign weights1[22][578] = 16'b1111111111111001;
    assign weights1[22][579] = 16'b1111111111111101;
    assign weights1[22][580] = 16'b1111111111110111;
    assign weights1[22][581] = 16'b0000000000000101;
    assign weights1[22][582] = 16'b0000000000000111;
    assign weights1[22][583] = 16'b0000000000001000;
    assign weights1[22][584] = 16'b0000000000001000;
    assign weights1[22][585] = 16'b0000000000000011;
    assign weights1[22][586] = 16'b1111111111111100;
    assign weights1[22][587] = 16'b1111111111111011;
    assign weights1[22][588] = 16'b1111111111110100;
    assign weights1[22][589] = 16'b1111111111110100;
    assign weights1[22][590] = 16'b1111111111100101;
    assign weights1[22][591] = 16'b1111111111110111;
    assign weights1[22][592] = 16'b1111111111111010;
    assign weights1[22][593] = 16'b0000000000000001;
    assign weights1[22][594] = 16'b0000000000000000;
    assign weights1[22][595] = 16'b1111111111111000;
    assign weights1[22][596] = 16'b1111111111111110;
    assign weights1[22][597] = 16'b1111111111111100;
    assign weights1[22][598] = 16'b1111111111111001;
    assign weights1[22][599] = 16'b1111111111100010;
    assign weights1[22][600] = 16'b1111111111111111;
    assign weights1[22][601] = 16'b1111111111101011;
    assign weights1[22][602] = 16'b1111111111111110;
    assign weights1[22][603] = 16'b1111111111111101;
    assign weights1[22][604] = 16'b0000000000000111;
    assign weights1[22][605] = 16'b1111111111111000;
    assign weights1[22][606] = 16'b0000000000000100;
    assign weights1[22][607] = 16'b0000000000000100;
    assign weights1[22][608] = 16'b1111111111110111;
    assign weights1[22][609] = 16'b0000000000000010;
    assign weights1[22][610] = 16'b0000000000000100;
    assign weights1[22][611] = 16'b0000000000000101;
    assign weights1[22][612] = 16'b1111111111111010;
    assign weights1[22][613] = 16'b0000000000000000;
    assign weights1[22][614] = 16'b0000000000000000;
    assign weights1[22][615] = 16'b0000000000000100;
    assign weights1[22][616] = 16'b1111111111110110;
    assign weights1[22][617] = 16'b1111111111110101;
    assign weights1[22][618] = 16'b1111111111110100;
    assign weights1[22][619] = 16'b1111111111110001;
    assign weights1[22][620] = 16'b1111111111111101;
    assign weights1[22][621] = 16'b0000000000001000;
    assign weights1[22][622] = 16'b1111111111101100;
    assign weights1[22][623] = 16'b1111111111111111;
    assign weights1[22][624] = 16'b1111111111110000;
    assign weights1[22][625] = 16'b1111111111110100;
    assign weights1[22][626] = 16'b0000000000010100;
    assign weights1[22][627] = 16'b0000000000011000;
    assign weights1[22][628] = 16'b1111111111111000;
    assign weights1[22][629] = 16'b0000000000000001;
    assign weights1[22][630] = 16'b1111111111110111;
    assign weights1[22][631] = 16'b0000000000001011;
    assign weights1[22][632] = 16'b1111111111110111;
    assign weights1[22][633] = 16'b1111111111110011;
    assign weights1[22][634] = 16'b1111111111111101;
    assign weights1[22][635] = 16'b1111111111110000;
    assign weights1[22][636] = 16'b1111111111111010;
    assign weights1[22][637] = 16'b1111111111110110;
    assign weights1[22][638] = 16'b1111111111101111;
    assign weights1[22][639] = 16'b0000000000001001;
    assign weights1[22][640] = 16'b1111111111111010;
    assign weights1[22][641] = 16'b1111111111111111;
    assign weights1[22][642] = 16'b1111111111110100;
    assign weights1[22][643] = 16'b1111111111111111;
    assign weights1[22][644] = 16'b1111111111111010;
    assign weights1[22][645] = 16'b1111111111111000;
    assign weights1[22][646] = 16'b1111111111110101;
    assign weights1[22][647] = 16'b1111111111100101;
    assign weights1[22][648] = 16'b1111111111101100;
    assign weights1[22][649] = 16'b1111111111101110;
    assign weights1[22][650] = 16'b1111111111110110;
    assign weights1[22][651] = 16'b1111111111101110;
    assign weights1[22][652] = 16'b1111111111111000;
    assign weights1[22][653] = 16'b1111111111111111;
    assign weights1[22][654] = 16'b1111111111110101;
    assign weights1[22][655] = 16'b1111111111110110;
    assign weights1[22][656] = 16'b1111111111111011;
    assign weights1[22][657] = 16'b1111111111101111;
    assign weights1[22][658] = 16'b1111111111111111;
    assign weights1[22][659] = 16'b1111111111111111;
    assign weights1[22][660] = 16'b1111111111111010;
    assign weights1[22][661] = 16'b1111111111110000;
    assign weights1[22][662] = 16'b1111111111111000;
    assign weights1[22][663] = 16'b0000000000000100;
    assign weights1[22][664] = 16'b0000000000011110;
    assign weights1[22][665] = 16'b0000000000000111;
    assign weights1[22][666] = 16'b0000000000001000;
    assign weights1[22][667] = 16'b1111111111111011;
    assign weights1[22][668] = 16'b0000000000000010;
    assign weights1[22][669] = 16'b1111111111111000;
    assign weights1[22][670] = 16'b1111111111111010;
    assign weights1[22][671] = 16'b0000000000000001;
    assign weights1[22][672] = 16'b1111111111110111;
    assign weights1[22][673] = 16'b1111111111101110;
    assign weights1[22][674] = 16'b1111111111111010;
    assign weights1[22][675] = 16'b1111111111110100;
    assign weights1[22][676] = 16'b1111111111110010;
    assign weights1[22][677] = 16'b1111111111110011;
    assign weights1[22][678] = 16'b1111111111110010;
    assign weights1[22][679] = 16'b1111111111111001;
    assign weights1[22][680] = 16'b0000000000000000;
    assign weights1[22][681] = 16'b0000000000000001;
    assign weights1[22][682] = 16'b1111111111110111;
    assign weights1[22][683] = 16'b1111111111111101;
    assign weights1[22][684] = 16'b1111111111110101;
    assign weights1[22][685] = 16'b0000000000010010;
    assign weights1[22][686] = 16'b1111111111111000;
    assign weights1[22][687] = 16'b1111111111111011;
    assign weights1[22][688] = 16'b1111111111111001;
    assign weights1[22][689] = 16'b0000000000000011;
    assign weights1[22][690] = 16'b0000000000001010;
    assign weights1[22][691] = 16'b1111111111110110;
    assign weights1[22][692] = 16'b1111111111110100;
    assign weights1[22][693] = 16'b0000000000001011;
    assign weights1[22][694] = 16'b1111111111111011;
    assign weights1[22][695] = 16'b0000000000000010;
    assign weights1[22][696] = 16'b1111111111110101;
    assign weights1[22][697] = 16'b0000000000000000;
    assign weights1[22][698] = 16'b1111111111111101;
    assign weights1[22][699] = 16'b0000000000000101;
    assign weights1[22][700] = 16'b1111111111111000;
    assign weights1[22][701] = 16'b1111111111111000;
    assign weights1[22][702] = 16'b1111111111110011;
    assign weights1[22][703] = 16'b1111111111110110;
    assign weights1[22][704] = 16'b0000000000000001;
    assign weights1[22][705] = 16'b1111111111111011;
    assign weights1[22][706] = 16'b1111111111101000;
    assign weights1[22][707] = 16'b1111111111100010;
    assign weights1[22][708] = 16'b1111111111110100;
    assign weights1[22][709] = 16'b1111111111110000;
    assign weights1[22][710] = 16'b1111111111111110;
    assign weights1[22][711] = 16'b1111111111101011;
    assign weights1[22][712] = 16'b1111111111111001;
    assign weights1[22][713] = 16'b1111111111111111;
    assign weights1[22][714] = 16'b1111111111100110;
    assign weights1[22][715] = 16'b0000000000010001;
    assign weights1[22][716] = 16'b1111111111110110;
    assign weights1[22][717] = 16'b0000000000000110;
    assign weights1[22][718] = 16'b0000000000000101;
    assign weights1[22][719] = 16'b0000000000000100;
    assign weights1[22][720] = 16'b0000000000000101;
    assign weights1[22][721] = 16'b1111111111111111;
    assign weights1[22][722] = 16'b1111111111111100;
    assign weights1[22][723] = 16'b1111111111111011;
    assign weights1[22][724] = 16'b1111111111110110;
    assign weights1[22][725] = 16'b0000000000000011;
    assign weights1[22][726] = 16'b0000000000000000;
    assign weights1[22][727] = 16'b0000000000000001;
    assign weights1[22][728] = 16'b1111111111111100;
    assign weights1[22][729] = 16'b1111111111111110;
    assign weights1[22][730] = 16'b1111111111110111;
    assign weights1[22][731] = 16'b0000000000000100;
    assign weights1[22][732] = 16'b1111111111110111;
    assign weights1[22][733] = 16'b1111111111110011;
    assign weights1[22][734] = 16'b1111111111101111;
    assign weights1[22][735] = 16'b1111111111101010;
    assign weights1[22][736] = 16'b1111111111101011;
    assign weights1[22][737] = 16'b1111111111100111;
    assign weights1[22][738] = 16'b1111111111100111;
    assign weights1[22][739] = 16'b1111111111101100;
    assign weights1[22][740] = 16'b1111111111110011;
    assign weights1[22][741] = 16'b1111111111101011;
    assign weights1[22][742] = 16'b0000000000000110;
    assign weights1[22][743] = 16'b1111111111111110;
    assign weights1[22][744] = 16'b1111111111111010;
    assign weights1[22][745] = 16'b0000000000000000;
    assign weights1[22][746] = 16'b1111111111101011;
    assign weights1[22][747] = 16'b1111111111111101;
    assign weights1[22][748] = 16'b0000000000000110;
    assign weights1[22][749] = 16'b0000000000001000;
    assign weights1[22][750] = 16'b1111111111110111;
    assign weights1[22][751] = 16'b0000000000000000;
    assign weights1[22][752] = 16'b0000000000001010;
    assign weights1[22][753] = 16'b0000000000001001;
    assign weights1[22][754] = 16'b0000000000000000;
    assign weights1[22][755] = 16'b0000000000000100;
    assign weights1[22][756] = 16'b1111111111111111;
    assign weights1[22][757] = 16'b1111111111111100;
    assign weights1[22][758] = 16'b1111111111111101;
    assign weights1[22][759] = 16'b1111111111110011;
    assign weights1[22][760] = 16'b0000000000000011;
    assign weights1[22][761] = 16'b1111111111111001;
    assign weights1[22][762] = 16'b1111111111101101;
    assign weights1[22][763] = 16'b1111111111111001;
    assign weights1[22][764] = 16'b0000000000000010;
    assign weights1[22][765] = 16'b0000000000000111;
    assign weights1[22][766] = 16'b1111111111111011;
    assign weights1[22][767] = 16'b0000000000010011;
    assign weights1[22][768] = 16'b0000000000010110;
    assign weights1[22][769] = 16'b0000000000011011;
    assign weights1[22][770] = 16'b0000000000001110;
    assign weights1[22][771] = 16'b0000000000001010;
    assign weights1[22][772] = 16'b0000000000010101;
    assign weights1[22][773] = 16'b0000000000010100;
    assign weights1[22][774] = 16'b0000000000010001;
    assign weights1[22][775] = 16'b0000000000001011;
    assign weights1[22][776] = 16'b0000000000011000;
    assign weights1[22][777] = 16'b0000000000011000;
    assign weights1[22][778] = 16'b0000000000010010;
    assign weights1[22][779] = 16'b0000000000010101;
    assign weights1[22][780] = 16'b0000000000010010;
    assign weights1[22][781] = 16'b0000000000001000;
    assign weights1[22][782] = 16'b0000000000000110;
    assign weights1[22][783] = 16'b0000000000000011;
    assign weights1[23][0] = 16'b0000000000000000;
    assign weights1[23][1] = 16'b1111111111111111;
    assign weights1[23][2] = 16'b1111111111111111;
    assign weights1[23][3] = 16'b0000000000000000;
    assign weights1[23][4] = 16'b0000000000000000;
    assign weights1[23][5] = 16'b0000000000000000;
    assign weights1[23][6] = 16'b0000000000000001;
    assign weights1[23][7] = 16'b0000000000000010;
    assign weights1[23][8] = 16'b1111111111111001;
    assign weights1[23][9] = 16'b1111111111111110;
    assign weights1[23][10] = 16'b0000000000000000;
    assign weights1[23][11] = 16'b1111111111111100;
    assign weights1[23][12] = 16'b1111111111111011;
    assign weights1[23][13] = 16'b1111111111111110;
    assign weights1[23][14] = 16'b0000000000000001;
    assign weights1[23][15] = 16'b1111111111111101;
    assign weights1[23][16] = 16'b1111111111111111;
    assign weights1[23][17] = 16'b0000000000000011;
    assign weights1[23][18] = 16'b1111111111111110;
    assign weights1[23][19] = 16'b1111111111111111;
    assign weights1[23][20] = 16'b1111111111111110;
    assign weights1[23][21] = 16'b1111111111111100;
    assign weights1[23][22] = 16'b1111111111111111;
    assign weights1[23][23] = 16'b1111111111111111;
    assign weights1[23][24] = 16'b0000000000000000;
    assign weights1[23][25] = 16'b1111111111111111;
    assign weights1[23][26] = 16'b0000000000000000;
    assign weights1[23][27] = 16'b0000000000000000;
    assign weights1[23][28] = 16'b1111111111111111;
    assign weights1[23][29] = 16'b1111111111111110;
    assign weights1[23][30] = 16'b1111111111111110;
    assign weights1[23][31] = 16'b1111111111111110;
    assign weights1[23][32] = 16'b1111111111111111;
    assign weights1[23][33] = 16'b1111111111111011;
    assign weights1[23][34] = 16'b0000000000000000;
    assign weights1[23][35] = 16'b0000000000000000;
    assign weights1[23][36] = 16'b1111111111110111;
    assign weights1[23][37] = 16'b1111111111111010;
    assign weights1[23][38] = 16'b1111111111111000;
    assign weights1[23][39] = 16'b1111111111111101;
    assign weights1[23][40] = 16'b1111111111111101;
    assign weights1[23][41] = 16'b1111111111111010;
    assign weights1[23][42] = 16'b0000000000000001;
    assign weights1[23][43] = 16'b1111111111111110;
    assign weights1[23][44] = 16'b0000000000000100;
    assign weights1[23][45] = 16'b0000000000000011;
    assign weights1[23][46] = 16'b1111111111110111;
    assign weights1[23][47] = 16'b1111111111111000;
    assign weights1[23][48] = 16'b1111111111110111;
    assign weights1[23][49] = 16'b1111111111111010;
    assign weights1[23][50] = 16'b1111111111111110;
    assign weights1[23][51] = 16'b1111111111111111;
    assign weights1[23][52] = 16'b0000000000000000;
    assign weights1[23][53] = 16'b1111111111111101;
    assign weights1[23][54] = 16'b0000000000000000;
    assign weights1[23][55] = 16'b0000000000000000;
    assign weights1[23][56] = 16'b1111111111111111;
    assign weights1[23][57] = 16'b1111111111111111;
    assign weights1[23][58] = 16'b1111111111111111;
    assign weights1[23][59] = 16'b1111111111111100;
    assign weights1[23][60] = 16'b1111111111111101;
    assign weights1[23][61] = 16'b1111111111111100;
    assign weights1[23][62] = 16'b1111111111111011;
    assign weights1[23][63] = 16'b0000000000000000;
    assign weights1[23][64] = 16'b1111111111110000;
    assign weights1[23][65] = 16'b1111111111110010;
    assign weights1[23][66] = 16'b1111111111101111;
    assign weights1[23][67] = 16'b1111111111110101;
    assign weights1[23][68] = 16'b1111111111111001;
    assign weights1[23][69] = 16'b0000000000000011;
    assign weights1[23][70] = 16'b1111111111111000;
    assign weights1[23][71] = 16'b0000000000000100;
    assign weights1[23][72] = 16'b0000000000001000;
    assign weights1[23][73] = 16'b0000000000000010;
    assign weights1[23][74] = 16'b0000000000000111;
    assign weights1[23][75] = 16'b1111111111110011;
    assign weights1[23][76] = 16'b1111111111101010;
    assign weights1[23][77] = 16'b1111111111110111;
    assign weights1[23][78] = 16'b1111111111111110;
    assign weights1[23][79] = 16'b1111111111111100;
    assign weights1[23][80] = 16'b0000000000000000;
    assign weights1[23][81] = 16'b0000000000000100;
    assign weights1[23][82] = 16'b0000000000000000;
    assign weights1[23][83] = 16'b0000000000000000;
    assign weights1[23][84] = 16'b1111111111111111;
    assign weights1[23][85] = 16'b1111111111111111;
    assign weights1[23][86] = 16'b1111111111111110;
    assign weights1[23][87] = 16'b1111111111111100;
    assign weights1[23][88] = 16'b1111111111111001;
    assign weights1[23][89] = 16'b1111111111111000;
    assign weights1[23][90] = 16'b1111111111110011;
    assign weights1[23][91] = 16'b1111111111101000;
    assign weights1[23][92] = 16'b1111111111101100;
    assign weights1[23][93] = 16'b1111111111101010;
    assign weights1[23][94] = 16'b1111111111111010;
    assign weights1[23][95] = 16'b1111111111110101;
    assign weights1[23][96] = 16'b1111111111100010;
    assign weights1[23][97] = 16'b1111111111011110;
    assign weights1[23][98] = 16'b1111111111110111;
    assign weights1[23][99] = 16'b1111111111110100;
    assign weights1[23][100] = 16'b1111111111100101;
    assign weights1[23][101] = 16'b1111111111101010;
    assign weights1[23][102] = 16'b1111111111110001;
    assign weights1[23][103] = 16'b1111111111111000;
    assign weights1[23][104] = 16'b1111111111110100;
    assign weights1[23][105] = 16'b1111111111111011;
    assign weights1[23][106] = 16'b1111111111111100;
    assign weights1[23][107] = 16'b1111111111101111;
    assign weights1[23][108] = 16'b0000000000000111;
    assign weights1[23][109] = 16'b1111111111111010;
    assign weights1[23][110] = 16'b1111111111111100;
    assign weights1[23][111] = 16'b0000000000000010;
    assign weights1[23][112] = 16'b1111111111111110;
    assign weights1[23][113] = 16'b1111111111111101;
    assign weights1[23][114] = 16'b0000000000000000;
    assign weights1[23][115] = 16'b1111111111111011;
    assign weights1[23][116] = 16'b1111111111111010;
    assign weights1[23][117] = 16'b1111111111111011;
    assign weights1[23][118] = 16'b1111111111111100;
    assign weights1[23][119] = 16'b0000000000001001;
    assign weights1[23][120] = 16'b0000000000000000;
    assign weights1[23][121] = 16'b1111111111101000;
    assign weights1[23][122] = 16'b1111111111101001;
    assign weights1[23][123] = 16'b1111111111101011;
    assign weights1[23][124] = 16'b1111111111101101;
    assign weights1[23][125] = 16'b1111111111111010;
    assign weights1[23][126] = 16'b1111111111111011;
    assign weights1[23][127] = 16'b0000000000001110;
    assign weights1[23][128] = 16'b0000000000001100;
    assign weights1[23][129] = 16'b0000000000010101;
    assign weights1[23][130] = 16'b0000000000000111;
    assign weights1[23][131] = 16'b0000000000010011;
    assign weights1[23][132] = 16'b1111111111111000;
    assign weights1[23][133] = 16'b1111111111110101;
    assign weights1[23][134] = 16'b1111111111111110;
    assign weights1[23][135] = 16'b1111111111101010;
    assign weights1[23][136] = 16'b1111111111111001;
    assign weights1[23][137] = 16'b1111111111111110;
    assign weights1[23][138] = 16'b0000000000000010;
    assign weights1[23][139] = 16'b0000000000000001;
    assign weights1[23][140] = 16'b1111111111111110;
    assign weights1[23][141] = 16'b1111111111111001;
    assign weights1[23][142] = 16'b1111111111111011;
    assign weights1[23][143] = 16'b1111111111110011;
    assign weights1[23][144] = 16'b1111111111110010;
    assign weights1[23][145] = 16'b1111111111110011;
    assign weights1[23][146] = 16'b1111111111111000;
    assign weights1[23][147] = 16'b0000000000000010;
    assign weights1[23][148] = 16'b1111111111111000;
    assign weights1[23][149] = 16'b1111111111101010;
    assign weights1[23][150] = 16'b0000000000000110;
    assign weights1[23][151] = 16'b1111111111110101;
    assign weights1[23][152] = 16'b1111111111110010;
    assign weights1[23][153] = 16'b0000000000000000;
    assign weights1[23][154] = 16'b1111111111101111;
    assign weights1[23][155] = 16'b0000000000001111;
    assign weights1[23][156] = 16'b0000000000010000;
    assign weights1[23][157] = 16'b0000000000000101;
    assign weights1[23][158] = 16'b1111111111110101;
    assign weights1[23][159] = 16'b0000000000001010;
    assign weights1[23][160] = 16'b1111111111111111;
    assign weights1[23][161] = 16'b1111111111111100;
    assign weights1[23][162] = 16'b1111111111111011;
    assign weights1[23][163] = 16'b1111111111110110;
    assign weights1[23][164] = 16'b1111111111110101;
    assign weights1[23][165] = 16'b1111111111111011;
    assign weights1[23][166] = 16'b1111111111111111;
    assign weights1[23][167] = 16'b1111111111111101;
    assign weights1[23][168] = 16'b1111111111111100;
    assign weights1[23][169] = 16'b1111111111110111;
    assign weights1[23][170] = 16'b1111111111110010;
    assign weights1[23][171] = 16'b1111111111110110;
    assign weights1[23][172] = 16'b1111111111101011;
    assign weights1[23][173] = 16'b1111111111110100;
    assign weights1[23][174] = 16'b1111111111111011;
    assign weights1[23][175] = 16'b1111111111111111;
    assign weights1[23][176] = 16'b0000000000001011;
    assign weights1[23][177] = 16'b1111111111111100;
    assign weights1[23][178] = 16'b1111111111101101;
    assign weights1[23][179] = 16'b1111111111101011;
    assign weights1[23][180] = 16'b0000000000000011;
    assign weights1[23][181] = 16'b1111111111111011;
    assign weights1[23][182] = 16'b0000000000000001;
    assign weights1[23][183] = 16'b1111111111110001;
    assign weights1[23][184] = 16'b1111111111110001;
    assign weights1[23][185] = 16'b1111111111110000;
    assign weights1[23][186] = 16'b0000000000001010;
    assign weights1[23][187] = 16'b0000000000010111;
    assign weights1[23][188] = 16'b0000000000000110;
    assign weights1[23][189] = 16'b0000000000000110;
    assign weights1[23][190] = 16'b0000000000000001;
    assign weights1[23][191] = 16'b0000000000000101;
    assign weights1[23][192] = 16'b1111111111111010;
    assign weights1[23][193] = 16'b0000000000001100;
    assign weights1[23][194] = 16'b1111111111111100;
    assign weights1[23][195] = 16'b0000000000001011;
    assign weights1[23][196] = 16'b1111111111111000;
    assign weights1[23][197] = 16'b1111111111111000;
    assign weights1[23][198] = 16'b1111111111111010;
    assign weights1[23][199] = 16'b0000000000000111;
    assign weights1[23][200] = 16'b1111111111110111;
    assign weights1[23][201] = 16'b0000000000000111;
    assign weights1[23][202] = 16'b0000000000000111;
    assign weights1[23][203] = 16'b0000000000000110;
    assign weights1[23][204] = 16'b0000000000000110;
    assign weights1[23][205] = 16'b1111111111010100;
    assign weights1[23][206] = 16'b1111111111111011;
    assign weights1[23][207] = 16'b1111111111110011;
    assign weights1[23][208] = 16'b0000000000000000;
    assign weights1[23][209] = 16'b1111111111110110;
    assign weights1[23][210] = 16'b1111111111111110;
    assign weights1[23][211] = 16'b0000000000000100;
    assign weights1[23][212] = 16'b1111111111111101;
    assign weights1[23][213] = 16'b1111111111111011;
    assign weights1[23][214] = 16'b0000000000001000;
    assign weights1[23][215] = 16'b1111111111111010;
    assign weights1[23][216] = 16'b1111111111110111;
    assign weights1[23][217] = 16'b0000000000010000;
    assign weights1[23][218] = 16'b0000000000010000;
    assign weights1[23][219] = 16'b0000000000001110;
    assign weights1[23][220] = 16'b0000000000000110;
    assign weights1[23][221] = 16'b1111111111111101;
    assign weights1[23][222] = 16'b0000000000001100;
    assign weights1[23][223] = 16'b0000000000001000;
    assign weights1[23][224] = 16'b1111111111111100;
    assign weights1[23][225] = 16'b1111111111111011;
    assign weights1[23][226] = 16'b1111111111111001;
    assign weights1[23][227] = 16'b1111111111110100;
    assign weights1[23][228] = 16'b1111111111111100;
    assign weights1[23][229] = 16'b1111111111110000;
    assign weights1[23][230] = 16'b1111111111111001;
    assign weights1[23][231] = 16'b0000000000011011;
    assign weights1[23][232] = 16'b1111111111111100;
    assign weights1[23][233] = 16'b1111111111111100;
    assign weights1[23][234] = 16'b1111111111111000;
    assign weights1[23][235] = 16'b1111111111111000;
    assign weights1[23][236] = 16'b0000000000001001;
    assign weights1[23][237] = 16'b0000000000001100;
    assign weights1[23][238] = 16'b1111111111111100;
    assign weights1[23][239] = 16'b0000000000001000;
    assign weights1[23][240] = 16'b1111111111111111;
    assign weights1[23][241] = 16'b1111111111111001;
    assign weights1[23][242] = 16'b0000000000000000;
    assign weights1[23][243] = 16'b0000000000001101;
    assign weights1[23][244] = 16'b0000000000000000;
    assign weights1[23][245] = 16'b1111111111111110;
    assign weights1[23][246] = 16'b0000000000001100;
    assign weights1[23][247] = 16'b0000000000000110;
    assign weights1[23][248] = 16'b1111111111111111;
    assign weights1[23][249] = 16'b1111111111110011;
    assign weights1[23][250] = 16'b0000000000010100;
    assign weights1[23][251] = 16'b0000000000000101;
    assign weights1[23][252] = 16'b1111111111111101;
    assign weights1[23][253] = 16'b1111111111110111;
    assign weights1[23][254] = 16'b1111111111110111;
    assign weights1[23][255] = 16'b1111111111101101;
    assign weights1[23][256] = 16'b1111111111110111;
    assign weights1[23][257] = 16'b1111111111110110;
    assign weights1[23][258] = 16'b0000000000000110;
    assign weights1[23][259] = 16'b0000000000010001;
    assign weights1[23][260] = 16'b0000000000010011;
    assign weights1[23][261] = 16'b0000000000010000;
    assign weights1[23][262] = 16'b1111111111100111;
    assign weights1[23][263] = 16'b1111111111101000;
    assign weights1[23][264] = 16'b1111111111101000;
    assign weights1[23][265] = 16'b1111111111111101;
    assign weights1[23][266] = 16'b1111111111111010;
    assign weights1[23][267] = 16'b0000000000000111;
    assign weights1[23][268] = 16'b0000000000000010;
    assign weights1[23][269] = 16'b0000000000000110;
    assign weights1[23][270] = 16'b1111111111110100;
    assign weights1[23][271] = 16'b1111111111110110;
    assign weights1[23][272] = 16'b0000000000000110;
    assign weights1[23][273] = 16'b0000000000001011;
    assign weights1[23][274] = 16'b1111111111111101;
    assign weights1[23][275] = 16'b0000000000011011;
    assign weights1[23][276] = 16'b0000000000000011;
    assign weights1[23][277] = 16'b0000000000010011;
    assign weights1[23][278] = 16'b0000000000001010;
    assign weights1[23][279] = 16'b0000000000000011;
    assign weights1[23][280] = 16'b1111111111111000;
    assign weights1[23][281] = 16'b0000000000000100;
    assign weights1[23][282] = 16'b0000000000000111;
    assign weights1[23][283] = 16'b1111111111110010;
    assign weights1[23][284] = 16'b1111111111110011;
    assign weights1[23][285] = 16'b0000000000000011;
    assign weights1[23][286] = 16'b1111111111111101;
    assign weights1[23][287] = 16'b1111111111111111;
    assign weights1[23][288] = 16'b0000000000010110;
    assign weights1[23][289] = 16'b0000000000000011;
    assign weights1[23][290] = 16'b0000000000010111;
    assign weights1[23][291] = 16'b0000000000000100;
    assign weights1[23][292] = 16'b1111111111110000;
    assign weights1[23][293] = 16'b1111111111111100;
    assign weights1[23][294] = 16'b1111111111110101;
    assign weights1[23][295] = 16'b1111111111111001;
    assign weights1[23][296] = 16'b1111111111110111;
    assign weights1[23][297] = 16'b0000000000000111;
    assign weights1[23][298] = 16'b1111111111110100;
    assign weights1[23][299] = 16'b1111111111111101;
    assign weights1[23][300] = 16'b0000000000010100;
    assign weights1[23][301] = 16'b1111111111111101;
    assign weights1[23][302] = 16'b1111111111101011;
    assign weights1[23][303] = 16'b0000000000001010;
    assign weights1[23][304] = 16'b0000000000010011;
    assign weights1[23][305] = 16'b1111111111100101;
    assign weights1[23][306] = 16'b0000000000000111;
    assign weights1[23][307] = 16'b1111111111111111;
    assign weights1[23][308] = 16'b1111111111111111;
    assign weights1[23][309] = 16'b0000000000000111;
    assign weights1[23][310] = 16'b0000000000000101;
    assign weights1[23][311] = 16'b0000000000000000;
    assign weights1[23][312] = 16'b1111111111111110;
    assign weights1[23][313] = 16'b1111111111111000;
    assign weights1[23][314] = 16'b0000000000001011;
    assign weights1[23][315] = 16'b0000000000000100;
    assign weights1[23][316] = 16'b1111111111111001;
    assign weights1[23][317] = 16'b1111111111111100;
    assign weights1[23][318] = 16'b1111111111110111;
    assign weights1[23][319] = 16'b0000000000001010;
    assign weights1[23][320] = 16'b0000000000000101;
    assign weights1[23][321] = 16'b1111111111101100;
    assign weights1[23][322] = 16'b1111111111111110;
    assign weights1[23][323] = 16'b1111111111101100;
    assign weights1[23][324] = 16'b1111111111110100;
    assign weights1[23][325] = 16'b1111111111111001;
    assign weights1[23][326] = 16'b0000000000001000;
    assign weights1[23][327] = 16'b0000000000000100;
    assign weights1[23][328] = 16'b1111111111111101;
    assign weights1[23][329] = 16'b1111111111101110;
    assign weights1[23][330] = 16'b0000000000010011;
    assign weights1[23][331] = 16'b0000000000010001;
    assign weights1[23][332] = 16'b1111111111111100;
    assign weights1[23][333] = 16'b1111111111111101;
    assign weights1[23][334] = 16'b0000000000001110;
    assign weights1[23][335] = 16'b0000000000001011;
    assign weights1[23][336] = 16'b0000000000000110;
    assign weights1[23][337] = 16'b0000000000000111;
    assign weights1[23][338] = 16'b0000000000000110;
    assign weights1[23][339] = 16'b0000000000001110;
    assign weights1[23][340] = 16'b0000000000010110;
    assign weights1[23][341] = 16'b0000000000010101;
    assign weights1[23][342] = 16'b1111111111111111;
    assign weights1[23][343] = 16'b0000000000011110;
    assign weights1[23][344] = 16'b0000000000001001;
    assign weights1[23][345] = 16'b1111111111110000;
    assign weights1[23][346] = 16'b1111111111110000;
    assign weights1[23][347] = 16'b0000000000000101;
    assign weights1[23][348] = 16'b1111111111100010;
    assign weights1[23][349] = 16'b1111111111100101;
    assign weights1[23][350] = 16'b1111111111011011;
    assign weights1[23][351] = 16'b1111111111101101;
    assign weights1[23][352] = 16'b1111111111100001;
    assign weights1[23][353] = 16'b1111111111110101;
    assign weights1[23][354] = 16'b1111111111110011;
    assign weights1[23][355] = 16'b1111111111101000;
    assign weights1[23][356] = 16'b0000000000001000;
    assign weights1[23][357] = 16'b1111111111110101;
    assign weights1[23][358] = 16'b1111111111111001;
    assign weights1[23][359] = 16'b1111111111110011;
    assign weights1[23][360] = 16'b0000000000000000;
    assign weights1[23][361] = 16'b0000000000001000;
    assign weights1[23][362] = 16'b0000000000001100;
    assign weights1[23][363] = 16'b1111111111111100;
    assign weights1[23][364] = 16'b1111111111111010;
    assign weights1[23][365] = 16'b1111111111111011;
    assign weights1[23][366] = 16'b1111111111111110;
    assign weights1[23][367] = 16'b0000000000000110;
    assign weights1[23][368] = 16'b0000000000010101;
    assign weights1[23][369] = 16'b1111111111111011;
    assign weights1[23][370] = 16'b1111111111101010;
    assign weights1[23][371] = 16'b1111111111101111;
    assign weights1[23][372] = 16'b0000000000000001;
    assign weights1[23][373] = 16'b0000000000001001;
    assign weights1[23][374] = 16'b1111111111110111;
    assign weights1[23][375] = 16'b1111111111101000;
    assign weights1[23][376] = 16'b1111111111100011;
    assign weights1[23][377] = 16'b1111111111100011;
    assign weights1[23][378] = 16'b1111111111101001;
    assign weights1[23][379] = 16'b1111111111100110;
    assign weights1[23][380] = 16'b1111111111011110;
    assign weights1[23][381] = 16'b1111111111110010;
    assign weights1[23][382] = 16'b0000000000000110;
    assign weights1[23][383] = 16'b0000000000001001;
    assign weights1[23][384] = 16'b0000000000001101;
    assign weights1[23][385] = 16'b0000000000001010;
    assign weights1[23][386] = 16'b0000000000010100;
    assign weights1[23][387] = 16'b1111111111110110;
    assign weights1[23][388] = 16'b0000000000010100;
    assign weights1[23][389] = 16'b0000000000010110;
    assign weights1[23][390] = 16'b1111111111111000;
    assign weights1[23][391] = 16'b1111111111011110;
    assign weights1[23][392] = 16'b1111111111110100;
    assign weights1[23][393] = 16'b1111111111101110;
    assign weights1[23][394] = 16'b1111111111110101;
    assign weights1[23][395] = 16'b1111111111111010;
    assign weights1[23][396] = 16'b0000000000000001;
    assign weights1[23][397] = 16'b1111111111110001;
    assign weights1[23][398] = 16'b0000000000001001;
    assign weights1[23][399] = 16'b1111111111100111;
    assign weights1[23][400] = 16'b1111111111110010;
    assign weights1[23][401] = 16'b1111111111101000;
    assign weights1[23][402] = 16'b1111111111011011;
    assign weights1[23][403] = 16'b1111111111010001;
    assign weights1[23][404] = 16'b1111111111001001;
    assign weights1[23][405] = 16'b0000000000000000;
    assign weights1[23][406] = 16'b1111111111110100;
    assign weights1[23][407] = 16'b1111111111110100;
    assign weights1[23][408] = 16'b1111111111110100;
    assign weights1[23][409] = 16'b1111111111110100;
    assign weights1[23][410] = 16'b1111111111010101;
    assign weights1[23][411] = 16'b1111111111101111;
    assign weights1[23][412] = 16'b0000000000000001;
    assign weights1[23][413] = 16'b0000000000100101;
    assign weights1[23][414] = 16'b0000000000010001;
    assign weights1[23][415] = 16'b0000000000011110;
    assign weights1[23][416] = 16'b0000000000101000;
    assign weights1[23][417] = 16'b0000000000010001;
    assign weights1[23][418] = 16'b1111111111101100;
    assign weights1[23][419] = 16'b1111111111010101;
    assign weights1[23][420] = 16'b1111111111110111;
    assign weights1[23][421] = 16'b1111111111101110;
    assign weights1[23][422] = 16'b1111111111100100;
    assign weights1[23][423] = 16'b1111111111011111;
    assign weights1[23][424] = 16'b1111111111100000;
    assign weights1[23][425] = 16'b1111111111100010;
    assign weights1[23][426] = 16'b1111111111101110;
    assign weights1[23][427] = 16'b1111111111101101;
    assign weights1[23][428] = 16'b1111111111010011;
    assign weights1[23][429] = 16'b1111111110110001;
    assign weights1[23][430] = 16'b1111111111001100;
    assign weights1[23][431] = 16'b1111111111010101;
    assign weights1[23][432] = 16'b1111111111111101;
    assign weights1[23][433] = 16'b1111111111111111;
    assign weights1[23][434] = 16'b0000000000000110;
    assign weights1[23][435] = 16'b1111111111111110;
    assign weights1[23][436] = 16'b1111111111100001;
    assign weights1[23][437] = 16'b1111111111101101;
    assign weights1[23][438] = 16'b0000000000000110;
    assign weights1[23][439] = 16'b1111111111101001;
    assign weights1[23][440] = 16'b1111111111111011;
    assign weights1[23][441] = 16'b0000000000010000;
    assign weights1[23][442] = 16'b0000000000101011;
    assign weights1[23][443] = 16'b0000000000101010;
    assign weights1[23][444] = 16'b0000000000001101;
    assign weights1[23][445] = 16'b1111111111000101;
    assign weights1[23][446] = 16'b1111111110110010;
    assign weights1[23][447] = 16'b1111111110110101;
    assign weights1[23][448] = 16'b1111111111101111;
    assign weights1[23][449] = 16'b1111111111101100;
    assign weights1[23][450] = 16'b1111111111010001;
    assign weights1[23][451] = 16'b1111111110111101;
    assign weights1[23][452] = 16'b1111111111010011;
    assign weights1[23][453] = 16'b1111111111010000;
    assign weights1[23][454] = 16'b1111111110111011;
    assign weights1[23][455] = 16'b1111111110111010;
    assign weights1[23][456] = 16'b1111111110011101;
    assign weights1[23][457] = 16'b1111111111001101;
    assign weights1[23][458] = 16'b1111111111010001;
    assign weights1[23][459] = 16'b1111111111111111;
    assign weights1[23][460] = 16'b0000000000010000;
    assign weights1[23][461] = 16'b0000000000010010;
    assign weights1[23][462] = 16'b0000000000010001;
    assign weights1[23][463] = 16'b0000000000010010;
    assign weights1[23][464] = 16'b1111111111110110;
    assign weights1[23][465] = 16'b1111111111101111;
    assign weights1[23][466] = 16'b1111111111110001;
    assign weights1[23][467] = 16'b1111111111110000;
    assign weights1[23][468] = 16'b1111111111111011;
    assign weights1[23][469] = 16'b0000000000001000;
    assign weights1[23][470] = 16'b1111111111111000;
    assign weights1[23][471] = 16'b1111111111001101;
    assign weights1[23][472] = 16'b1111111110110100;
    assign weights1[23][473] = 16'b1111111110010110;
    assign weights1[23][474] = 16'b1111111110101011;
    assign weights1[23][475] = 16'b1111111110110011;
    assign weights1[23][476] = 16'b1111111111101100;
    assign weights1[23][477] = 16'b1111111111011110;
    assign weights1[23][478] = 16'b1111111111001000;
    assign weights1[23][479] = 16'b1111111110110000;
    assign weights1[23][480] = 16'b1111111110111000;
    assign weights1[23][481] = 16'b1111111110100011;
    assign weights1[23][482] = 16'b1111111110010110;
    assign weights1[23][483] = 16'b1111111110011011;
    assign weights1[23][484] = 16'b1111111111010011;
    assign weights1[23][485] = 16'b1111111111110111;
    assign weights1[23][486] = 16'b0000000000000100;
    assign weights1[23][487] = 16'b0000000000011001;
    assign weights1[23][488] = 16'b0000000000011000;
    assign weights1[23][489] = 16'b0000000000010111;
    assign weights1[23][490] = 16'b0000000000000010;
    assign weights1[23][491] = 16'b0000000000011000;
    assign weights1[23][492] = 16'b0000000000000110;
    assign weights1[23][493] = 16'b1111111111110101;
    assign weights1[23][494] = 16'b1111111111011111;
    assign weights1[23][495] = 16'b1111111111010101;
    assign weights1[23][496] = 16'b1111111110110000;
    assign weights1[23][497] = 16'b1111111110101010;
    assign weights1[23][498] = 16'b1111111101111100;
    assign weights1[23][499] = 16'b1111111101101101;
    assign weights1[23][500] = 16'b1111111101111011;
    assign weights1[23][501] = 16'b1111111110100100;
    assign weights1[23][502] = 16'b1111111110100011;
    assign weights1[23][503] = 16'b1111111110110110;
    assign weights1[23][504] = 16'b1111111111101011;
    assign weights1[23][505] = 16'b1111111111011001;
    assign weights1[23][506] = 16'b1111111111001011;
    assign weights1[23][507] = 16'b1111111110111000;
    assign weights1[23][508] = 16'b1111111110110010;
    assign weights1[23][509] = 16'b1111111110100101;
    assign weights1[23][510] = 16'b1111111111010000;
    assign weights1[23][511] = 16'b1111111111100100;
    assign weights1[23][512] = 16'b1111111111111110;
    assign weights1[23][513] = 16'b0000000000011001;
    assign weights1[23][514] = 16'b0000000000011110;
    assign weights1[23][515] = 16'b0000000000100010;
    assign weights1[23][516] = 16'b0000000000000101;
    assign weights1[23][517] = 16'b0000000000010100;
    assign weights1[23][518] = 16'b0000000000000000;
    assign weights1[23][519] = 16'b0000000000001001;
    assign weights1[23][520] = 16'b1111111111111101;
    assign weights1[23][521] = 16'b1111111111100001;
    assign weights1[23][522] = 16'b1111111111010111;
    assign weights1[23][523] = 16'b1111111110110111;
    assign weights1[23][524] = 16'b1111111101111011;
    assign weights1[23][525] = 16'b1111111100111010;
    assign weights1[23][526] = 16'b1111111100101101;
    assign weights1[23][527] = 16'b1111111101011110;
    assign weights1[23][528] = 16'b1111111101110110;
    assign weights1[23][529] = 16'b1111111110100010;
    assign weights1[23][530] = 16'b1111111110100110;
    assign weights1[23][531] = 16'b1111111110110001;
    assign weights1[23][532] = 16'b1111111111101011;
    assign weights1[23][533] = 16'b1111111111100000;
    assign weights1[23][534] = 16'b1111111111010001;
    assign weights1[23][535] = 16'b1111111111010010;
    assign weights1[23][536] = 16'b1111111111001011;
    assign weights1[23][537] = 16'b1111111111011111;
    assign weights1[23][538] = 16'b1111111111100101;
    assign weights1[23][539] = 16'b0000000000010000;
    assign weights1[23][540] = 16'b0000000000011011;
    assign weights1[23][541] = 16'b0000000000011111;
    assign weights1[23][542] = 16'b1111111111111101;
    assign weights1[23][543] = 16'b0000000000010111;
    assign weights1[23][544] = 16'b0000000000010110;
    assign weights1[23][545] = 16'b0000000000010011;
    assign weights1[23][546] = 16'b0000000000010111;
    assign weights1[23][547] = 16'b1111111111111110;
    assign weights1[23][548] = 16'b0000000000000110;
    assign weights1[23][549] = 16'b1111111111111110;
    assign weights1[23][550] = 16'b1111111111011010;
    assign weights1[23][551] = 16'b1111111111000100;
    assign weights1[23][552] = 16'b1111111110000111;
    assign weights1[23][553] = 16'b1111111101101010;
    assign weights1[23][554] = 16'b1111111101101001;
    assign weights1[23][555] = 16'b1111111101111110;
    assign weights1[23][556] = 16'b1111111110000100;
    assign weights1[23][557] = 16'b1111111110011111;
    assign weights1[23][558] = 16'b1111111110100101;
    assign weights1[23][559] = 16'b1111111111000000;
    assign weights1[23][560] = 16'b1111111111101101;
    assign weights1[23][561] = 16'b1111111111100100;
    assign weights1[23][562] = 16'b1111111111011100;
    assign weights1[23][563] = 16'b1111111111100010;
    assign weights1[23][564] = 16'b1111111111111011;
    assign weights1[23][565] = 16'b0000000000000010;
    assign weights1[23][566] = 16'b0000000000100100;
    assign weights1[23][567] = 16'b0000000000100101;
    assign weights1[23][568] = 16'b0000000000001111;
    assign weights1[23][569] = 16'b0000000000011110;
    assign weights1[23][570] = 16'b0000000000100001;
    assign weights1[23][571] = 16'b0000000000001001;
    assign weights1[23][572] = 16'b0000000000000111;
    assign weights1[23][573] = 16'b0000000000010100;
    assign weights1[23][574] = 16'b0000000000010111;
    assign weights1[23][575] = 16'b0000000000010000;
    assign weights1[23][576] = 16'b0000000000000001;
    assign weights1[23][577] = 16'b0000000000010000;
    assign weights1[23][578] = 16'b1111111111110010;
    assign weights1[23][579] = 16'b1111111111011001;
    assign weights1[23][580] = 16'b0000000000000010;
    assign weights1[23][581] = 16'b1111111111011111;
    assign weights1[23][582] = 16'b1111111111001111;
    assign weights1[23][583] = 16'b1111111110101100;
    assign weights1[23][584] = 16'b1111111110110000;
    assign weights1[23][585] = 16'b1111111110110110;
    assign weights1[23][586] = 16'b1111111110111010;
    assign weights1[23][587] = 16'b1111111111001100;
    assign weights1[23][588] = 16'b1111111111110100;
    assign weights1[23][589] = 16'b1111111111110011;
    assign weights1[23][590] = 16'b1111111111111110;
    assign weights1[23][591] = 16'b0000000000000111;
    assign weights1[23][592] = 16'b0000000000001010;
    assign weights1[23][593] = 16'b0000000000011111;
    assign weights1[23][594] = 16'b0000000000101100;
    assign weights1[23][595] = 16'b0000000000000111;
    assign weights1[23][596] = 16'b0000000000010000;
    assign weights1[23][597] = 16'b0000000000001001;
    assign weights1[23][598] = 16'b0000000000011111;
    assign weights1[23][599] = 16'b0000000000100001;
    assign weights1[23][600] = 16'b0000000000101101;
    assign weights1[23][601] = 16'b0000000000100110;
    assign weights1[23][602] = 16'b0000000000001010;
    assign weights1[23][603] = 16'b0000000000111000;
    assign weights1[23][604] = 16'b0000000000100000;
    assign weights1[23][605] = 16'b0000000000100011;
    assign weights1[23][606] = 16'b0000000000111110;
    assign weights1[23][607] = 16'b0000000000101001;
    assign weights1[23][608] = 16'b0000000000101100;
    assign weights1[23][609] = 16'b0000000000101101;
    assign weights1[23][610] = 16'b0000000000100011;
    assign weights1[23][611] = 16'b0000000000001000;
    assign weights1[23][612] = 16'b1111111111011100;
    assign weights1[23][613] = 16'b1111111111010111;
    assign weights1[23][614] = 16'b1111111111011000;
    assign weights1[23][615] = 16'b1111111111100001;
    assign weights1[23][616] = 16'b0000000000000111;
    assign weights1[23][617] = 16'b0000000000001110;
    assign weights1[23][618] = 16'b0000000000001111;
    assign weights1[23][619] = 16'b0000000000010100;
    assign weights1[23][620] = 16'b0000000000010000;
    assign weights1[23][621] = 16'b0000000000100010;
    assign weights1[23][622] = 16'b0000000000001001;
    assign weights1[23][623] = 16'b0000000000000001;
    assign weights1[23][624] = 16'b0000000000011001;
    assign weights1[23][625] = 16'b0000000000010101;
    assign weights1[23][626] = 16'b0000000000011110;
    assign weights1[23][627] = 16'b0000000000011000;
    assign weights1[23][628] = 16'b0000000000101010;
    assign weights1[23][629] = 16'b0000000000110001;
    assign weights1[23][630] = 16'b0000000000100000;
    assign weights1[23][631] = 16'b0000000000101110;
    assign weights1[23][632] = 16'b0000000000100111;
    assign weights1[23][633] = 16'b0000000000101110;
    assign weights1[23][634] = 16'b0000000001001101;
    assign weights1[23][635] = 16'b0000000000110111;
    assign weights1[23][636] = 16'b0000000000111011;
    assign weights1[23][637] = 16'b0000000001010111;
    assign weights1[23][638] = 16'b0000000001000101;
    assign weights1[23][639] = 16'b0000000000100001;
    assign weights1[23][640] = 16'b0000000000010011;
    assign weights1[23][641] = 16'b1111111111110011;
    assign weights1[23][642] = 16'b1111111111111001;
    assign weights1[23][643] = 16'b1111111111110011;
    assign weights1[23][644] = 16'b0000000000001011;
    assign weights1[23][645] = 16'b0000000000011011;
    assign weights1[23][646] = 16'b0000000000011001;
    assign weights1[23][647] = 16'b0000000000010011;
    assign weights1[23][648] = 16'b0000000000100101;
    assign weights1[23][649] = 16'b0000000000010010;
    assign weights1[23][650] = 16'b0000000000000100;
    assign weights1[23][651] = 16'b0000000000001010;
    assign weights1[23][652] = 16'b0000000000011111;
    assign weights1[23][653] = 16'b0000000000001100;
    assign weights1[23][654] = 16'b0000000000011110;
    assign weights1[23][655] = 16'b0000000000010001;
    assign weights1[23][656] = 16'b0000000000011110;
    assign weights1[23][657] = 16'b0000000000100011;
    assign weights1[23][658] = 16'b0000000000011011;
    assign weights1[23][659] = 16'b0000000000100110;
    assign weights1[23][660] = 16'b0000000001000110;
    assign weights1[23][661] = 16'b0000000000010100;
    assign weights1[23][662] = 16'b0000000000100001;
    assign weights1[23][663] = 16'b0000000001001000;
    assign weights1[23][664] = 16'b0000000000111110;
    assign weights1[23][665] = 16'b0000000000101111;
    assign weights1[23][666] = 16'b0000000001010100;
    assign weights1[23][667] = 16'b0000000001000000;
    assign weights1[23][668] = 16'b0000000000101111;
    assign weights1[23][669] = 16'b0000000000011001;
    assign weights1[23][670] = 16'b0000000000001111;
    assign weights1[23][671] = 16'b0000000000001011;
    assign weights1[23][672] = 16'b0000000000000001;
    assign weights1[23][673] = 16'b0000000000000111;
    assign weights1[23][674] = 16'b0000000000000001;
    assign weights1[23][675] = 16'b0000000000000100;
    assign weights1[23][676] = 16'b0000000000001010;
    assign weights1[23][677] = 16'b0000000000010011;
    assign weights1[23][678] = 16'b1111111111111110;
    assign weights1[23][679] = 16'b1111111111111000;
    assign weights1[23][680] = 16'b0000000000001000;
    assign weights1[23][681] = 16'b0000000000010111;
    assign weights1[23][682] = 16'b0000000000000101;
    assign weights1[23][683] = 16'b0000000000011110;
    assign weights1[23][684] = 16'b0000000000100000;
    assign weights1[23][685] = 16'b0000000000010100;
    assign weights1[23][686] = 16'b0000000000010101;
    assign weights1[23][687] = 16'b0000000000011110;
    assign weights1[23][688] = 16'b0000000000000111;
    assign weights1[23][689] = 16'b0000000000110011;
    assign weights1[23][690] = 16'b0000000000101101;
    assign weights1[23][691] = 16'b0000000000100011;
    assign weights1[23][692] = 16'b0000000000100110;
    assign weights1[23][693] = 16'b0000000000101011;
    assign weights1[23][694] = 16'b0000000001011111;
    assign weights1[23][695] = 16'b0000000000110111;
    assign weights1[23][696] = 16'b0000000000101011;
    assign weights1[23][697] = 16'b0000000000101000;
    assign weights1[23][698] = 16'b0000000000011110;
    assign weights1[23][699] = 16'b0000000000001100;
    assign weights1[23][700] = 16'b0000000000000001;
    assign weights1[23][701] = 16'b0000000000000100;
    assign weights1[23][702] = 16'b0000000000000000;
    assign weights1[23][703] = 16'b0000000000001001;
    assign weights1[23][704] = 16'b0000000000010100;
    assign weights1[23][705] = 16'b0000000000011111;
    assign weights1[23][706] = 16'b0000000000010100;
    assign weights1[23][707] = 16'b0000000000010011;
    assign weights1[23][708] = 16'b0000000000001010;
    assign weights1[23][709] = 16'b0000000000001101;
    assign weights1[23][710] = 16'b0000000000001011;
    assign weights1[23][711] = 16'b1111111111110100;
    assign weights1[23][712] = 16'b0000000000001011;
    assign weights1[23][713] = 16'b0000000000010111;
    assign weights1[23][714] = 16'b0000000000001010;
    assign weights1[23][715] = 16'b0000000000011000;
    assign weights1[23][716] = 16'b0000000000001000;
    assign weights1[23][717] = 16'b0000000000011000;
    assign weights1[23][718] = 16'b0000000000010110;
    assign weights1[23][719] = 16'b0000000000100011;
    assign weights1[23][720] = 16'b0000000000110010;
    assign weights1[23][721] = 16'b0000000000001101;
    assign weights1[23][722] = 16'b0000000000101111;
    assign weights1[23][723] = 16'b0000000000110111;
    assign weights1[23][724] = 16'b0000000000110010;
    assign weights1[23][725] = 16'b0000000000100100;
    assign weights1[23][726] = 16'b0000000000011001;
    assign weights1[23][727] = 16'b0000000000000111;
    assign weights1[23][728] = 16'b0000000000000000;
    assign weights1[23][729] = 16'b1111111111111111;
    assign weights1[23][730] = 16'b0000000000000110;
    assign weights1[23][731] = 16'b0000000000001110;
    assign weights1[23][732] = 16'b0000000000000000;
    assign weights1[23][733] = 16'b0000000000000100;
    assign weights1[23][734] = 16'b0000000000011011;
    assign weights1[23][735] = 16'b0000000000011001;
    assign weights1[23][736] = 16'b0000000000010100;
    assign weights1[23][737] = 16'b0000000000010100;
    assign weights1[23][738] = 16'b0000000000000010;
    assign weights1[23][739] = 16'b0000000000010000;
    assign weights1[23][740] = 16'b0000000000001011;
    assign weights1[23][741] = 16'b0000000000000101;
    assign weights1[23][742] = 16'b0000000000001111;
    assign weights1[23][743] = 16'b0000000000000111;
    assign weights1[23][744] = 16'b0000000000010110;
    assign weights1[23][745] = 16'b0000000000000010;
    assign weights1[23][746] = 16'b0000000000001111;
    assign weights1[23][747] = 16'b0000000000001111;
    assign weights1[23][748] = 16'b0000000000001110;
    assign weights1[23][749] = 16'b0000000000011010;
    assign weights1[23][750] = 16'b0000000000111110;
    assign weights1[23][751] = 16'b0000000000110001;
    assign weights1[23][752] = 16'b0000000000101010;
    assign weights1[23][753] = 16'b0000000000010010;
    assign weights1[23][754] = 16'b0000000000001011;
    assign weights1[23][755] = 16'b0000000000000100;
    assign weights1[23][756] = 16'b0000000000000010;
    assign weights1[23][757] = 16'b1111111111111111;
    assign weights1[23][758] = 16'b1111111111111111;
    assign weights1[23][759] = 16'b0000000000000001;
    assign weights1[23][760] = 16'b1111111111111001;
    assign weights1[23][761] = 16'b0000000000001010;
    assign weights1[23][762] = 16'b0000000000010000;
    assign weights1[23][763] = 16'b1111111111111101;
    assign weights1[23][764] = 16'b0000000000001111;
    assign weights1[23][765] = 16'b0000000000001011;
    assign weights1[23][766] = 16'b1111111111111011;
    assign weights1[23][767] = 16'b0000000000000110;
    assign weights1[23][768] = 16'b1111111111111110;
    assign weights1[23][769] = 16'b1111111111111111;
    assign weights1[23][770] = 16'b1111111111111011;
    assign weights1[23][771] = 16'b0000000000010011;
    assign weights1[23][772] = 16'b0000000000010000;
    assign weights1[23][773] = 16'b0000000000010110;
    assign weights1[23][774] = 16'b0000000000000110;
    assign weights1[23][775] = 16'b1111111111111100;
    assign weights1[23][776] = 16'b0000000000010001;
    assign weights1[23][777] = 16'b0000000000101001;
    assign weights1[23][778] = 16'b0000000000100110;
    assign weights1[23][779] = 16'b0000000000011101;
    assign weights1[23][780] = 16'b0000000000010111;
    assign weights1[23][781] = 16'b0000000000001000;
    assign weights1[23][782] = 16'b0000000000000100;
    assign weights1[23][783] = 16'b0000000000000100;
    assign weights1[24][0] = 16'b0000000000000000;
    assign weights1[24][1] = 16'b0000000000000000;
    assign weights1[24][2] = 16'b0000000000000001;
    assign weights1[24][3] = 16'b0000000000000010;
    assign weights1[24][4] = 16'b0000000000000111;
    assign weights1[24][5] = 16'b0000000000000101;
    assign weights1[24][6] = 16'b0000000000000101;
    assign weights1[24][7] = 16'b1111111111110000;
    assign weights1[24][8] = 16'b1111111111011100;
    assign weights1[24][9] = 16'b1111111111001001;
    assign weights1[24][10] = 16'b1111111110110111;
    assign weights1[24][11] = 16'b1111111110111010;
    assign weights1[24][12] = 16'b1111111111001111;
    assign weights1[24][13] = 16'b1111111111110011;
    assign weights1[24][14] = 16'b0000000000011001;
    assign weights1[24][15] = 16'b0000000000100011;
    assign weights1[24][16] = 16'b0000000000100101;
    assign weights1[24][17] = 16'b0000000000011110;
    assign weights1[24][18] = 16'b1111111111111110;
    assign weights1[24][19] = 16'b1111111111011011;
    assign weights1[24][20] = 16'b1111111111001000;
    assign weights1[24][21] = 16'b1111111111000011;
    assign weights1[24][22] = 16'b1111111111001100;
    assign weights1[24][23] = 16'b1111111111011011;
    assign weights1[24][24] = 16'b1111111111110111;
    assign weights1[24][25] = 16'b0000000000000011;
    assign weights1[24][26] = 16'b0000000000000010;
    assign weights1[24][27] = 16'b1111111111111111;
    assign weights1[24][28] = 16'b0000000000000000;
    assign weights1[24][29] = 16'b0000000000000000;
    assign weights1[24][30] = 16'b0000000000000011;
    assign weights1[24][31] = 16'b0000000000000111;
    assign weights1[24][32] = 16'b0000000000001000;
    assign weights1[24][33] = 16'b0000000000000101;
    assign weights1[24][34] = 16'b1111111111111101;
    assign weights1[24][35] = 16'b1111111111101101;
    assign weights1[24][36] = 16'b1111111111010010;
    assign weights1[24][37] = 16'b1111111110110011;
    assign weights1[24][38] = 16'b1111111110100000;
    assign weights1[24][39] = 16'b1111111110101011;
    assign weights1[24][40] = 16'b1111111111011000;
    assign weights1[24][41] = 16'b0000000000000100;
    assign weights1[24][42] = 16'b0000000000100100;
    assign weights1[24][43] = 16'b0000000000101110;
    assign weights1[24][44] = 16'b0000000000011100;
    assign weights1[24][45] = 16'b0000000000000111;
    assign weights1[24][46] = 16'b1111111111011111;
    assign weights1[24][47] = 16'b1111111110101110;
    assign weights1[24][48] = 16'b1111111110010111;
    assign weights1[24][49] = 16'b1111111110101100;
    assign weights1[24][50] = 16'b1111111111000011;
    assign weights1[24][51] = 16'b1111111111010110;
    assign weights1[24][52] = 16'b1111111111110101;
    assign weights1[24][53] = 16'b0000000000000010;
    assign weights1[24][54] = 16'b0000000000000111;
    assign weights1[24][55] = 16'b0000000000000011;
    assign weights1[24][56] = 16'b0000000000000000;
    assign weights1[24][57] = 16'b0000000000000001;
    assign weights1[24][58] = 16'b0000000000000000;
    assign weights1[24][59] = 16'b0000000000001010;
    assign weights1[24][60] = 16'b0000000000001001;
    assign weights1[24][61] = 16'b0000000000001110;
    assign weights1[24][62] = 16'b0000000000000001;
    assign weights1[24][63] = 16'b1111111111110010;
    assign weights1[24][64] = 16'b1111111110111011;
    assign weights1[24][65] = 16'b1111111110011110;
    assign weights1[24][66] = 16'b1111111110000101;
    assign weights1[24][67] = 16'b1111111110010101;
    assign weights1[24][68] = 16'b1111111111100111;
    assign weights1[24][69] = 16'b0000000000101110;
    assign weights1[24][70] = 16'b0000000000101111;
    assign weights1[24][71] = 16'b0000000000101100;
    assign weights1[24][72] = 16'b0000000000101010;
    assign weights1[24][73] = 16'b0000000000010100;
    assign weights1[24][74] = 16'b1111111111010000;
    assign weights1[24][75] = 16'b1111111110001011;
    assign weights1[24][76] = 16'b1111111101110111;
    assign weights1[24][77] = 16'b1111111110011000;
    assign weights1[24][78] = 16'b1111111111001011;
    assign weights1[24][79] = 16'b1111111111100110;
    assign weights1[24][80] = 16'b1111111111110101;
    assign weights1[24][81] = 16'b0000000000000010;
    assign weights1[24][82] = 16'b0000000000000011;
    assign weights1[24][83] = 16'b0000000000000100;
    assign weights1[24][84] = 16'b0000000000000000;
    assign weights1[24][85] = 16'b0000000000000001;
    assign weights1[24][86] = 16'b0000000000010000;
    assign weights1[24][87] = 16'b0000000000010110;
    assign weights1[24][88] = 16'b0000000000011110;
    assign weights1[24][89] = 16'b0000000000011111;
    assign weights1[24][90] = 16'b0000000000010100;
    assign weights1[24][91] = 16'b1111111111111011;
    assign weights1[24][92] = 16'b1111111110111001;
    assign weights1[24][93] = 16'b1111111110011000;
    assign weights1[24][94] = 16'b1111111110000011;
    assign weights1[24][95] = 16'b1111111110010110;
    assign weights1[24][96] = 16'b1111111111011111;
    assign weights1[24][97] = 16'b0000000000101000;
    assign weights1[24][98] = 16'b0000000000111111;
    assign weights1[24][99] = 16'b0000000000101111;
    assign weights1[24][100] = 16'b0000000000001110;
    assign weights1[24][101] = 16'b0000000000100000;
    assign weights1[24][102] = 16'b1111111110111010;
    assign weights1[24][103] = 16'b1111111101100001;
    assign weights1[24][104] = 16'b1111111101100111;
    assign weights1[24][105] = 16'b1111111110011111;
    assign weights1[24][106] = 16'b1111111111001000;
    assign weights1[24][107] = 16'b1111111111101001;
    assign weights1[24][108] = 16'b0000000000000111;
    assign weights1[24][109] = 16'b0000000000010111;
    assign weights1[24][110] = 16'b0000000000010101;
    assign weights1[24][111] = 16'b0000000000001000;
    assign weights1[24][112] = 16'b0000000000000000;
    assign weights1[24][113] = 16'b0000000000001000;
    assign weights1[24][114] = 16'b0000000000010101;
    assign weights1[24][115] = 16'b0000000000011110;
    assign weights1[24][116] = 16'b0000000000100110;
    assign weights1[24][117] = 16'b0000000000100001;
    assign weights1[24][118] = 16'b0000000000010100;
    assign weights1[24][119] = 16'b1111111111111111;
    assign weights1[24][120] = 16'b1111111110111010;
    assign weights1[24][121] = 16'b1111111101111111;
    assign weights1[24][122] = 16'b1111111101010101;
    assign weights1[24][123] = 16'b1111111110100110;
    assign weights1[24][124] = 16'b1111111111011110;
    assign weights1[24][125] = 16'b0000000001001011;
    assign weights1[24][126] = 16'b0000000000101110;
    assign weights1[24][127] = 16'b0000000000100001;
    assign weights1[24][128] = 16'b0000000000110101;
    assign weights1[24][129] = 16'b1111111111011110;
    assign weights1[24][130] = 16'b1111111110011001;
    assign weights1[24][131] = 16'b1111111101000111;
    assign weights1[24][132] = 16'b1111111101010111;
    assign weights1[24][133] = 16'b1111111110110100;
    assign weights1[24][134] = 16'b1111111111111100;
    assign weights1[24][135] = 16'b0000000000001011;
    assign weights1[24][136] = 16'b0000000000100001;
    assign weights1[24][137] = 16'b0000000000101100;
    assign weights1[24][138] = 16'b0000000000100000;
    assign weights1[24][139] = 16'b0000000000010010;
    assign weights1[24][140] = 16'b0000000000000010;
    assign weights1[24][141] = 16'b0000000000000110;
    assign weights1[24][142] = 16'b0000000000001010;
    assign weights1[24][143] = 16'b0000000000011010;
    assign weights1[24][144] = 16'b0000000000100011;
    assign weights1[24][145] = 16'b0000000000100101;
    assign weights1[24][146] = 16'b0000000000011101;
    assign weights1[24][147] = 16'b0000000000001110;
    assign weights1[24][148] = 16'b1111111111010001;
    assign weights1[24][149] = 16'b1111111110011011;
    assign weights1[24][150] = 16'b1111111101100001;
    assign weights1[24][151] = 16'b1111111111000101;
    assign weights1[24][152] = 16'b0000000000010010;
    assign weights1[24][153] = 16'b0000000000101000;
    assign weights1[24][154] = 16'b0000000000111000;
    assign weights1[24][155] = 16'b0000000000111001;
    assign weights1[24][156] = 16'b0000000000000010;
    assign weights1[24][157] = 16'b1111111111000100;
    assign weights1[24][158] = 16'b1111111101100100;
    assign weights1[24][159] = 16'b1111111101001100;
    assign weights1[24][160] = 16'b1111111101111101;
    assign weights1[24][161] = 16'b1111111111111011;
    assign weights1[24][162] = 16'b0000000000011011;
    assign weights1[24][163] = 16'b0000000000010011;
    assign weights1[24][164] = 16'b0000000000011000;
    assign weights1[24][165] = 16'b0000000000101100;
    assign weights1[24][166] = 16'b0000000000010101;
    assign weights1[24][167] = 16'b0000000000010110;
    assign weights1[24][168] = 16'b1111111111111100;
    assign weights1[24][169] = 16'b0000000000000011;
    assign weights1[24][170] = 16'b0000000000000011;
    assign weights1[24][171] = 16'b0000000000000010;
    assign weights1[24][172] = 16'b0000000000010101;
    assign weights1[24][173] = 16'b0000000000101100;
    assign weights1[24][174] = 16'b0000000000101101;
    assign weights1[24][175] = 16'b0000000000100101;
    assign weights1[24][176] = 16'b1111111111011001;
    assign weights1[24][177] = 16'b1111111101111010;
    assign weights1[24][178] = 16'b1111111101110100;
    assign weights1[24][179] = 16'b1111111111110110;
    assign weights1[24][180] = 16'b0000000000001001;
    assign weights1[24][181] = 16'b0000000000100010;
    assign weights1[24][182] = 16'b0000000000100001;
    assign weights1[24][183] = 16'b0000000000100100;
    assign weights1[24][184] = 16'b0000000000001001;
    assign weights1[24][185] = 16'b1111111110111111;
    assign weights1[24][186] = 16'b1111111101010001;
    assign weights1[24][187] = 16'b1111111101010010;
    assign weights1[24][188] = 16'b1111111111011001;
    assign weights1[24][189] = 16'b0000000000110101;
    assign weights1[24][190] = 16'b0000000000101100;
    assign weights1[24][191] = 16'b0000000000110111;
    assign weights1[24][192] = 16'b0000000000011011;
    assign weights1[24][193] = 16'b0000000000011010;
    assign weights1[24][194] = 16'b0000000000011011;
    assign weights1[24][195] = 16'b0000000000011101;
    assign weights1[24][196] = 16'b0000000000000011;
    assign weights1[24][197] = 16'b1111111111111111;
    assign weights1[24][198] = 16'b0000000000000100;
    assign weights1[24][199] = 16'b0000000000001001;
    assign weights1[24][200] = 16'b1111111111111101;
    assign weights1[24][201] = 16'b0000000000011100;
    assign weights1[24][202] = 16'b0000000000100110;
    assign weights1[24][203] = 16'b0000000000110110;
    assign weights1[24][204] = 16'b1111111111001001;
    assign weights1[24][205] = 16'b1111111110011101;
    assign weights1[24][206] = 16'b1111111110110011;
    assign weights1[24][207] = 16'b1111111111101101;
    assign weights1[24][208] = 16'b0000000000000110;
    assign weights1[24][209] = 16'b0000000000100010;
    assign weights1[24][210] = 16'b0000000000110000;
    assign weights1[24][211] = 16'b0000000000011001;
    assign weights1[24][212] = 16'b1111111111110001;
    assign weights1[24][213] = 16'b1111111110100000;
    assign weights1[24][214] = 16'b1111111101010011;
    assign weights1[24][215] = 16'b1111111110100011;
    assign weights1[24][216] = 16'b0000000000000001;
    assign weights1[24][217] = 16'b0000000000101101;
    assign weights1[24][218] = 16'b0000000000100000;
    assign weights1[24][219] = 16'b0000000000101000;
    assign weights1[24][220] = 16'b0000000000011000;
    assign weights1[24][221] = 16'b0000000000000000;
    assign weights1[24][222] = 16'b0000000000001110;
    assign weights1[24][223] = 16'b0000000000001000;
    assign weights1[24][224] = 16'b0000000000000001;
    assign weights1[24][225] = 16'b1111111111111000;
    assign weights1[24][226] = 16'b1111111111111001;
    assign weights1[24][227] = 16'b1111111111111100;
    assign weights1[24][228] = 16'b0000000000001111;
    assign weights1[24][229] = 16'b0000000000011001;
    assign weights1[24][230] = 16'b0000000000011011;
    assign weights1[24][231] = 16'b0000000000100100;
    assign weights1[24][232] = 16'b1111111111011010;
    assign weights1[24][233] = 16'b1111111111000001;
    assign weights1[24][234] = 16'b1111111111001101;
    assign weights1[24][235] = 16'b1111111111001111;
    assign weights1[24][236] = 16'b0000000000010101;
    assign weights1[24][237] = 16'b0000000000100001;
    assign weights1[24][238] = 16'b0000000000101010;
    assign weights1[24][239] = 16'b0000000000010010;
    assign weights1[24][240] = 16'b1111111111111101;
    assign weights1[24][241] = 16'b1111111110001101;
    assign weights1[24][242] = 16'b1111111100111100;
    assign weights1[24][243] = 16'b1111111111110011;
    assign weights1[24][244] = 16'b0000000000111111;
    assign weights1[24][245] = 16'b0000000000010001;
    assign weights1[24][246] = 16'b0000000000011111;
    assign weights1[24][247] = 16'b0000000000000101;
    assign weights1[24][248] = 16'b0000000000001100;
    assign weights1[24][249] = 16'b0000000000011001;
    assign weights1[24][250] = 16'b0000000000001101;
    assign weights1[24][251] = 16'b0000000000001000;
    assign weights1[24][252] = 16'b1111111111111011;
    assign weights1[24][253] = 16'b1111111111111010;
    assign weights1[24][254] = 16'b0000000000000110;
    assign weights1[24][255] = 16'b1111111111111000;
    assign weights1[24][256] = 16'b1111111111101111;
    assign weights1[24][257] = 16'b0000000000011111;
    assign weights1[24][258] = 16'b0000000000110100;
    assign weights1[24][259] = 16'b0000000000100100;
    assign weights1[24][260] = 16'b1111111111101000;
    assign weights1[24][261] = 16'b1111111111001011;
    assign weights1[24][262] = 16'b1111111111000101;
    assign weights1[24][263] = 16'b0000000000000000;
    assign weights1[24][264] = 16'b0000000000000011;
    assign weights1[24][265] = 16'b0000000000011000;
    assign weights1[24][266] = 16'b0000000000100000;
    assign weights1[24][267] = 16'b0000000000010000;
    assign weights1[24][268] = 16'b1111111111110011;
    assign weights1[24][269] = 16'b1111111110000010;
    assign weights1[24][270] = 16'b1111111110110110;
    assign weights1[24][271] = 16'b0000000000011000;
    assign weights1[24][272] = 16'b0000000000011110;
    assign weights1[24][273] = 16'b0000000000100111;
    assign weights1[24][274] = 16'b0000000000000001;
    assign weights1[24][275] = 16'b0000000000010101;
    assign weights1[24][276] = 16'b0000000000001100;
    assign weights1[24][277] = 16'b0000000000100100;
    assign weights1[24][278] = 16'b0000000000001111;
    assign weights1[24][279] = 16'b0000000000010000;
    assign weights1[24][280] = 16'b1111111111111100;
    assign weights1[24][281] = 16'b0000000000000001;
    assign weights1[24][282] = 16'b1111111111110101;
    assign weights1[24][283] = 16'b0000000000000011;
    assign weights1[24][284] = 16'b1111111111101000;
    assign weights1[24][285] = 16'b0000000000000010;
    assign weights1[24][286] = 16'b0000000000001110;
    assign weights1[24][287] = 16'b0000000000011101;
    assign weights1[24][288] = 16'b0000000000001001;
    assign weights1[24][289] = 16'b1111111111011100;
    assign weights1[24][290] = 16'b1111111111011111;
    assign weights1[24][291] = 16'b1111111111101000;
    assign weights1[24][292] = 16'b1111111111111110;
    assign weights1[24][293] = 16'b0000000000010011;
    assign weights1[24][294] = 16'b0000000000001101;
    assign weights1[24][295] = 16'b0000000000010011;
    assign weights1[24][296] = 16'b1111111111100010;
    assign weights1[24][297] = 16'b1111111110100010;
    assign weights1[24][298] = 16'b1111111111010101;
    assign weights1[24][299] = 16'b0000000000001110;
    assign weights1[24][300] = 16'b0000000000100110;
    assign weights1[24][301] = 16'b0000000000001001;
    assign weights1[24][302] = 16'b0000000000011100;
    assign weights1[24][303] = 16'b0000000000000010;
    assign weights1[24][304] = 16'b0000000000000111;
    assign weights1[24][305] = 16'b0000000000011100;
    assign weights1[24][306] = 16'b0000000000010100;
    assign weights1[24][307] = 16'b1111111111110110;
    assign weights1[24][308] = 16'b1111111111111111;
    assign weights1[24][309] = 16'b0000000000000100;
    assign weights1[24][310] = 16'b1111111111111100;
    assign weights1[24][311] = 16'b0000000000000100;
    assign weights1[24][312] = 16'b1111111111111110;
    assign weights1[24][313] = 16'b1111111111111110;
    assign weights1[24][314] = 16'b0000000000001100;
    assign weights1[24][315] = 16'b0000000000001101;
    assign weights1[24][316] = 16'b1111111111111000;
    assign weights1[24][317] = 16'b1111111111101010;
    assign weights1[24][318] = 16'b1111111111100100;
    assign weights1[24][319] = 16'b1111111111110110;
    assign weights1[24][320] = 16'b1111111111111110;
    assign weights1[24][321] = 16'b1111111111111010;
    assign weights1[24][322] = 16'b0000000000001011;
    assign weights1[24][323] = 16'b0000000000000011;
    assign weights1[24][324] = 16'b1111111111011000;
    assign weights1[24][325] = 16'b1111111111011100;
    assign weights1[24][326] = 16'b1111111111100101;
    assign weights1[24][327] = 16'b0000000000100101;
    assign weights1[24][328] = 16'b0000000000001011;
    assign weights1[24][329] = 16'b0000000000010110;
    assign weights1[24][330] = 16'b0000000000001000;
    assign weights1[24][331] = 16'b0000000000001001;
    assign weights1[24][332] = 16'b0000000000000010;
    assign weights1[24][333] = 16'b0000000000011010;
    assign weights1[24][334] = 16'b0000000000000000;
    assign weights1[24][335] = 16'b1111111111110110;
    assign weights1[24][336] = 16'b1111111111111011;
    assign weights1[24][337] = 16'b1111111111111101;
    assign weights1[24][338] = 16'b0000000000001111;
    assign weights1[24][339] = 16'b0000000000001000;
    assign weights1[24][340] = 16'b0000000000000111;
    assign weights1[24][341] = 16'b1111111111101111;
    assign weights1[24][342] = 16'b1111111111110100;
    assign weights1[24][343] = 16'b0000000000000010;
    assign weights1[24][344] = 16'b0000000000010110;
    assign weights1[24][345] = 16'b1111111111110000;
    assign weights1[24][346] = 16'b0000000000001100;
    assign weights1[24][347] = 16'b1111111111110010;
    assign weights1[24][348] = 16'b1111111111111101;
    assign weights1[24][349] = 16'b1111111111111111;
    assign weights1[24][350] = 16'b0000000000001001;
    assign weights1[24][351] = 16'b1111111111111111;
    assign weights1[24][352] = 16'b1111111111001111;
    assign weights1[24][353] = 16'b1111111111101001;
    assign weights1[24][354] = 16'b1111111111111010;
    assign weights1[24][355] = 16'b0000000000001000;
    assign weights1[24][356] = 16'b0000000000000100;
    assign weights1[24][357] = 16'b0000000000010000;
    assign weights1[24][358] = 16'b1111111111110011;
    assign weights1[24][359] = 16'b0000000000001001;
    assign weights1[24][360] = 16'b1111111111110000;
    assign weights1[24][361] = 16'b0000000000000100;
    assign weights1[24][362] = 16'b1111111111101001;
    assign weights1[24][363] = 16'b1111111111100110;
    assign weights1[24][364] = 16'b1111111111111100;
    assign weights1[24][365] = 16'b1111111111111111;
    assign weights1[24][366] = 16'b1111111111111110;
    assign weights1[24][367] = 16'b1111111111111111;
    assign weights1[24][368] = 16'b0000000000001001;
    assign weights1[24][369] = 16'b0000000000000011;
    assign weights1[24][370] = 16'b1111111111111101;
    assign weights1[24][371] = 16'b0000000000000011;
    assign weights1[24][372] = 16'b0000000000001000;
    assign weights1[24][373] = 16'b1111111111101010;
    assign weights1[24][374] = 16'b0000000000000010;
    assign weights1[24][375] = 16'b1111111111101110;
    assign weights1[24][376] = 16'b1111111111111111;
    assign weights1[24][377] = 16'b0000000000001000;
    assign weights1[24][378] = 16'b1111111111111001;
    assign weights1[24][379] = 16'b1111111111110010;
    assign weights1[24][380] = 16'b1111111111101011;
    assign weights1[24][381] = 16'b0000000000001001;
    assign weights1[24][382] = 16'b0000000000001001;
    assign weights1[24][383] = 16'b0000000000001101;
    assign weights1[24][384] = 16'b0000000000011011;
    assign weights1[24][385] = 16'b0000000000000100;
    assign weights1[24][386] = 16'b0000000000001101;
    assign weights1[24][387] = 16'b0000000000001010;
    assign weights1[24][388] = 16'b1111111111111001;
    assign weights1[24][389] = 16'b1111111111010000;
    assign weights1[24][390] = 16'b1111111111011100;
    assign weights1[24][391] = 16'b1111111111100100;
    assign weights1[24][392] = 16'b1111111111111010;
    assign weights1[24][393] = 16'b0000000000000011;
    assign weights1[24][394] = 16'b1111111111111110;
    assign weights1[24][395] = 16'b0000000000000100;
    assign weights1[24][396] = 16'b0000000000000011;
    assign weights1[24][397] = 16'b0000000000011011;
    assign weights1[24][398] = 16'b0000000000001101;
    assign weights1[24][399] = 16'b1111111111111010;
    assign weights1[24][400] = 16'b0000000000000111;
    assign weights1[24][401] = 16'b0000000000000110;
    assign weights1[24][402] = 16'b0000000000001101;
    assign weights1[24][403] = 16'b1111111111111000;
    assign weights1[24][404] = 16'b1111111111111101;
    assign weights1[24][405] = 16'b0000000000000010;
    assign weights1[24][406] = 16'b0000000000001000;
    assign weights1[24][407] = 16'b1111111111101100;
    assign weights1[24][408] = 16'b0000000000000011;
    assign weights1[24][409] = 16'b1111111111111110;
    assign weights1[24][410] = 16'b0000000000010000;
    assign weights1[24][411] = 16'b1111111111101110;
    assign weights1[24][412] = 16'b0000000000001010;
    assign weights1[24][413] = 16'b1111111111111101;
    assign weights1[24][414] = 16'b0000000000001110;
    assign weights1[24][415] = 16'b1111111111110010;
    assign weights1[24][416] = 16'b1111111111100110;
    assign weights1[24][417] = 16'b0000000000000010;
    assign weights1[24][418] = 16'b0000000000000000;
    assign weights1[24][419] = 16'b1111111111111010;
    assign weights1[24][420] = 16'b0000000000000010;
    assign weights1[24][421] = 16'b0000000000000011;
    assign weights1[24][422] = 16'b1111111111110111;
    assign weights1[24][423] = 16'b1111111111111101;
    assign weights1[24][424] = 16'b1111111111110011;
    assign weights1[24][425] = 16'b1111111111111010;
    assign weights1[24][426] = 16'b1111111111110110;
    assign weights1[24][427] = 16'b0000000000000111;
    assign weights1[24][428] = 16'b0000000000000110;
    assign weights1[24][429] = 16'b0000000000000001;
    assign weights1[24][430] = 16'b1111111111111110;
    assign weights1[24][431] = 16'b1111111111111101;
    assign weights1[24][432] = 16'b1111111111111110;
    assign weights1[24][433] = 16'b1111111111110111;
    assign weights1[24][434] = 16'b0000000000001110;
    assign weights1[24][435] = 16'b0000000000000111;
    assign weights1[24][436] = 16'b0000000000000101;
    assign weights1[24][437] = 16'b1111111111110111;
    assign weights1[24][438] = 16'b0000000000011000;
    assign weights1[24][439] = 16'b1111111111111100;
    assign weights1[24][440] = 16'b0000000000000101;
    assign weights1[24][441] = 16'b1111111111111000;
    assign weights1[24][442] = 16'b1111111111110000;
    assign weights1[24][443] = 16'b0000000000001101;
    assign weights1[24][444] = 16'b0000000000000000;
    assign weights1[24][445] = 16'b1111111111111110;
    assign weights1[24][446] = 16'b1111111111111101;
    assign weights1[24][447] = 16'b1111111111111010;
    assign weights1[24][448] = 16'b1111111111111010;
    assign weights1[24][449] = 16'b1111111111110110;
    assign weights1[24][450] = 16'b0000000000000001;
    assign weights1[24][451] = 16'b0000000000000100;
    assign weights1[24][452] = 16'b0000000000000000;
    assign weights1[24][453] = 16'b0000000000010001;
    assign weights1[24][454] = 16'b0000000000000111;
    assign weights1[24][455] = 16'b1111111111111001;
    assign weights1[24][456] = 16'b0000000000001101;
    assign weights1[24][457] = 16'b1111111111101111;
    assign weights1[24][458] = 16'b0000000000000100;
    assign weights1[24][459] = 16'b0000000000000010;
    assign weights1[24][460] = 16'b1111111111110110;
    assign weights1[24][461] = 16'b1111111111111100;
    assign weights1[24][462] = 16'b0000000000000010;
    assign weights1[24][463] = 16'b0000000000001011;
    assign weights1[24][464] = 16'b1111111111110010;
    assign weights1[24][465] = 16'b1111111111110111;
    assign weights1[24][466] = 16'b0000000000001010;
    assign weights1[24][467] = 16'b1111111111100110;
    assign weights1[24][468] = 16'b0000000000000000;
    assign weights1[24][469] = 16'b1111111111111010;
    assign weights1[24][470] = 16'b1111111111100110;
    assign weights1[24][471] = 16'b1111111111111001;
    assign weights1[24][472] = 16'b1111111111111010;
    assign weights1[24][473] = 16'b1111111111111011;
    assign weights1[24][474] = 16'b0000000000000011;
    assign weights1[24][475] = 16'b1111111111110111;
    assign weights1[24][476] = 16'b1111111111110110;
    assign weights1[24][477] = 16'b1111111111111100;
    assign weights1[24][478] = 16'b0000000000001111;
    assign weights1[24][479] = 16'b1111111111111100;
    assign weights1[24][480] = 16'b0000000000001110;
    assign weights1[24][481] = 16'b0000000000000011;
    assign weights1[24][482] = 16'b0000000000000110;
    assign weights1[24][483] = 16'b0000000000000100;
    assign weights1[24][484] = 16'b1111111111111110;
    assign weights1[24][485] = 16'b0000000000001010;
    assign weights1[24][486] = 16'b0000000000000111;
    assign weights1[24][487] = 16'b1111111111110101;
    assign weights1[24][488] = 16'b1111111111111000;
    assign weights1[24][489] = 16'b0000000000001110;
    assign weights1[24][490] = 16'b0000000000000101;
    assign weights1[24][491] = 16'b0000000000001111;
    assign weights1[24][492] = 16'b0000000000001111;
    assign weights1[24][493] = 16'b1111111111111010;
    assign weights1[24][494] = 16'b0000000000000101;
    assign weights1[24][495] = 16'b0000000000011100;
    assign weights1[24][496] = 16'b1111111111101111;
    assign weights1[24][497] = 16'b0000000000000001;
    assign weights1[24][498] = 16'b0000000000000110;
    assign weights1[24][499] = 16'b0000000000001011;
    assign weights1[24][500] = 16'b0000000000000001;
    assign weights1[24][501] = 16'b1111111111101110;
    assign weights1[24][502] = 16'b0000000000000111;
    assign weights1[24][503] = 16'b0000000000001101;
    assign weights1[24][504] = 16'b1111111111111001;
    assign weights1[24][505] = 16'b1111111111110001;
    assign weights1[24][506] = 16'b0000000000001100;
    assign weights1[24][507] = 16'b0000000000000101;
    assign weights1[24][508] = 16'b0000000000000111;
    assign weights1[24][509] = 16'b0000000000000111;
    assign weights1[24][510] = 16'b1111111111101110;
    assign weights1[24][511] = 16'b1111111111111010;
    assign weights1[24][512] = 16'b0000000000001011;
    assign weights1[24][513] = 16'b1111111111101111;
    assign weights1[24][514] = 16'b0000000000000000;
    assign weights1[24][515] = 16'b1111111111111100;
    assign weights1[24][516] = 16'b0000000000000111;
    assign weights1[24][517] = 16'b0000000000001000;
    assign weights1[24][518] = 16'b0000000000001011;
    assign weights1[24][519] = 16'b0000000000000001;
    assign weights1[24][520] = 16'b1111111111111110;
    assign weights1[24][521] = 16'b0000000000000000;
    assign weights1[24][522] = 16'b1111111111110111;
    assign weights1[24][523] = 16'b0000000000000111;
    assign weights1[24][524] = 16'b0000000000000100;
    assign weights1[24][525] = 16'b0000000000000110;
    assign weights1[24][526] = 16'b1111111111111010;
    assign weights1[24][527] = 16'b0000000000010011;
    assign weights1[24][528] = 16'b1111111111111010;
    assign weights1[24][529] = 16'b1111111111111100;
    assign weights1[24][530] = 16'b1111111111111110;
    assign weights1[24][531] = 16'b0000000000000001;
    assign weights1[24][532] = 16'b1111111111111110;
    assign weights1[24][533] = 16'b1111111111110111;
    assign weights1[24][534] = 16'b1111111111111111;
    assign weights1[24][535] = 16'b0000000000010011;
    assign weights1[24][536] = 16'b0000000000000101;
    assign weights1[24][537] = 16'b1111111111110110;
    assign weights1[24][538] = 16'b0000000000001011;
    assign weights1[24][539] = 16'b0000000000000111;
    assign weights1[24][540] = 16'b1111111111110110;
    assign weights1[24][541] = 16'b1111111111101111;
    assign weights1[24][542] = 16'b1111111111111101;
    assign weights1[24][543] = 16'b1111111111111100;
    assign weights1[24][544] = 16'b0000000000001011;
    assign weights1[24][545] = 16'b0000000000000000;
    assign weights1[24][546] = 16'b0000000000010100;
    assign weights1[24][547] = 16'b1111111111110100;
    assign weights1[24][548] = 16'b0000000000010011;
    assign weights1[24][549] = 16'b0000000000000011;
    assign weights1[24][550] = 16'b0000000000001100;
    assign weights1[24][551] = 16'b0000000000000110;
    assign weights1[24][552] = 16'b1111111111111010;
    assign weights1[24][553] = 16'b1111111111110101;
    assign weights1[24][554] = 16'b0000000000000001;
    assign weights1[24][555] = 16'b0000000000001010;
    assign weights1[24][556] = 16'b0000000000011001;
    assign weights1[24][557] = 16'b0000000000001000;
    assign weights1[24][558] = 16'b1111111111111111;
    assign weights1[24][559] = 16'b1111111111111001;
    assign weights1[24][560] = 16'b0000000000000000;
    assign weights1[24][561] = 16'b0000000000000010;
    assign weights1[24][562] = 16'b1111111111111000;
    assign weights1[24][563] = 16'b0000000000000110;
    assign weights1[24][564] = 16'b0000000000000011;
    assign weights1[24][565] = 16'b1111111111111100;
    assign weights1[24][566] = 16'b0000000000001111;
    assign weights1[24][567] = 16'b1111111111111010;
    assign weights1[24][568] = 16'b0000000000001101;
    assign weights1[24][569] = 16'b1111111111111001;
    assign weights1[24][570] = 16'b1111111111111101;
    assign weights1[24][571] = 16'b0000000000001010;
    assign weights1[24][572] = 16'b0000000000000011;
    assign weights1[24][573] = 16'b0000000000001001;
    assign weights1[24][574] = 16'b0000000000001011;
    assign weights1[24][575] = 16'b0000000000001001;
    assign weights1[24][576] = 16'b0000000000000011;
    assign weights1[24][577] = 16'b1111111111111011;
    assign weights1[24][578] = 16'b1111111111111111;
    assign weights1[24][579] = 16'b1111111111110100;
    assign weights1[24][580] = 16'b0000000000010110;
    assign weights1[24][581] = 16'b0000000000000100;
    assign weights1[24][582] = 16'b1111111111101010;
    assign weights1[24][583] = 16'b1111111111111100;
    assign weights1[24][584] = 16'b1111111111110110;
    assign weights1[24][585] = 16'b1111111111110011;
    assign weights1[24][586] = 16'b1111111111111011;
    assign weights1[24][587] = 16'b0000000000000001;
    assign weights1[24][588] = 16'b0000000000000000;
    assign weights1[24][589] = 16'b0000000000001011;
    assign weights1[24][590] = 16'b0000000000000110;
    assign weights1[24][591] = 16'b1111111111111100;
    assign weights1[24][592] = 16'b1111111111111111;
    assign weights1[24][593] = 16'b1111111111110010;
    assign weights1[24][594] = 16'b0000000000000000;
    assign weights1[24][595] = 16'b1111111111110000;
    assign weights1[24][596] = 16'b1111111111100011;
    assign weights1[24][597] = 16'b0000000000001111;
    assign weights1[24][598] = 16'b1111111111110100;
    assign weights1[24][599] = 16'b1111111111110011;
    assign weights1[24][600] = 16'b1111111111111110;
    assign weights1[24][601] = 16'b1111111111111000;
    assign weights1[24][602] = 16'b0000000000000011;
    assign weights1[24][603] = 16'b0000000000000000;
    assign weights1[24][604] = 16'b1111111111110110;
    assign weights1[24][605] = 16'b0000000000001001;
    assign weights1[24][606] = 16'b1111111111111111;
    assign weights1[24][607] = 16'b1111111111110010;
    assign weights1[24][608] = 16'b1111111111101111;
    assign weights1[24][609] = 16'b0000000000010001;
    assign weights1[24][610] = 16'b0000000000001000;
    assign weights1[24][611] = 16'b0000000000001010;
    assign weights1[24][612] = 16'b1111111111111011;
    assign weights1[24][613] = 16'b0000000000011100;
    assign weights1[24][614] = 16'b1111111111111000;
    assign weights1[24][615] = 16'b1111111111110111;
    assign weights1[24][616] = 16'b0000000000000100;
    assign weights1[24][617] = 16'b1111111111111101;
    assign weights1[24][618] = 16'b0000000000001110;
    assign weights1[24][619] = 16'b0000000000000000;
    assign weights1[24][620] = 16'b0000000000000110;
    assign weights1[24][621] = 16'b1111111111110111;
    assign weights1[24][622] = 16'b0000000000010000;
    assign weights1[24][623] = 16'b0000000000000000;
    assign weights1[24][624] = 16'b1111111111111111;
    assign weights1[24][625] = 16'b1111111111100101;
    assign weights1[24][626] = 16'b1111111111101001;
    assign weights1[24][627] = 16'b1111111111111001;
    assign weights1[24][628] = 16'b0000000000010010;
    assign weights1[24][629] = 16'b1111111111110011;
    assign weights1[24][630] = 16'b1111111111101111;
    assign weights1[24][631] = 16'b0000000000000101;
    assign weights1[24][632] = 16'b0000000000001100;
    assign weights1[24][633] = 16'b0000000000000001;
    assign weights1[24][634] = 16'b0000000000000100;
    assign weights1[24][635] = 16'b0000000000000101;
    assign weights1[24][636] = 16'b1111111111110011;
    assign weights1[24][637] = 16'b1111111111111011;
    assign weights1[24][638] = 16'b0000000000000101;
    assign weights1[24][639] = 16'b0000000000000000;
    assign weights1[24][640] = 16'b1111111111111000;
    assign weights1[24][641] = 16'b1111111111110100;
    assign weights1[24][642] = 16'b1111111111111010;
    assign weights1[24][643] = 16'b1111111111111010;
    assign weights1[24][644] = 16'b0000000000000101;
    assign weights1[24][645] = 16'b0000000000000010;
    assign weights1[24][646] = 16'b0000000000000110;
    assign weights1[24][647] = 16'b1111111111111101;
    assign weights1[24][648] = 16'b1111111111111110;
    assign weights1[24][649] = 16'b0000000000000011;
    assign weights1[24][650] = 16'b0000000000001010;
    assign weights1[24][651] = 16'b0000000000000101;
    assign weights1[24][652] = 16'b0000000000000011;
    assign weights1[24][653] = 16'b0000000000010111;
    assign weights1[24][654] = 16'b0000000000001000;
    assign weights1[24][655] = 16'b1111111111111001;
    assign weights1[24][656] = 16'b1111111111101000;
    assign weights1[24][657] = 16'b0000000000000101;
    assign weights1[24][658] = 16'b1111111111110001;
    assign weights1[24][659] = 16'b0000000000000011;
    assign weights1[24][660] = 16'b1111111111110001;
    assign weights1[24][661] = 16'b0000000000001001;
    assign weights1[24][662] = 16'b1111111111111000;
    assign weights1[24][663] = 16'b0000000000010101;
    assign weights1[24][664] = 16'b1111111111111111;
    assign weights1[24][665] = 16'b1111111111111000;
    assign weights1[24][666] = 16'b1111111111101011;
    assign weights1[24][667] = 16'b1111111111111100;
    assign weights1[24][668] = 16'b1111111111101111;
    assign weights1[24][669] = 16'b1111111111111001;
    assign weights1[24][670] = 16'b0000000000000001;
    assign weights1[24][671] = 16'b1111111111110101;
    assign weights1[24][672] = 16'b0000000000001000;
    assign weights1[24][673] = 16'b0000000000001001;
    assign weights1[24][674] = 16'b0000000000000100;
    assign weights1[24][675] = 16'b1111111111111001;
    assign weights1[24][676] = 16'b1111111111111000;
    assign weights1[24][677] = 16'b0000000000000000;
    assign weights1[24][678] = 16'b0000000000000001;
    assign weights1[24][679] = 16'b0000000000000000;
    assign weights1[24][680] = 16'b1111111111111001;
    assign weights1[24][681] = 16'b0000000000000100;
    assign weights1[24][682] = 16'b0000000000000010;
    assign weights1[24][683] = 16'b0000000000000000;
    assign weights1[24][684] = 16'b1111111111111000;
    assign weights1[24][685] = 16'b1111111111111111;
    assign weights1[24][686] = 16'b1111111111101011;
    assign weights1[24][687] = 16'b1111111111101001;
    assign weights1[24][688] = 16'b1111111111111000;
    assign weights1[24][689] = 16'b1111111111101101;
    assign weights1[24][690] = 16'b0000000000001101;
    assign weights1[24][691] = 16'b0000000000000110;
    assign weights1[24][692] = 16'b1111111111111000;
    assign weights1[24][693] = 16'b0000000000000100;
    assign weights1[24][694] = 16'b0000000000000100;
    assign weights1[24][695] = 16'b0000000000001011;
    assign weights1[24][696] = 16'b1111111111110100;
    assign weights1[24][697] = 16'b1111111111111110;
    assign weights1[24][698] = 16'b0000000000000000;
    assign weights1[24][699] = 16'b1111111111111100;
    assign weights1[24][700] = 16'b0000000000001001;
    assign weights1[24][701] = 16'b0000000000000010;
    assign weights1[24][702] = 16'b0000000000000100;
    assign weights1[24][703] = 16'b1111111111111111;
    assign weights1[24][704] = 16'b1111111111110101;
    assign weights1[24][705] = 16'b1111111111111101;
    assign weights1[24][706] = 16'b1111111111110110;
    assign weights1[24][707] = 16'b1111111111111001;
    assign weights1[24][708] = 16'b1111111111110010;
    assign weights1[24][709] = 16'b0000000000000000;
    assign weights1[24][710] = 16'b0000000000000011;
    assign weights1[24][711] = 16'b0000000000001000;
    assign weights1[24][712] = 16'b1111111111110110;
    assign weights1[24][713] = 16'b1111111111101110;
    assign weights1[24][714] = 16'b1111111111110000;
    assign weights1[24][715] = 16'b0000000000000000;
    assign weights1[24][716] = 16'b1111111111110101;
    assign weights1[24][717] = 16'b1111111111110001;
    assign weights1[24][718] = 16'b1111111111111101;
    assign weights1[24][719] = 16'b1111111111111001;
    assign weights1[24][720] = 16'b0000000000000010;
    assign weights1[24][721] = 16'b1111111111101000;
    assign weights1[24][722] = 16'b0000000000000001;
    assign weights1[24][723] = 16'b0000000000000110;
    assign weights1[24][724] = 16'b1111111111111110;
    assign weights1[24][725] = 16'b1111111111110101;
    assign weights1[24][726] = 16'b1111111111111000;
    assign weights1[24][727] = 16'b1111111111111100;
    assign weights1[24][728] = 16'b0000000000000000;
    assign weights1[24][729] = 16'b0000000000000010;
    assign weights1[24][730] = 16'b0000000000000001;
    assign weights1[24][731] = 16'b1111111111110011;
    assign weights1[24][732] = 16'b1111111111111101;
    assign weights1[24][733] = 16'b1111111111110101;
    assign weights1[24][734] = 16'b1111111111110111;
    assign weights1[24][735] = 16'b1111111111111110;
    assign weights1[24][736] = 16'b1111111111111000;
    assign weights1[24][737] = 16'b0000000000000001;
    assign weights1[24][738] = 16'b1111111111110011;
    assign weights1[24][739] = 16'b1111111111111010;
    assign weights1[24][740] = 16'b1111111111111110;
    assign weights1[24][741] = 16'b1111111111111000;
    assign weights1[24][742] = 16'b0000000000000110;
    assign weights1[24][743] = 16'b1111111111110111;
    assign weights1[24][744] = 16'b0000000000000000;
    assign weights1[24][745] = 16'b1111111111110111;
    assign weights1[24][746] = 16'b1111111111111010;
    assign weights1[24][747] = 16'b1111111111110111;
    assign weights1[24][748] = 16'b0000000000000001;
    assign weights1[24][749] = 16'b0000000000001110;
    assign weights1[24][750] = 16'b0000000000001001;
    assign weights1[24][751] = 16'b0000000000001100;
    assign weights1[24][752] = 16'b1111111111110011;
    assign weights1[24][753] = 16'b1111111111110110;
    assign weights1[24][754] = 16'b1111111111110110;
    assign weights1[24][755] = 16'b0000000000000011;
    assign weights1[24][756] = 16'b1111111111111101;
    assign weights1[24][757] = 16'b1111111111111111;
    assign weights1[24][758] = 16'b1111111111111110;
    assign weights1[24][759] = 16'b1111111111111010;
    assign weights1[24][760] = 16'b1111111111101110;
    assign weights1[24][761] = 16'b1111111111111110;
    assign weights1[24][762] = 16'b1111111111111101;
    assign weights1[24][763] = 16'b1111111111101110;
    assign weights1[24][764] = 16'b1111111111111011;
    assign weights1[24][765] = 16'b1111111111111000;
    assign weights1[24][766] = 16'b1111111111110011;
    assign weights1[24][767] = 16'b1111111111110011;
    assign weights1[24][768] = 16'b0000000000000100;
    assign weights1[24][769] = 16'b1111111111111010;
    assign weights1[24][770] = 16'b1111111111111100;
    assign weights1[24][771] = 16'b1111111111111111;
    assign weights1[24][772] = 16'b1111111111111111;
    assign weights1[24][773] = 16'b1111111111111110;
    assign weights1[24][774] = 16'b1111111111111000;
    assign weights1[24][775] = 16'b1111111111101101;
    assign weights1[24][776] = 16'b1111111111101011;
    assign weights1[24][777] = 16'b1111111111110101;
    assign weights1[24][778] = 16'b1111111111110011;
    assign weights1[24][779] = 16'b1111111111111010;
    assign weights1[24][780] = 16'b1111111111110111;
    assign weights1[24][781] = 16'b1111111111111000;
    assign weights1[24][782] = 16'b1111111111111001;
    assign weights1[24][783] = 16'b0000000000000100;
    assign weights1[25][0] = 16'b0000000000000000;
    assign weights1[25][1] = 16'b0000000000000000;
    assign weights1[25][2] = 16'b1111111111111110;
    assign weights1[25][3] = 16'b1111111111111110;
    assign weights1[25][4] = 16'b1111111111111110;
    assign weights1[25][5] = 16'b1111111111110111;
    assign weights1[25][6] = 16'b1111111111110000;
    assign weights1[25][7] = 16'b1111111111100110;
    assign weights1[25][8] = 16'b1111111111100100;
    assign weights1[25][9] = 16'b1111111111011011;
    assign weights1[25][10] = 16'b1111111111001110;
    assign weights1[25][11] = 16'b1111111111010100;
    assign weights1[25][12] = 16'b1111111111011000;
    assign weights1[25][13] = 16'b1111111111100111;
    assign weights1[25][14] = 16'b1111111111100100;
    assign weights1[25][15] = 16'b1111111111111100;
    assign weights1[25][16] = 16'b0000000000001110;
    assign weights1[25][17] = 16'b0000000000000111;
    assign weights1[25][18] = 16'b0000000000011011;
    assign weights1[25][19] = 16'b0000000000010000;
    assign weights1[25][20] = 16'b0000000000011001;
    assign weights1[25][21] = 16'b0000000000010010;
    assign weights1[25][22] = 16'b0000000000011111;
    assign weights1[25][23] = 16'b0000000000011111;
    assign weights1[25][24] = 16'b0000000000011001;
    assign weights1[25][25] = 16'b0000000000010010;
    assign weights1[25][26] = 16'b0000000000001010;
    assign weights1[25][27] = 16'b0000000000000101;
    assign weights1[25][28] = 16'b0000000000000000;
    assign weights1[25][29] = 16'b1111111111111110;
    assign weights1[25][30] = 16'b1111111111111100;
    assign weights1[25][31] = 16'b1111111111111100;
    assign weights1[25][32] = 16'b1111111111110101;
    assign weights1[25][33] = 16'b1111111111110110;
    assign weights1[25][34] = 16'b1111111111101001;
    assign weights1[25][35] = 16'b1111111111011111;
    assign weights1[25][36] = 16'b1111111111010110;
    assign weights1[25][37] = 16'b1111111111001110;
    assign weights1[25][38] = 16'b1111111111010001;
    assign weights1[25][39] = 16'b1111111111101010;
    assign weights1[25][40] = 16'b1111111111100110;
    assign weights1[25][41] = 16'b1111111111110111;
    assign weights1[25][42] = 16'b1111111111111110;
    assign weights1[25][43] = 16'b0000000000000100;
    assign weights1[25][44] = 16'b0000000000010110;
    assign weights1[25][45] = 16'b0000000000010011;
    assign weights1[25][46] = 16'b0000000000010101;
    assign weights1[25][47] = 16'b0000000000010110;
    assign weights1[25][48] = 16'b0000000000010101;
    assign weights1[25][49] = 16'b0000000000100000;
    assign weights1[25][50] = 16'b0000000000011110;
    assign weights1[25][51] = 16'b0000000000011100;
    assign weights1[25][52] = 16'b0000000000011101;
    assign weights1[25][53] = 16'b0000000000010101;
    assign weights1[25][54] = 16'b0000000000001001;
    assign weights1[25][55] = 16'b0000000000000011;
    assign weights1[25][56] = 16'b0000000000000000;
    assign weights1[25][57] = 16'b1111111111111100;
    assign weights1[25][58] = 16'b1111111111111001;
    assign weights1[25][59] = 16'b1111111111110111;
    assign weights1[25][60] = 16'b1111111111101111;
    assign weights1[25][61] = 16'b1111111111110000;
    assign weights1[25][62] = 16'b1111111111100010;
    assign weights1[25][63] = 16'b1111111111011101;
    assign weights1[25][64] = 16'b1111111111011001;
    assign weights1[25][65] = 16'b1111111111001110;
    assign weights1[25][66] = 16'b1111111111100111;
    assign weights1[25][67] = 16'b1111111111101111;
    assign weights1[25][68] = 16'b0000000000000010;
    assign weights1[25][69] = 16'b1111111111110101;
    assign weights1[25][70] = 16'b0000000000000110;
    assign weights1[25][71] = 16'b0000000000010111;
    assign weights1[25][72] = 16'b1111111111111101;
    assign weights1[25][73] = 16'b0000000000011011;
    assign weights1[25][74] = 16'b0000000000001110;
    assign weights1[25][75] = 16'b0000000000011001;
    assign weights1[25][76] = 16'b0000000000101010;
    assign weights1[25][77] = 16'b0000000000100001;
    assign weights1[25][78] = 16'b0000000000100100;
    assign weights1[25][79] = 16'b0000000000100111;
    assign weights1[25][80] = 16'b0000000000011011;
    assign weights1[25][81] = 16'b0000000000010010;
    assign weights1[25][82] = 16'b0000000000010001;
    assign weights1[25][83] = 16'b0000000000000110;
    assign weights1[25][84] = 16'b1111111111111110;
    assign weights1[25][85] = 16'b1111111111111010;
    assign weights1[25][86] = 16'b1111111111110100;
    assign weights1[25][87] = 16'b1111111111101110;
    assign weights1[25][88] = 16'b1111111111101000;
    assign weights1[25][89] = 16'b1111111111110000;
    assign weights1[25][90] = 16'b1111111111100100;
    assign weights1[25][91] = 16'b1111111111010101;
    assign weights1[25][92] = 16'b1111111111110010;
    assign weights1[25][93] = 16'b1111111111101000;
    assign weights1[25][94] = 16'b0000000000000111;
    assign weights1[25][95] = 16'b0000000000010000;
    assign weights1[25][96] = 16'b1111111111111110;
    assign weights1[25][97] = 16'b0000000000001000;
    assign weights1[25][98] = 16'b1111111111111100;
    assign weights1[25][99] = 16'b0000000000001011;
    assign weights1[25][100] = 16'b0000000000001010;
    assign weights1[25][101] = 16'b0000000000010011;
    assign weights1[25][102] = 16'b0000000000011010;
    assign weights1[25][103] = 16'b0000000000001001;
    assign weights1[25][104] = 16'b0000000000010011;
    assign weights1[25][105] = 16'b0000000000011010;
    assign weights1[25][106] = 16'b0000000000011011;
    assign weights1[25][107] = 16'b0000000000010001;
    assign weights1[25][108] = 16'b0000000000001111;
    assign weights1[25][109] = 16'b0000000000001011;
    assign weights1[25][110] = 16'b0000000000010100;
    assign weights1[25][111] = 16'b0000000000001001;
    assign weights1[25][112] = 16'b1111111111111011;
    assign weights1[25][113] = 16'b1111111111110100;
    assign weights1[25][114] = 16'b1111111111101101;
    assign weights1[25][115] = 16'b1111111111100100;
    assign weights1[25][116] = 16'b1111111111100101;
    assign weights1[25][117] = 16'b1111111111110001;
    assign weights1[25][118] = 16'b1111111111100100;
    assign weights1[25][119] = 16'b1111111111110011;
    assign weights1[25][120] = 16'b1111111111110101;
    assign weights1[25][121] = 16'b0000000000010011;
    assign weights1[25][122] = 16'b0000000000011111;
    assign weights1[25][123] = 16'b0000000000101001;
    assign weights1[25][124] = 16'b1111111111111111;
    assign weights1[25][125] = 16'b0000000000011111;
    assign weights1[25][126] = 16'b0000000000100100;
    assign weights1[25][127] = 16'b0000000000011000;
    assign weights1[25][128] = 16'b0000000000011001;
    assign weights1[25][129] = 16'b0000000000010101;
    assign weights1[25][130] = 16'b0000000000100000;
    assign weights1[25][131] = 16'b0000000000001100;
    assign weights1[25][132] = 16'b0000000000001000;
    assign weights1[25][133] = 16'b0000000000011010;
    assign weights1[25][134] = 16'b0000000000001011;
    assign weights1[25][135] = 16'b0000000000011011;
    assign weights1[25][136] = 16'b0000000000011100;
    assign weights1[25][137] = 16'b0000000000011000;
    assign weights1[25][138] = 16'b0000000000100111;
    assign weights1[25][139] = 16'b0000000000010101;
    assign weights1[25][140] = 16'b1111111111111010;
    assign weights1[25][141] = 16'b1111111111101111;
    assign weights1[25][142] = 16'b1111111111100111;
    assign weights1[25][143] = 16'b1111111111011110;
    assign weights1[25][144] = 16'b1111111111100110;
    assign weights1[25][145] = 16'b1111111111101001;
    assign weights1[25][146] = 16'b1111111111111111;
    assign weights1[25][147] = 16'b1111111111111100;
    assign weights1[25][148] = 16'b0000000000100101;
    assign weights1[25][149] = 16'b0000000000101000;
    assign weights1[25][150] = 16'b0000000000110100;
    assign weights1[25][151] = 16'b0000000000011101;
    assign weights1[25][152] = 16'b0000000000111101;
    assign weights1[25][153] = 16'b0000000000100001;
    assign weights1[25][154] = 16'b0000000000010001;
    assign weights1[25][155] = 16'b0000000000101000;
    assign weights1[25][156] = 16'b0000000000010001;
    assign weights1[25][157] = 16'b0000000000010111;
    assign weights1[25][158] = 16'b0000000000011010;
    assign weights1[25][159] = 16'b0000000000011101;
    assign weights1[25][160] = 16'b0000000000100110;
    assign weights1[25][161] = 16'b0000000000100010;
    assign weights1[25][162] = 16'b0000000000011110;
    assign weights1[25][163] = 16'b0000000000101011;
    assign weights1[25][164] = 16'b0000000000111100;
    assign weights1[25][165] = 16'b0000000000110000;
    assign weights1[25][166] = 16'b0000000000100100;
    assign weights1[25][167] = 16'b0000000000100010;
    assign weights1[25][168] = 16'b1111111111110111;
    assign weights1[25][169] = 16'b1111111111101110;
    assign weights1[25][170] = 16'b1111111111100010;
    assign weights1[25][171] = 16'b1111111111101001;
    assign weights1[25][172] = 16'b1111111111101101;
    assign weights1[25][173] = 16'b1111111111111110;
    assign weights1[25][174] = 16'b1111111111110101;
    assign weights1[25][175] = 16'b0000000000001101;
    assign weights1[25][176] = 16'b0000000000011110;
    assign weights1[25][177] = 16'b0000000001000010;
    assign weights1[25][178] = 16'b0000000001000101;
    assign weights1[25][179] = 16'b0000000001000001;
    assign weights1[25][180] = 16'b0000000000111100;
    assign weights1[25][181] = 16'b0000000000011111;
    assign weights1[25][182] = 16'b0000000000010101;
    assign weights1[25][183] = 16'b0000000000100001;
    assign weights1[25][184] = 16'b0000000001000000;
    assign weights1[25][185] = 16'b0000000000010000;
    assign weights1[25][186] = 16'b0000000000011110;
    assign weights1[25][187] = 16'b0000000000100100;
    assign weights1[25][188] = 16'b0000000000010011;
    assign weights1[25][189] = 16'b0000000000100100;
    assign weights1[25][190] = 16'b0000000000101111;
    assign weights1[25][191] = 16'b0000000000100110;
    assign weights1[25][192] = 16'b0000000000100101;
    assign weights1[25][193] = 16'b0000000000101000;
    assign weights1[25][194] = 16'b0000000000101100;
    assign weights1[25][195] = 16'b0000000000100101;
    assign weights1[25][196] = 16'b1111111111110100;
    assign weights1[25][197] = 16'b1111111111101100;
    assign weights1[25][198] = 16'b1111111111101010;
    assign weights1[25][199] = 16'b1111111111110110;
    assign weights1[25][200] = 16'b1111111111110101;
    assign weights1[25][201] = 16'b0000000000000101;
    assign weights1[25][202] = 16'b0000000000001000;
    assign weights1[25][203] = 16'b0000000000011110;
    assign weights1[25][204] = 16'b0000000000100101;
    assign weights1[25][205] = 16'b0000000000100010;
    assign weights1[25][206] = 16'b0000000000111010;
    assign weights1[25][207] = 16'b0000000001000011;
    assign weights1[25][208] = 16'b0000000001000110;
    assign weights1[25][209] = 16'b0000000000100010;
    assign weights1[25][210] = 16'b0000000000101011;
    assign weights1[25][211] = 16'b0000000000011111;
    assign weights1[25][212] = 16'b0000000000010101;
    assign weights1[25][213] = 16'b0000000000011110;
    assign weights1[25][214] = 16'b0000000000011111;
    assign weights1[25][215] = 16'b0000000000011110;
    assign weights1[25][216] = 16'b0000000000101000;
    assign weights1[25][217] = 16'b0000000000000001;
    assign weights1[25][218] = 16'b0000000000000111;
    assign weights1[25][219] = 16'b1111111111111101;
    assign weights1[25][220] = 16'b0000000000100010;
    assign weights1[25][221] = 16'b0000000000011100;
    assign weights1[25][222] = 16'b0000000000100110;
    assign weights1[25][223] = 16'b0000000000101011;
    assign weights1[25][224] = 16'b1111111111101100;
    assign weights1[25][225] = 16'b1111111111101010;
    assign weights1[25][226] = 16'b1111111111110100;
    assign weights1[25][227] = 16'b1111111111101000;
    assign weights1[25][228] = 16'b1111111111011011;
    assign weights1[25][229] = 16'b0000000000011010;
    assign weights1[25][230] = 16'b0000000000001001;
    assign weights1[25][231] = 16'b0000000000100011;
    assign weights1[25][232] = 16'b0000000000100011;
    assign weights1[25][233] = 16'b0000000000101101;
    assign weights1[25][234] = 16'b0000000001000001;
    assign weights1[25][235] = 16'b0000000001001000;
    assign weights1[25][236] = 16'b0000000000111100;
    assign weights1[25][237] = 16'b0000000000011100;
    assign weights1[25][238] = 16'b0000000001000010;
    assign weights1[25][239] = 16'b0000000001001000;
    assign weights1[25][240] = 16'b0000000000100000;
    assign weights1[25][241] = 16'b0000000000011011;
    assign weights1[25][242] = 16'b0000000000010011;
    assign weights1[25][243] = 16'b1111111111111001;
    assign weights1[25][244] = 16'b0000000000001001;
    assign weights1[25][245] = 16'b1111111111010101;
    assign weights1[25][246] = 16'b0000000000000111;
    assign weights1[25][247] = 16'b0000000000000000;
    assign weights1[25][248] = 16'b0000000000010001;
    assign weights1[25][249] = 16'b0000000000001011;
    assign weights1[25][250] = 16'b0000000000010101;
    assign weights1[25][251] = 16'b0000000000100010;
    assign weights1[25][252] = 16'b1111111111101101;
    assign weights1[25][253] = 16'b1111111111110001;
    assign weights1[25][254] = 16'b1111111111111101;
    assign weights1[25][255] = 16'b0000000000000101;
    assign weights1[25][256] = 16'b1111111111110110;
    assign weights1[25][257] = 16'b0000000000001010;
    assign weights1[25][258] = 16'b0000000000001101;
    assign weights1[25][259] = 16'b0000000000010001;
    assign weights1[25][260] = 16'b0000000000110010;
    assign weights1[25][261] = 16'b0000000000110001;
    assign weights1[25][262] = 16'b0000000001010011;
    assign weights1[25][263] = 16'b0000000000101110;
    assign weights1[25][264] = 16'b0000000000000101;
    assign weights1[25][265] = 16'b1111111111100010;
    assign weights1[25][266] = 16'b1111111111100100;
    assign weights1[25][267] = 16'b0000000000011110;
    assign weights1[25][268] = 16'b0000000000011010;
    assign weights1[25][269] = 16'b1111111111101110;
    assign weights1[25][270] = 16'b1111111111101101;
    assign weights1[25][271] = 16'b1111111111110100;
    assign weights1[25][272] = 16'b1111111111111011;
    assign weights1[25][273] = 16'b1111111111111010;
    assign weights1[25][274] = 16'b1111111111110011;
    assign weights1[25][275] = 16'b1111111111110011;
    assign weights1[25][276] = 16'b0000000000001010;
    assign weights1[25][277] = 16'b0000000000010010;
    assign weights1[25][278] = 16'b0000000000001111;
    assign weights1[25][279] = 16'b0000000000010100;
    assign weights1[25][280] = 16'b1111111111110000;
    assign weights1[25][281] = 16'b1111111111110101;
    assign weights1[25][282] = 16'b0000000000000101;
    assign weights1[25][283] = 16'b0000000000001011;
    assign weights1[25][284] = 16'b0000000000001010;
    assign weights1[25][285] = 16'b0000000000001010;
    assign weights1[25][286] = 16'b0000000000001100;
    assign weights1[25][287] = 16'b0000000000000010;
    assign weights1[25][288] = 16'b0000000000010011;
    assign weights1[25][289] = 16'b0000000000100010;
    assign weights1[25][290] = 16'b0000000001000101;
    assign weights1[25][291] = 16'b0000000000110011;
    assign weights1[25][292] = 16'b1111111111100000;
    assign weights1[25][293] = 16'b1111111110000010;
    assign weights1[25][294] = 16'b1111111110000010;
    assign weights1[25][295] = 16'b1111111111011000;
    assign weights1[25][296] = 16'b1111111111101000;
    assign weights1[25][297] = 16'b1111111111110101;
    assign weights1[25][298] = 16'b1111111111100100;
    assign weights1[25][299] = 16'b1111111111100110;
    assign weights1[25][300] = 16'b1111111111110000;
    assign weights1[25][301] = 16'b1111111111111011;
    assign weights1[25][302] = 16'b1111111111011111;
    assign weights1[25][303] = 16'b0000000000000000;
    assign weights1[25][304] = 16'b1111111111111111;
    assign weights1[25][305] = 16'b0000000000001100;
    assign weights1[25][306] = 16'b0000000000001101;
    assign weights1[25][307] = 16'b0000000000010100;
    assign weights1[25][308] = 16'b1111111111111001;
    assign weights1[25][309] = 16'b0000000000000110;
    assign weights1[25][310] = 16'b0000000000010110;
    assign weights1[25][311] = 16'b0000000000010111;
    assign weights1[25][312] = 16'b0000000000011010;
    assign weights1[25][313] = 16'b0000000000010001;
    assign weights1[25][314] = 16'b0000000000011000;
    assign weights1[25][315] = 16'b0000000000010111;
    assign weights1[25][316] = 16'b0000000000010101;
    assign weights1[25][317] = 16'b0000000000001101;
    assign weights1[25][318] = 16'b0000000000101100;
    assign weights1[25][319] = 16'b0000000000000100;
    assign weights1[25][320] = 16'b1111111110111000;
    assign weights1[25][321] = 16'b1111111101110101;
    assign weights1[25][322] = 16'b1111111101110110;
    assign weights1[25][323] = 16'b1111111111000001;
    assign weights1[25][324] = 16'b0000000000000000;
    assign weights1[25][325] = 16'b1111111111011001;
    assign weights1[25][326] = 16'b1111111111100100;
    assign weights1[25][327] = 16'b1111111111010010;
    assign weights1[25][328] = 16'b1111111111100110;
    assign weights1[25][329] = 16'b1111111111100011;
    assign weights1[25][330] = 16'b1111111111100011;
    assign weights1[25][331] = 16'b1111111111101111;
    assign weights1[25][332] = 16'b1111111111111010;
    assign weights1[25][333] = 16'b1111111111111110;
    assign weights1[25][334] = 16'b0000000000011000;
    assign weights1[25][335] = 16'b0000000000010100;
    assign weights1[25][336] = 16'b1111111111111011;
    assign weights1[25][337] = 16'b0000000000010101;
    assign weights1[25][338] = 16'b0000000000011011;
    assign weights1[25][339] = 16'b0000000000100001;
    assign weights1[25][340] = 16'b0000000000100101;
    assign weights1[25][341] = 16'b0000000000010011;
    assign weights1[25][342] = 16'b0000000000000110;
    assign weights1[25][343] = 16'b0000000000011100;
    assign weights1[25][344] = 16'b0000000000010001;
    assign weights1[25][345] = 16'b0000000000001100;
    assign weights1[25][346] = 16'b0000000000011001;
    assign weights1[25][347] = 16'b0000000000011100;
    assign weights1[25][348] = 16'b1111111111010100;
    assign weights1[25][349] = 16'b1111111110101000;
    assign weights1[25][350] = 16'b1111111110011111;
    assign weights1[25][351] = 16'b1111111111100010;
    assign weights1[25][352] = 16'b1111111111110010;
    assign weights1[25][353] = 16'b1111111111110001;
    assign weights1[25][354] = 16'b1111111111110101;
    assign weights1[25][355] = 16'b1111111111010111;
    assign weights1[25][356] = 16'b1111111111110111;
    assign weights1[25][357] = 16'b1111111111011101;
    assign weights1[25][358] = 16'b1111111111101100;
    assign weights1[25][359] = 16'b1111111111110011;
    assign weights1[25][360] = 16'b1111111111110010;
    assign weights1[25][361] = 16'b0000000000000001;
    assign weights1[25][362] = 16'b0000000000001001;
    assign weights1[25][363] = 16'b0000000000010101;
    assign weights1[25][364] = 16'b1111111111111000;
    assign weights1[25][365] = 16'b0000000000001001;
    assign weights1[25][366] = 16'b0000000000010110;
    assign weights1[25][367] = 16'b0000000000100010;
    assign weights1[25][368] = 16'b0000000000110000;
    assign weights1[25][369] = 16'b0000000000001101;
    assign weights1[25][370] = 16'b0000000000001110;
    assign weights1[25][371] = 16'b0000000000101111;
    assign weights1[25][372] = 16'b1111111111110001;
    assign weights1[25][373] = 16'b0000000000011100;
    assign weights1[25][374] = 16'b0000000000010010;
    assign weights1[25][375] = 16'b0000000000000110;
    assign weights1[25][376] = 16'b1111111111000110;
    assign weights1[25][377] = 16'b1111111110110011;
    assign weights1[25][378] = 16'b1111111110011010;
    assign weights1[25][379] = 16'b1111111110111101;
    assign weights1[25][380] = 16'b1111111111100011;
    assign weights1[25][381] = 16'b1111111111111010;
    assign weights1[25][382] = 16'b1111111111111111;
    assign weights1[25][383] = 16'b1111111111011011;
    assign weights1[25][384] = 16'b1111111111111110;
    assign weights1[25][385] = 16'b1111111111101110;
    assign weights1[25][386] = 16'b1111111111110100;
    assign weights1[25][387] = 16'b1111111111111111;
    assign weights1[25][388] = 16'b1111111111110100;
    assign weights1[25][389] = 16'b1111111111110111;
    assign weights1[25][390] = 16'b0000000000010010;
    assign weights1[25][391] = 16'b0000000000011000;
    assign weights1[25][392] = 16'b0000000000000100;
    assign weights1[25][393] = 16'b0000000000001110;
    assign weights1[25][394] = 16'b0000000000011010;
    assign weights1[25][395] = 16'b0000000000010011;
    assign weights1[25][396] = 16'b0000000000100010;
    assign weights1[25][397] = 16'b0000000000001000;
    assign weights1[25][398] = 16'b1111111111111101;
    assign weights1[25][399] = 16'b0000000000000110;
    assign weights1[25][400] = 16'b0000000000001010;
    assign weights1[25][401] = 16'b0000000000011010;
    assign weights1[25][402] = 16'b0000000000000011;
    assign weights1[25][403] = 16'b1111111111011111;
    assign weights1[25][404] = 16'b1111111111011101;
    assign weights1[25][405] = 16'b1111111110110000;
    assign weights1[25][406] = 16'b1111111110111111;
    assign weights1[25][407] = 16'b1111111111001011;
    assign weights1[25][408] = 16'b1111111111110100;
    assign weights1[25][409] = 16'b1111111111011010;
    assign weights1[25][410] = 16'b1111111111101011;
    assign weights1[25][411] = 16'b1111111111110100;
    assign weights1[25][412] = 16'b1111111111111001;
    assign weights1[25][413] = 16'b0000000000000111;
    assign weights1[25][414] = 16'b1111111111111011;
    assign weights1[25][415] = 16'b1111111111110010;
    assign weights1[25][416] = 16'b1111111111110101;
    assign weights1[25][417] = 16'b1111111111111101;
    assign weights1[25][418] = 16'b0000000000011100;
    assign weights1[25][419] = 16'b0000000000011011;
    assign weights1[25][420] = 16'b1111111111111101;
    assign weights1[25][421] = 16'b0000000000000010;
    assign weights1[25][422] = 16'b0000000000001111;
    assign weights1[25][423] = 16'b0000000000011101;
    assign weights1[25][424] = 16'b1111111111111001;
    assign weights1[25][425] = 16'b0000000000000111;
    assign weights1[25][426] = 16'b1111111111111001;
    assign weights1[25][427] = 16'b0000000000000010;
    assign weights1[25][428] = 16'b0000000000010100;
    assign weights1[25][429] = 16'b1111111111110001;
    assign weights1[25][430] = 16'b0000000000001000;
    assign weights1[25][431] = 16'b1111111111101011;
    assign weights1[25][432] = 16'b1111111111001111;
    assign weights1[25][433] = 16'b1111111111000000;
    assign weights1[25][434] = 16'b1111111110110100;
    assign weights1[25][435] = 16'b1111111111010001;
    assign weights1[25][436] = 16'b1111111111011101;
    assign weights1[25][437] = 16'b1111111111101000;
    assign weights1[25][438] = 16'b1111111111111000;
    assign weights1[25][439] = 16'b0000000000000000;
    assign weights1[25][440] = 16'b0000000000000001;
    assign weights1[25][441] = 16'b0000000000000110;
    assign weights1[25][442] = 16'b1111111111110001;
    assign weights1[25][443] = 16'b1111111111110001;
    assign weights1[25][444] = 16'b1111111111100011;
    assign weights1[25][445] = 16'b1111111111110111;
    assign weights1[25][446] = 16'b0000000000001110;
    assign weights1[25][447] = 16'b0000000000001101;
    assign weights1[25][448] = 16'b1111111111111111;
    assign weights1[25][449] = 16'b0000000000001001;
    assign weights1[25][450] = 16'b0000000000000101;
    assign weights1[25][451] = 16'b0000000000001011;
    assign weights1[25][452] = 16'b1111111111011110;
    assign weights1[25][453] = 16'b0000000000000100;
    assign weights1[25][454] = 16'b1111111111110100;
    assign weights1[25][455] = 16'b1111111111110011;
    assign weights1[25][456] = 16'b1111111111111010;
    assign weights1[25][457] = 16'b1111111111101001;
    assign weights1[25][458] = 16'b1111111111110101;
    assign weights1[25][459] = 16'b1111111111100001;
    assign weights1[25][460] = 16'b1111111111100000;
    assign weights1[25][461] = 16'b1111111110110000;
    assign weights1[25][462] = 16'b1111111111000010;
    assign weights1[25][463] = 16'b1111111111101101;
    assign weights1[25][464] = 16'b1111111111011010;
    assign weights1[25][465] = 16'b1111111111100100;
    assign weights1[25][466] = 16'b1111111111101001;
    assign weights1[25][467] = 16'b1111111111101110;
    assign weights1[25][468] = 16'b1111111111111101;
    assign weights1[25][469] = 16'b0000000000001000;
    assign weights1[25][470] = 16'b0000000000000000;
    assign weights1[25][471] = 16'b1111111111100111;
    assign weights1[25][472] = 16'b1111111111101010;
    assign weights1[25][473] = 16'b1111111111110010;
    assign weights1[25][474] = 16'b1111111111111111;
    assign weights1[25][475] = 16'b0000000000000000;
    assign weights1[25][476] = 16'b0000000000000111;
    assign weights1[25][477] = 16'b0000000000000101;
    assign weights1[25][478] = 16'b0000000000000000;
    assign weights1[25][479] = 16'b0000000000001001;
    assign weights1[25][480] = 16'b1111111111110110;
    assign weights1[25][481] = 16'b0000000000001010;
    assign weights1[25][482] = 16'b1111111111101101;
    assign weights1[25][483] = 16'b1111111111101011;
    assign weights1[25][484] = 16'b1111111111110011;
    assign weights1[25][485] = 16'b1111111111100101;
    assign weights1[25][486] = 16'b1111111111101111;
    assign weights1[25][487] = 16'b1111111111101011;
    assign weights1[25][488] = 16'b1111111111010111;
    assign weights1[25][489] = 16'b1111111111000110;
    assign weights1[25][490] = 16'b1111111110111110;
    assign weights1[25][491] = 16'b1111111111010000;
    assign weights1[25][492] = 16'b0000000000000100;
    assign weights1[25][493] = 16'b1111111111101011;
    assign weights1[25][494] = 16'b0000000000001010;
    assign weights1[25][495] = 16'b1111111111110011;
    assign weights1[25][496] = 16'b0000000000001000;
    assign weights1[25][497] = 16'b1111111111110110;
    assign weights1[25][498] = 16'b1111111111011001;
    assign weights1[25][499] = 16'b1111111111100110;
    assign weights1[25][500] = 16'b1111111111100101;
    assign weights1[25][501] = 16'b1111111111101100;
    assign weights1[25][502] = 16'b1111111111111010;
    assign weights1[25][503] = 16'b1111111111111010;
    assign weights1[25][504] = 16'b0000000000000111;
    assign weights1[25][505] = 16'b0000000000000011;
    assign weights1[25][506] = 16'b1111111111111111;
    assign weights1[25][507] = 16'b0000000000000110;
    assign weights1[25][508] = 16'b1111111111110001;
    assign weights1[25][509] = 16'b0000000000000010;
    assign weights1[25][510] = 16'b1111111111111001;
    assign weights1[25][511] = 16'b1111111111111001;
    assign weights1[25][512] = 16'b1111111111111000;
    assign weights1[25][513] = 16'b1111111111111001;
    assign weights1[25][514] = 16'b1111111111111110;
    assign weights1[25][515] = 16'b1111111111101101;
    assign weights1[25][516] = 16'b1111111111100010;
    assign weights1[25][517] = 16'b1111111111011001;
    assign weights1[25][518] = 16'b1111111111011100;
    assign weights1[25][519] = 16'b1111111111101111;
    assign weights1[25][520] = 16'b1111111111001000;
    assign weights1[25][521] = 16'b1111111111111000;
    assign weights1[25][522] = 16'b0000000000000001;
    assign weights1[25][523] = 16'b0000000000000001;
    assign weights1[25][524] = 16'b1111111111111010;
    assign weights1[25][525] = 16'b1111111111111101;
    assign weights1[25][526] = 16'b0000000000000001;
    assign weights1[25][527] = 16'b1111111111101001;
    assign weights1[25][528] = 16'b1111111111101101;
    assign weights1[25][529] = 16'b1111111111110011;
    assign weights1[25][530] = 16'b1111111111110000;
    assign weights1[25][531] = 16'b1111111111110100;
    assign weights1[25][532] = 16'b0000000000000101;
    assign weights1[25][533] = 16'b0000000000000000;
    assign weights1[25][534] = 16'b1111111111110110;
    assign weights1[25][535] = 16'b0000000000000100;
    assign weights1[25][536] = 16'b1111111111101110;
    assign weights1[25][537] = 16'b1111111111110010;
    assign weights1[25][538] = 16'b1111111111101001;
    assign weights1[25][539] = 16'b1111111111100111;
    assign weights1[25][540] = 16'b1111111111111000;
    assign weights1[25][541] = 16'b1111111111111110;
    assign weights1[25][542] = 16'b1111111111101100;
    assign weights1[25][543] = 16'b1111111111110000;
    assign weights1[25][544] = 16'b1111111111100011;
    assign weights1[25][545] = 16'b1111111111001000;
    assign weights1[25][546] = 16'b1111111111111010;
    assign weights1[25][547] = 16'b1111111111111110;
    assign weights1[25][548] = 16'b1111111111100010;
    assign weights1[25][549] = 16'b0000000000001101;
    assign weights1[25][550] = 16'b0000000000000101;
    assign weights1[25][551] = 16'b1111111111101111;
    assign weights1[25][552] = 16'b0000000000001111;
    assign weights1[25][553] = 16'b1111111111111100;
    assign weights1[25][554] = 16'b1111111111111110;
    assign weights1[25][555] = 16'b1111111111101110;
    assign weights1[25][556] = 16'b1111111111111111;
    assign weights1[25][557] = 16'b1111111111110000;
    assign weights1[25][558] = 16'b1111111111101001;
    assign weights1[25][559] = 16'b1111111111110000;
    assign weights1[25][560] = 16'b0000000000000001;
    assign weights1[25][561] = 16'b1111111111111011;
    assign weights1[25][562] = 16'b1111111111111001;
    assign weights1[25][563] = 16'b0000000000000000;
    assign weights1[25][564] = 16'b0000000000000010;
    assign weights1[25][565] = 16'b0000000000000100;
    assign weights1[25][566] = 16'b1111111111111110;
    assign weights1[25][567] = 16'b1111111111100111;
    assign weights1[25][568] = 16'b0000000000000100;
    assign weights1[25][569] = 16'b1111111111110101;
    assign weights1[25][570] = 16'b1111111111110101;
    assign weights1[25][571] = 16'b1111111111111100;
    assign weights1[25][572] = 16'b1111111111100010;
    assign weights1[25][573] = 16'b1111111111101010;
    assign weights1[25][574] = 16'b1111111111110011;
    assign weights1[25][575] = 16'b1111111111101010;
    assign weights1[25][576] = 16'b0000000000000001;
    assign weights1[25][577] = 16'b0000000000001010;
    assign weights1[25][578] = 16'b0000000000000000;
    assign weights1[25][579] = 16'b0000000000001000;
    assign weights1[25][580] = 16'b1111111111101001;
    assign weights1[25][581] = 16'b0000000000010000;
    assign weights1[25][582] = 16'b1111111111111001;
    assign weights1[25][583] = 16'b1111111111101111;
    assign weights1[25][584] = 16'b1111111111011100;
    assign weights1[25][585] = 16'b1111111111101110;
    assign weights1[25][586] = 16'b1111111111101100;
    assign weights1[25][587] = 16'b1111111111110100;
    assign weights1[25][588] = 16'b0000000000001000;
    assign weights1[25][589] = 16'b0000000000001111;
    assign weights1[25][590] = 16'b0000000000001110;
    assign weights1[25][591] = 16'b1111111111110101;
    assign weights1[25][592] = 16'b1111111111111001;
    assign weights1[25][593] = 16'b1111111111111101;
    assign weights1[25][594] = 16'b1111111111111101;
    assign weights1[25][595] = 16'b1111111111110011;
    assign weights1[25][596] = 16'b1111111111110100;
    assign weights1[25][597] = 16'b0000000000001111;
    assign weights1[25][598] = 16'b0000000000001100;
    assign weights1[25][599] = 16'b0000000000001100;
    assign weights1[25][600] = 16'b0000000000001100;
    assign weights1[25][601] = 16'b1111111111101110;
    assign weights1[25][602] = 16'b0000000000000001;
    assign weights1[25][603] = 16'b0000000000001001;
    assign weights1[25][604] = 16'b0000000000000110;
    assign weights1[25][605] = 16'b1111111111010001;
    assign weights1[25][606] = 16'b1111111111101000;
    assign weights1[25][607] = 16'b1111111111100110;
    assign weights1[25][608] = 16'b1111111111110111;
    assign weights1[25][609] = 16'b1111111111111001;
    assign weights1[25][610] = 16'b1111111111100101;
    assign weights1[25][611] = 16'b1111111111101010;
    assign weights1[25][612] = 16'b1111111111100110;
    assign weights1[25][613] = 16'b1111111111110010;
    assign weights1[25][614] = 16'b1111111111110101;
    assign weights1[25][615] = 16'b1111111111110110;
    assign weights1[25][616] = 16'b0000000000000111;
    assign weights1[25][617] = 16'b0000000000001110;
    assign weights1[25][618] = 16'b0000000000001001;
    assign weights1[25][619] = 16'b1111111111110111;
    assign weights1[25][620] = 16'b1111111111110111;
    assign weights1[25][621] = 16'b1111111111110001;
    assign weights1[25][622] = 16'b1111111111100001;
    assign weights1[25][623] = 16'b1111111111110110;
    assign weights1[25][624] = 16'b0000000000000111;
    assign weights1[25][625] = 16'b1111111111110010;
    assign weights1[25][626] = 16'b0000000000000001;
    assign weights1[25][627] = 16'b1111111111101101;
    assign weights1[25][628] = 16'b1111111111111110;
    assign weights1[25][629] = 16'b0000000000011000;
    assign weights1[25][630] = 16'b0000000000010101;
    assign weights1[25][631] = 16'b0000000000000110;
    assign weights1[25][632] = 16'b0000000000010110;
    assign weights1[25][633] = 16'b1111111111101111;
    assign weights1[25][634] = 16'b0000000000001110;
    assign weights1[25][635] = 16'b1111111111100010;
    assign weights1[25][636] = 16'b0000000000000101;
    assign weights1[25][637] = 16'b1111111111110111;
    assign weights1[25][638] = 16'b1111111111101011;
    assign weights1[25][639] = 16'b1111111111011011;
    assign weights1[25][640] = 16'b1111111111011011;
    assign weights1[25][641] = 16'b1111111111100110;
    assign weights1[25][642] = 16'b1111111111110011;
    assign weights1[25][643] = 16'b1111111111111000;
    assign weights1[25][644] = 16'b0000000000001000;
    assign weights1[25][645] = 16'b0000000000001001;
    assign weights1[25][646] = 16'b1111111111111111;
    assign weights1[25][647] = 16'b0000000000000100;
    assign weights1[25][648] = 16'b1111111111111111;
    assign weights1[25][649] = 16'b1111111111111110;
    assign weights1[25][650] = 16'b1111111111101010;
    assign weights1[25][651] = 16'b1111111111110111;
    assign weights1[25][652] = 16'b1111111111110011;
    assign weights1[25][653] = 16'b1111111111101011;
    assign weights1[25][654] = 16'b1111111111111101;
    assign weights1[25][655] = 16'b1111111111111010;
    assign weights1[25][656] = 16'b1111111111111011;
    assign weights1[25][657] = 16'b1111111111111010;
    assign weights1[25][658] = 16'b0000000000011111;
    assign weights1[25][659] = 16'b1111111111101100;
    assign weights1[25][660] = 16'b0000000000000111;
    assign weights1[25][661] = 16'b1111111111111110;
    assign weights1[25][662] = 16'b1111111111101110;
    assign weights1[25][663] = 16'b1111111111110011;
    assign weights1[25][664] = 16'b1111111111100111;
    assign weights1[25][665] = 16'b1111111111101101;
    assign weights1[25][666] = 16'b1111111111110110;
    assign weights1[25][667] = 16'b1111111111100110;
    assign weights1[25][668] = 16'b1111111111100011;
    assign weights1[25][669] = 16'b1111111111101110;
    assign weights1[25][670] = 16'b1111111111110110;
    assign weights1[25][671] = 16'b1111111111111010;
    assign weights1[25][672] = 16'b0000000000000111;
    assign weights1[25][673] = 16'b0000000000001011;
    assign weights1[25][674] = 16'b0000000000001011;
    assign weights1[25][675] = 16'b0000000000001001;
    assign weights1[25][676] = 16'b0000000000001101;
    assign weights1[25][677] = 16'b1111111111111111;
    assign weights1[25][678] = 16'b1111111111110110;
    assign weights1[25][679] = 16'b1111111111101001;
    assign weights1[25][680] = 16'b1111111111101110;
    assign weights1[25][681] = 16'b0000000000000000;
    assign weights1[25][682] = 16'b1111111111101101;
    assign weights1[25][683] = 16'b0000000000000000;
    assign weights1[25][684] = 16'b1111111111111011;
    assign weights1[25][685] = 16'b0000000000001011;
    assign weights1[25][686] = 16'b1111111111110011;
    assign weights1[25][687] = 16'b0000000000000010;
    assign weights1[25][688] = 16'b1111111111110010;
    assign weights1[25][689] = 16'b0000000000001101;
    assign weights1[25][690] = 16'b1111111111110110;
    assign weights1[25][691] = 16'b1111111111100011;
    assign weights1[25][692] = 16'b1111111111011111;
    assign weights1[25][693] = 16'b1111111111101011;
    assign weights1[25][694] = 16'b1111111111100100;
    assign weights1[25][695] = 16'b1111111111011110;
    assign weights1[25][696] = 16'b1111111111101101;
    assign weights1[25][697] = 16'b1111111111110001;
    assign weights1[25][698] = 16'b1111111111111100;
    assign weights1[25][699] = 16'b1111111111111110;
    assign weights1[25][700] = 16'b0000000000000011;
    assign weights1[25][701] = 16'b0000000000000001;
    assign weights1[25][702] = 16'b0000000000001101;
    assign weights1[25][703] = 16'b0000000000010000;
    assign weights1[25][704] = 16'b0000000000010100;
    assign weights1[25][705] = 16'b1111111111110110;
    assign weights1[25][706] = 16'b0000000000000111;
    assign weights1[25][707] = 16'b0000000000000001;
    assign weights1[25][708] = 16'b1111111111110011;
    assign weights1[25][709] = 16'b1111111111101111;
    assign weights1[25][710] = 16'b1111111111100111;
    assign weights1[25][711] = 16'b1111111111111010;
    assign weights1[25][712] = 16'b0000000000000011;
    assign weights1[25][713] = 16'b0000000000000100;
    assign weights1[25][714] = 16'b0000000000000000;
    assign weights1[25][715] = 16'b0000000000010100;
    assign weights1[25][716] = 16'b1111111111110001;
    assign weights1[25][717] = 16'b1111111111110110;
    assign weights1[25][718] = 16'b1111111111110111;
    assign weights1[25][719] = 16'b1111111111100110;
    assign weights1[25][720] = 16'b1111111111100000;
    assign weights1[25][721] = 16'b1111111111101001;
    assign weights1[25][722] = 16'b1111111111101010;
    assign weights1[25][723] = 16'b1111111111101100;
    assign weights1[25][724] = 16'b1111111111110100;
    assign weights1[25][725] = 16'b1111111111111010;
    assign weights1[25][726] = 16'b1111111111111100;
    assign weights1[25][727] = 16'b1111111111111101;
    assign weights1[25][728] = 16'b0000000000000010;
    assign weights1[25][729] = 16'b0000000000000000;
    assign weights1[25][730] = 16'b0000000000000000;
    assign weights1[25][731] = 16'b0000000000000110;
    assign weights1[25][732] = 16'b0000000000001101;
    assign weights1[25][733] = 16'b0000000000000010;
    assign weights1[25][734] = 16'b0000000000001110;
    assign weights1[25][735] = 16'b0000000000010001;
    assign weights1[25][736] = 16'b0000000000010011;
    assign weights1[25][737] = 16'b0000000000010011;
    assign weights1[25][738] = 16'b0000000000001110;
    assign weights1[25][739] = 16'b0000000000100011;
    assign weights1[25][740] = 16'b0000000000001111;
    assign weights1[25][741] = 16'b0000000000011100;
    assign weights1[25][742] = 16'b0000000000010010;
    assign weights1[25][743] = 16'b0000000000001011;
    assign weights1[25][744] = 16'b0000000000000110;
    assign weights1[25][745] = 16'b0000000000001000;
    assign weights1[25][746] = 16'b1111111111111011;
    assign weights1[25][747] = 16'b0000000000000011;
    assign weights1[25][748] = 16'b1111111111111010;
    assign weights1[25][749] = 16'b1111111111110010;
    assign weights1[25][750] = 16'b1111111111110000;
    assign weights1[25][751] = 16'b1111111111110010;
    assign weights1[25][752] = 16'b1111111111110110;
    assign weights1[25][753] = 16'b1111111111111101;
    assign weights1[25][754] = 16'b0000000000000000;
    assign weights1[25][755] = 16'b0000000000000000;
    assign weights1[25][756] = 16'b0000000000000001;
    assign weights1[25][757] = 16'b0000000000000000;
    assign weights1[25][758] = 16'b1111111111111100;
    assign weights1[25][759] = 16'b1111111111111010;
    assign weights1[25][760] = 16'b0000000000000000;
    assign weights1[25][761] = 16'b1111111111111101;
    assign weights1[25][762] = 16'b0000000000000010;
    assign weights1[25][763] = 16'b0000000000001101;
    assign weights1[25][764] = 16'b0000000000001100;
    assign weights1[25][765] = 16'b0000000000010010;
    assign weights1[25][766] = 16'b0000000000000011;
    assign weights1[25][767] = 16'b0000000000000101;
    assign weights1[25][768] = 16'b0000000000000000;
    assign weights1[25][769] = 16'b0000000000000010;
    assign weights1[25][770] = 16'b0000000000001000;
    assign weights1[25][771] = 16'b0000000000001000;
    assign weights1[25][772] = 16'b1111111111111100;
    assign weights1[25][773] = 16'b1111111111111100;
    assign weights1[25][774] = 16'b1111111111110011;
    assign weights1[25][775] = 16'b1111111111111011;
    assign weights1[25][776] = 16'b1111111111111000;
    assign weights1[25][777] = 16'b1111111111110100;
    assign weights1[25][778] = 16'b1111111111110011;
    assign weights1[25][779] = 16'b1111111111111010;
    assign weights1[25][780] = 16'b1111111111111111;
    assign weights1[25][781] = 16'b0000000000000000;
    assign weights1[25][782] = 16'b0000000000000000;
    assign weights1[25][783] = 16'b0000000000000000;
    assign weights1[26][0] = 16'b1111111111111111;
    assign weights1[26][1] = 16'b1111111111111111;
    assign weights1[26][2] = 16'b1111111111111110;
    assign weights1[26][3] = 16'b1111111111111111;
    assign weights1[26][4] = 16'b0000000000000001;
    assign weights1[26][5] = 16'b1111111111111110;
    assign weights1[26][6] = 16'b0000000000000001;
    assign weights1[26][7] = 16'b1111111111111101;
    assign weights1[26][8] = 16'b1111111111101110;
    assign weights1[26][9] = 16'b1111111111101111;
    assign weights1[26][10] = 16'b1111111111110011;
    assign weights1[26][11] = 16'b1111111111110011;
    assign weights1[26][12] = 16'b1111111111101010;
    assign weights1[26][13] = 16'b1111111111111001;
    assign weights1[26][14] = 16'b1111111111101011;
    assign weights1[26][15] = 16'b1111111111110011;
    assign weights1[26][16] = 16'b1111111111101011;
    assign weights1[26][17] = 16'b1111111111101010;
    assign weights1[26][18] = 16'b1111111111101011;
    assign weights1[26][19] = 16'b1111111111101101;
    assign weights1[26][20] = 16'b1111111111101100;
    assign weights1[26][21] = 16'b1111111111101110;
    assign weights1[26][22] = 16'b1111111111110011;
    assign weights1[26][23] = 16'b1111111111110010;
    assign weights1[26][24] = 16'b1111111111110001;
    assign weights1[26][25] = 16'b1111111111111010;
    assign weights1[26][26] = 16'b1111111111111100;
    assign weights1[26][27] = 16'b1111111111111110;
    assign weights1[26][28] = 16'b1111111111111110;
    assign weights1[26][29] = 16'b1111111111111110;
    assign weights1[26][30] = 16'b1111111111111110;
    assign weights1[26][31] = 16'b1111111111111010;
    assign weights1[26][32] = 16'b0000000000000001;
    assign weights1[26][33] = 16'b0000000000000010;
    assign weights1[26][34] = 16'b0000000000000111;
    assign weights1[26][35] = 16'b0000000000000000;
    assign weights1[26][36] = 16'b1111111111111101;
    assign weights1[26][37] = 16'b1111111111110000;
    assign weights1[26][38] = 16'b1111111111101111;
    assign weights1[26][39] = 16'b1111111111101110;
    assign weights1[26][40] = 16'b1111111111111111;
    assign weights1[26][41] = 16'b1111111111111011;
    assign weights1[26][42] = 16'b1111111111111111;
    assign weights1[26][43] = 16'b1111111111101011;
    assign weights1[26][44] = 16'b0000000000000010;
    assign weights1[26][45] = 16'b1111111111100011;
    assign weights1[26][46] = 16'b1111111111011101;
    assign weights1[26][47] = 16'b1111111111110001;
    assign weights1[26][48] = 16'b1111111111101011;
    assign weights1[26][49] = 16'b1111111111100000;
    assign weights1[26][50] = 16'b1111111111101010;
    assign weights1[26][51] = 16'b1111111111110101;
    assign weights1[26][52] = 16'b1111111111110010;
    assign weights1[26][53] = 16'b1111111111110100;
    assign weights1[26][54] = 16'b1111111111110011;
    assign weights1[26][55] = 16'b1111111111111100;
    assign weights1[26][56] = 16'b1111111111111101;
    assign weights1[26][57] = 16'b0000000000000000;
    assign weights1[26][58] = 16'b0000000000000001;
    assign weights1[26][59] = 16'b1111111111111111;
    assign weights1[26][60] = 16'b0000000000000010;
    assign weights1[26][61] = 16'b0000000000000100;
    assign weights1[26][62] = 16'b0000000000010001;
    assign weights1[26][63] = 16'b1111111111111100;
    assign weights1[26][64] = 16'b0000000000000011;
    assign weights1[26][65] = 16'b0000000000001100;
    assign weights1[26][66] = 16'b0000000000001110;
    assign weights1[26][67] = 16'b0000000000000000;
    assign weights1[26][68] = 16'b1111111111111010;
    assign weights1[26][69] = 16'b0000000000001011;
    assign weights1[26][70] = 16'b0000000000000101;
    assign weights1[26][71] = 16'b1111111111111011;
    assign weights1[26][72] = 16'b0000000000000011;
    assign weights1[26][73] = 16'b1111111111111001;
    assign weights1[26][74] = 16'b1111111111100000;
    assign weights1[26][75] = 16'b1111111111110100;
    assign weights1[26][76] = 16'b1111111111101110;
    assign weights1[26][77] = 16'b1111111111100011;
    assign weights1[26][78] = 16'b1111111111110101;
    assign weights1[26][79] = 16'b1111111111101101;
    assign weights1[26][80] = 16'b1111111111110100;
    assign weights1[26][81] = 16'b1111111111111001;
    assign weights1[26][82] = 16'b1111111111110001;
    assign weights1[26][83] = 16'b1111111111110101;
    assign weights1[26][84] = 16'b1111111111111110;
    assign weights1[26][85] = 16'b0000000000000010;
    assign weights1[26][86] = 16'b1111111111111111;
    assign weights1[26][87] = 16'b0000000000000101;
    assign weights1[26][88] = 16'b0000000000001011;
    assign weights1[26][89] = 16'b1111111111111001;
    assign weights1[26][90] = 16'b1111111111111100;
    assign weights1[26][91] = 16'b1111111111111111;
    assign weights1[26][92] = 16'b1111111111111001;
    assign weights1[26][93] = 16'b1111111111110011;
    assign weights1[26][94] = 16'b1111111111110100;
    assign weights1[26][95] = 16'b0000000000001010;
    assign weights1[26][96] = 16'b1111111111110000;
    assign weights1[26][97] = 16'b1111111111110011;
    assign weights1[26][98] = 16'b1111111111011111;
    assign weights1[26][99] = 16'b1111111111111111;
    assign weights1[26][100] = 16'b1111111111111100;
    assign weights1[26][101] = 16'b1111111111110110;
    assign weights1[26][102] = 16'b1111111111111111;
    assign weights1[26][103] = 16'b0000000000000100;
    assign weights1[26][104] = 16'b1111111111101010;
    assign weights1[26][105] = 16'b1111111111110011;
    assign weights1[26][106] = 16'b1111111111101001;
    assign weights1[26][107] = 16'b1111111111100110;
    assign weights1[26][108] = 16'b1111111111101011;
    assign weights1[26][109] = 16'b1111111111101110;
    assign weights1[26][110] = 16'b1111111111100111;
    assign weights1[26][111] = 16'b1111111111110110;
    assign weights1[26][112] = 16'b0000000000000000;
    assign weights1[26][113] = 16'b0000000000000110;
    assign weights1[26][114] = 16'b1111111111111100;
    assign weights1[26][115] = 16'b1111111111111101;
    assign weights1[26][116] = 16'b1111111111101110;
    assign weights1[26][117] = 16'b1111111111110110;
    assign weights1[26][118] = 16'b1111111111101101;
    assign weights1[26][119] = 16'b1111111111111100;
    assign weights1[26][120] = 16'b1111111111111100;
    assign weights1[26][121] = 16'b0000000000001011;
    assign weights1[26][122] = 16'b0000000000000110;
    assign weights1[26][123] = 16'b1111111111111010;
    assign weights1[26][124] = 16'b0000000000101100;
    assign weights1[26][125] = 16'b1111111111111100;
    assign weights1[26][126] = 16'b0000000000000010;
    assign weights1[26][127] = 16'b0000000000000101;
    assign weights1[26][128] = 16'b1111111111101110;
    assign weights1[26][129] = 16'b1111111111100111;
    assign weights1[26][130] = 16'b1111111111101111;
    assign weights1[26][131] = 16'b1111111111101111;
    assign weights1[26][132] = 16'b0000000000000001;
    assign weights1[26][133] = 16'b1111111111110101;
    assign weights1[26][134] = 16'b1111111111110100;
    assign weights1[26][135] = 16'b1111111111101011;
    assign weights1[26][136] = 16'b0000000000001001;
    assign weights1[26][137] = 16'b1111111111110010;
    assign weights1[26][138] = 16'b1111111111110001;
    assign weights1[26][139] = 16'b1111111111111011;
    assign weights1[26][140] = 16'b0000000000000010;
    assign weights1[26][141] = 16'b1111111111111110;
    assign weights1[26][142] = 16'b1111111111111101;
    assign weights1[26][143] = 16'b1111111111111100;
    assign weights1[26][144] = 16'b1111111111110111;
    assign weights1[26][145] = 16'b1111111111101110;
    assign weights1[26][146] = 16'b0000000000000010;
    assign weights1[26][147] = 16'b1111111111110000;
    assign weights1[26][148] = 16'b1111111111111011;
    assign weights1[26][149] = 16'b0000000000000101;
    assign weights1[26][150] = 16'b1111111111111010;
    assign weights1[26][151] = 16'b1111111111110111;
    assign weights1[26][152] = 16'b1111111111111001;
    assign weights1[26][153] = 16'b1111111111111001;
    assign weights1[26][154] = 16'b0000000000000011;
    assign weights1[26][155] = 16'b0000000000010111;
    assign weights1[26][156] = 16'b1111111111110110;
    assign weights1[26][157] = 16'b1111111111110010;
    assign weights1[26][158] = 16'b0000000000010000;
    assign weights1[26][159] = 16'b0000000000000001;
    assign weights1[26][160] = 16'b0000000000000011;
    assign weights1[26][161] = 16'b0000000000000100;
    assign weights1[26][162] = 16'b0000000000100101;
    assign weights1[26][163] = 16'b0000000000000011;
    assign weights1[26][164] = 16'b0000000000000010;
    assign weights1[26][165] = 16'b1111111111111110;
    assign weights1[26][166] = 16'b1111111111111101;
    assign weights1[26][167] = 16'b0000000000000010;
    assign weights1[26][168] = 16'b1111111111111111;
    assign weights1[26][169] = 16'b1111111111110100;
    assign weights1[26][170] = 16'b1111111111110111;
    assign weights1[26][171] = 16'b1111111111101111;
    assign weights1[26][172] = 16'b1111111111110111;
    assign weights1[26][173] = 16'b1111111111111101;
    assign weights1[26][174] = 16'b1111111111110110;
    assign weights1[26][175] = 16'b1111111111111000;
    assign weights1[26][176] = 16'b0000000000000001;
    assign weights1[26][177] = 16'b1111111111011001;
    assign weights1[26][178] = 16'b1111111111101001;
    assign weights1[26][179] = 16'b1111111111110000;
    assign weights1[26][180] = 16'b0000000000001011;
    assign weights1[26][181] = 16'b1111111111101011;
    assign weights1[26][182] = 16'b1111111111111001;
    assign weights1[26][183] = 16'b1111111111101100;
    assign weights1[26][184] = 16'b0000000000000001;
    assign weights1[26][185] = 16'b1111111111111000;
    assign weights1[26][186] = 16'b1111111111110110;
    assign weights1[26][187] = 16'b1111111111110000;
    assign weights1[26][188] = 16'b1111111111101110;
    assign weights1[26][189] = 16'b0000000000000100;
    assign weights1[26][190] = 16'b1111111111101100;
    assign weights1[26][191] = 16'b1111111111110001;
    assign weights1[26][192] = 16'b1111111111111101;
    assign weights1[26][193] = 16'b1111111111101001;
    assign weights1[26][194] = 16'b1111111111111001;
    assign weights1[26][195] = 16'b1111111111111101;
    assign weights1[26][196] = 16'b1111111111111010;
    assign weights1[26][197] = 16'b1111111111110001;
    assign weights1[26][198] = 16'b1111111111111001;
    assign weights1[26][199] = 16'b1111111111011110;
    assign weights1[26][200] = 16'b1111111111100110;
    assign weights1[26][201] = 16'b1111111111101001;
    assign weights1[26][202] = 16'b1111111111101011;
    assign weights1[26][203] = 16'b1111111111100111;
    assign weights1[26][204] = 16'b1111111111111000;
    assign weights1[26][205] = 16'b1111111111100101;
    assign weights1[26][206] = 16'b1111111111100010;
    assign weights1[26][207] = 16'b1111111111101100;
    assign weights1[26][208] = 16'b1111111111010101;
    assign weights1[26][209] = 16'b1111111111101001;
    assign weights1[26][210] = 16'b1111111111110101;
    assign weights1[26][211] = 16'b1111111111101010;
    assign weights1[26][212] = 16'b1111111111101001;
    assign weights1[26][213] = 16'b0000000000001110;
    assign weights1[26][214] = 16'b1111111111111000;
    assign weights1[26][215] = 16'b1111111111101011;
    assign weights1[26][216] = 16'b1111111111110111;
    assign weights1[26][217] = 16'b1111111111101000;
    assign weights1[26][218] = 16'b0000000000011001;
    assign weights1[26][219] = 16'b1111111111100010;
    assign weights1[26][220] = 16'b0000000000000000;
    assign weights1[26][221] = 16'b1111111111110110;
    assign weights1[26][222] = 16'b0000000000000010;
    assign weights1[26][223] = 16'b1111111111100111;
    assign weights1[26][224] = 16'b1111111111110101;
    assign weights1[26][225] = 16'b1111111111101101;
    assign weights1[26][226] = 16'b1111111111110000;
    assign weights1[26][227] = 16'b1111111111101001;
    assign weights1[26][228] = 16'b1111111111101000;
    assign weights1[26][229] = 16'b1111111111011111;
    assign weights1[26][230] = 16'b1111111111101100;
    assign weights1[26][231] = 16'b1111111111110101;
    assign weights1[26][232] = 16'b1111111111011000;
    assign weights1[26][233] = 16'b1111111111010010;
    assign weights1[26][234] = 16'b1111111111111100;
    assign weights1[26][235] = 16'b1111111111100000;
    assign weights1[26][236] = 16'b1111111111110100;
    assign weights1[26][237] = 16'b1111111111110100;
    assign weights1[26][238] = 16'b1111111111011100;
    assign weights1[26][239] = 16'b0000000000000101;
    assign weights1[26][240] = 16'b1111111111111101;
    assign weights1[26][241] = 16'b1111111111100000;
    assign weights1[26][242] = 16'b1111111111111001;
    assign weights1[26][243] = 16'b0000000000001001;
    assign weights1[26][244] = 16'b0000000000001110;
    assign weights1[26][245] = 16'b1111111111110001;
    assign weights1[26][246] = 16'b1111111111111100;
    assign weights1[26][247] = 16'b1111111111111011;
    assign weights1[26][248] = 16'b0000000000000010;
    assign weights1[26][249] = 16'b0000000000001111;
    assign weights1[26][250] = 16'b1111111111110100;
    assign weights1[26][251] = 16'b1111111111100110;
    assign weights1[26][252] = 16'b1111111111101110;
    assign weights1[26][253] = 16'b1111111111101010;
    assign weights1[26][254] = 16'b1111111111101000;
    assign weights1[26][255] = 16'b1111111111101001;
    assign weights1[26][256] = 16'b1111111111100000;
    assign weights1[26][257] = 16'b1111111111100111;
    assign weights1[26][258] = 16'b1111111111001101;
    assign weights1[26][259] = 16'b1111111111001000;
    assign weights1[26][260] = 16'b1111111111000100;
    assign weights1[26][261] = 16'b1111111111110001;
    assign weights1[26][262] = 16'b1111111111101101;
    assign weights1[26][263] = 16'b1111111111010010;
    assign weights1[26][264] = 16'b1111111111100000;
    assign weights1[26][265] = 16'b1111111111111110;
    assign weights1[26][266] = 16'b1111111111101100;
    assign weights1[26][267] = 16'b1111111111011010;
    assign weights1[26][268] = 16'b1111111111111010;
    assign weights1[26][269] = 16'b1111111111100100;
    assign weights1[26][270] = 16'b1111111111100111;
    assign weights1[26][271] = 16'b1111111111101010;
    assign weights1[26][272] = 16'b1111111111111011;
    assign weights1[26][273] = 16'b1111111111110010;
    assign weights1[26][274] = 16'b1111111111110101;
    assign weights1[26][275] = 16'b1111111111110000;
    assign weights1[26][276] = 16'b0000000000000010;
    assign weights1[26][277] = 16'b0000000000001110;
    assign weights1[26][278] = 16'b1111111111110001;
    assign weights1[26][279] = 16'b1111111111010110;
    assign weights1[26][280] = 16'b1111111111101100;
    assign weights1[26][281] = 16'b1111111111100000;
    assign weights1[26][282] = 16'b1111111111100111;
    assign weights1[26][283] = 16'b1111111111010101;
    assign weights1[26][284] = 16'b1111111111001111;
    assign weights1[26][285] = 16'b1111111111001111;
    assign weights1[26][286] = 16'b1111111111010101;
    assign weights1[26][287] = 16'b1111111111001111;
    assign weights1[26][288] = 16'b1111111110110100;
    assign weights1[26][289] = 16'b1111111111001110;
    assign weights1[26][290] = 16'b1111111111000110;
    assign weights1[26][291] = 16'b1111111111010111;
    assign weights1[26][292] = 16'b1111111111010011;
    assign weights1[26][293] = 16'b1111111111001111;
    assign weights1[26][294] = 16'b1111111111010111;
    assign weights1[26][295] = 16'b1111111111010100;
    assign weights1[26][296] = 16'b1111111111101011;
    assign weights1[26][297] = 16'b1111111111110000;
    assign weights1[26][298] = 16'b1111111111101111;
    assign weights1[26][299] = 16'b1111111111100110;
    assign weights1[26][300] = 16'b1111111111010000;
    assign weights1[26][301] = 16'b1111111111111101;
    assign weights1[26][302] = 16'b1111111111110000;
    assign weights1[26][303] = 16'b1111111111011101;
    assign weights1[26][304] = 16'b1111111111100000;
    assign weights1[26][305] = 16'b1111111111111010;
    assign weights1[26][306] = 16'b1111111111100010;
    assign weights1[26][307] = 16'b1111111111001111;
    assign weights1[26][308] = 16'b1111111111101100;
    assign weights1[26][309] = 16'b1111111111011111;
    assign weights1[26][310] = 16'b1111111111001010;
    assign weights1[26][311] = 16'b1111111110111011;
    assign weights1[26][312] = 16'b1111111111100000;
    assign weights1[26][313] = 16'b1111111111101100;
    assign weights1[26][314] = 16'b1111111111001110;
    assign weights1[26][315] = 16'b1111111111100111;
    assign weights1[26][316] = 16'b1111111111010010;
    assign weights1[26][317] = 16'b1111111111000000;
    assign weights1[26][318] = 16'b1111111111001011;
    assign weights1[26][319] = 16'b1111111111011011;
    assign weights1[26][320] = 16'b1111111111010100;
    assign weights1[26][321] = 16'b1111111111001011;
    assign weights1[26][322] = 16'b1111111111000011;
    assign weights1[26][323] = 16'b1111111111000010;
    assign weights1[26][324] = 16'b1111111111001100;
    assign weights1[26][325] = 16'b1111111111010011;
    assign weights1[26][326] = 16'b1111111111000001;
    assign weights1[26][327] = 16'b1111111111100000;
    assign weights1[26][328] = 16'b1111111111001110;
    assign weights1[26][329] = 16'b1111111111010100;
    assign weights1[26][330] = 16'b1111111111010010;
    assign weights1[26][331] = 16'b1111111111100010;
    assign weights1[26][332] = 16'b1111111111001111;
    assign weights1[26][333] = 16'b1111111111100001;
    assign weights1[26][334] = 16'b1111111111001100;
    assign weights1[26][335] = 16'b1111111111010010;
    assign weights1[26][336] = 16'b1111111111101011;
    assign weights1[26][337] = 16'b1111111111100100;
    assign weights1[26][338] = 16'b1111111111001111;
    assign weights1[26][339] = 16'b1111111111011001;
    assign weights1[26][340] = 16'b1111111111010100;
    assign weights1[26][341] = 16'b1111111111110111;
    assign weights1[26][342] = 16'b1111111111010100;
    assign weights1[26][343] = 16'b1111111111011011;
    assign weights1[26][344] = 16'b1111111111111010;
    assign weights1[26][345] = 16'b1111111111000111;
    assign weights1[26][346] = 16'b1111111111101001;
    assign weights1[26][347] = 16'b1111111111001100;
    assign weights1[26][348] = 16'b1111111111010111;
    assign weights1[26][349] = 16'b1111111110110101;
    assign weights1[26][350] = 16'b1111111110101110;
    assign weights1[26][351] = 16'b1111111110101100;
    assign weights1[26][352] = 16'b1111111111010101;
    assign weights1[26][353] = 16'b1111111111001010;
    assign weights1[26][354] = 16'b1111111111001010;
    assign weights1[26][355] = 16'b1111111111011010;
    assign weights1[26][356] = 16'b1111111111100110;
    assign weights1[26][357] = 16'b1111111110111111;
    assign weights1[26][358] = 16'b1111111111000010;
    assign weights1[26][359] = 16'b1111111110111011;
    assign weights1[26][360] = 16'b1111111111001101;
    assign weights1[26][361] = 16'b1111111111000001;
    assign weights1[26][362] = 16'b1111111111000001;
    assign weights1[26][363] = 16'b1111111111000100;
    assign weights1[26][364] = 16'b1111111111101110;
    assign weights1[26][365] = 16'b1111111111101110;
    assign weights1[26][366] = 16'b1111111111101011;
    assign weights1[26][367] = 16'b1111111111101101;
    assign weights1[26][368] = 16'b1111111111110001;
    assign weights1[26][369] = 16'b1111111111110000;
    assign weights1[26][370] = 16'b1111111111111010;
    assign weights1[26][371] = 16'b1111111111010110;
    assign weights1[26][372] = 16'b0000000000000100;
    assign weights1[26][373] = 16'b0000000000000011;
    assign weights1[26][374] = 16'b0000000000000001;
    assign weights1[26][375] = 16'b1111111111101101;
    assign weights1[26][376] = 16'b1111111111111000;
    assign weights1[26][377] = 16'b1111111111101110;
    assign weights1[26][378] = 16'b1111111111101101;
    assign weights1[26][379] = 16'b1111111111011111;
    assign weights1[26][380] = 16'b1111111111010111;
    assign weights1[26][381] = 16'b1111111111001001;
    assign weights1[26][382] = 16'b1111111110111110;
    assign weights1[26][383] = 16'b1111111111010000;
    assign weights1[26][384] = 16'b1111111110111111;
    assign weights1[26][385] = 16'b1111111110111001;
    assign weights1[26][386] = 16'b1111111110110101;
    assign weights1[26][387] = 16'b1111111110110011;
    assign weights1[26][388] = 16'b1111111111011000;
    assign weights1[26][389] = 16'b1111111110110111;
    assign weights1[26][390] = 16'b1111111111000100;
    assign weights1[26][391] = 16'b1111111111000100;
    assign weights1[26][392] = 16'b1111111111111011;
    assign weights1[26][393] = 16'b1111111111110101;
    assign weights1[26][394] = 16'b0000000000000100;
    assign weights1[26][395] = 16'b0000000000000111;
    assign weights1[26][396] = 16'b0000000000100010;
    assign weights1[26][397] = 16'b0000000000011011;
    assign weights1[26][398] = 16'b1111111111111110;
    assign weights1[26][399] = 16'b0000000000100001;
    assign weights1[26][400] = 16'b1111111111111011;
    assign weights1[26][401] = 16'b0000000000001010;
    assign weights1[26][402] = 16'b0000000000010000;
    assign weights1[26][403] = 16'b0000000000000001;
    assign weights1[26][404] = 16'b0000000000010100;
    assign weights1[26][405] = 16'b0000000000000010;
    assign weights1[26][406] = 16'b0000000000000011;
    assign weights1[26][407] = 16'b0000000000000111;
    assign weights1[26][408] = 16'b0000000000000111;
    assign weights1[26][409] = 16'b1111111111101101;
    assign weights1[26][410] = 16'b1111111111100001;
    assign weights1[26][411] = 16'b1111111111001000;
    assign weights1[26][412] = 16'b1111111111001111;
    assign weights1[26][413] = 16'b1111111111000001;
    assign weights1[26][414] = 16'b1111111111010101;
    assign weights1[26][415] = 16'b1111111110111101;
    assign weights1[26][416] = 16'b1111111110110001;
    assign weights1[26][417] = 16'b1111111110111000;
    assign weights1[26][418] = 16'b1111111111001000;
    assign weights1[26][419] = 16'b1111111111010000;
    assign weights1[26][420] = 16'b0000000000001011;
    assign weights1[26][421] = 16'b0000000000011010;
    assign weights1[26][422] = 16'b0000000000011010;
    assign weights1[26][423] = 16'b0000000000101111;
    assign weights1[26][424] = 16'b0000000000011011;
    assign weights1[26][425] = 16'b0000000000111001;
    assign weights1[26][426] = 16'b0000000000101110;
    assign weights1[26][427] = 16'b0000000000101111;
    assign weights1[26][428] = 16'b0000000000100001;
    assign weights1[26][429] = 16'b0000000000100100;
    assign weights1[26][430] = 16'b0000000000101010;
    assign weights1[26][431] = 16'b0000000000110011;
    assign weights1[26][432] = 16'b0000000000101010;
    assign weights1[26][433] = 16'b0000000000011011;
    assign weights1[26][434] = 16'b0000000000001010;
    assign weights1[26][435] = 16'b0000000000010000;
    assign weights1[26][436] = 16'b0000000000010011;
    assign weights1[26][437] = 16'b0000000000100011;
    assign weights1[26][438] = 16'b1111111111110100;
    assign weights1[26][439] = 16'b0000000000001100;
    assign weights1[26][440] = 16'b1111111111111001;
    assign weights1[26][441] = 16'b1111111111100101;
    assign weights1[26][442] = 16'b1111111111100100;
    assign weights1[26][443] = 16'b1111111111100000;
    assign weights1[26][444] = 16'b1111111111111100;
    assign weights1[26][445] = 16'b1111111111100111;
    assign weights1[26][446] = 16'b1111111111011111;
    assign weights1[26][447] = 16'b1111111111011010;
    assign weights1[26][448] = 16'b0000000000010011;
    assign weights1[26][449] = 16'b0000000000100010;
    assign weights1[26][450] = 16'b0000000000100110;
    assign weights1[26][451] = 16'b0000000001001001;
    assign weights1[26][452] = 16'b0000000000110111;
    assign weights1[26][453] = 16'b0000000000101011;
    assign weights1[26][454] = 16'b0000000000110110;
    assign weights1[26][455] = 16'b0000000000100111;
    assign weights1[26][456] = 16'b0000000000101111;
    assign weights1[26][457] = 16'b0000000000110110;
    assign weights1[26][458] = 16'b0000000000110100;
    assign weights1[26][459] = 16'b0000000000111000;
    assign weights1[26][460] = 16'b0000000000101010;
    assign weights1[26][461] = 16'b0000000000100111;
    assign weights1[26][462] = 16'b0000000000101100;
    assign weights1[26][463] = 16'b0000000000101111;
    assign weights1[26][464] = 16'b0000000000100001;
    assign weights1[26][465] = 16'b0000000000101010;
    assign weights1[26][466] = 16'b0000000000100001;
    assign weights1[26][467] = 16'b0000000000011010;
    assign weights1[26][468] = 16'b0000000000101011;
    assign weights1[26][469] = 16'b0000000001010001;
    assign weights1[26][470] = 16'b0000000000100110;
    assign weights1[26][471] = 16'b0000000000010101;
    assign weights1[26][472] = 16'b0000000000010110;
    assign weights1[26][473] = 16'b0000000000010010;
    assign weights1[26][474] = 16'b1111111111111100;
    assign weights1[26][475] = 16'b1111111111111101;
    assign weights1[26][476] = 16'b0000000000011110;
    assign weights1[26][477] = 16'b0000000000110011;
    assign weights1[26][478] = 16'b0000000000101100;
    assign weights1[26][479] = 16'b0000000000110111;
    assign weights1[26][480] = 16'b0000000000011111;
    assign weights1[26][481] = 16'b0000000000110010;
    assign weights1[26][482] = 16'b0000000001000000;
    assign weights1[26][483] = 16'b0000000000100110;
    assign weights1[26][484] = 16'b0000000001001001;
    assign weights1[26][485] = 16'b0000000000100110;
    assign weights1[26][486] = 16'b0000000000101111;
    assign weights1[26][487] = 16'b0000000000101010;
    assign weights1[26][488] = 16'b0000000000110010;
    assign weights1[26][489] = 16'b0000000000110011;
    assign weights1[26][490] = 16'b0000000000110101;
    assign weights1[26][491] = 16'b0000000000111010;
    assign weights1[26][492] = 16'b0000000000110111;
    assign weights1[26][493] = 16'b0000000000110110;
    assign weights1[26][494] = 16'b0000000000111010;
    assign weights1[26][495] = 16'b0000000000101010;
    assign weights1[26][496] = 16'b0000000000101100;
    assign weights1[26][497] = 16'b0000000000011011;
    assign weights1[26][498] = 16'b0000000000011110;
    assign weights1[26][499] = 16'b0000000001000000;
    assign weights1[26][500] = 16'b0000000000110111;
    assign weights1[26][501] = 16'b0000000001001110;
    assign weights1[26][502] = 16'b0000000000100001;
    assign weights1[26][503] = 16'b0000000000011001;
    assign weights1[26][504] = 16'b0000000000100101;
    assign weights1[26][505] = 16'b0000000000101100;
    assign weights1[26][506] = 16'b0000000000010110;
    assign weights1[26][507] = 16'b0000000000011110;
    assign weights1[26][508] = 16'b0000000000101001;
    assign weights1[26][509] = 16'b0000000000101110;
    assign weights1[26][510] = 16'b0000000000011101;
    assign weights1[26][511] = 16'b0000000000011010;
    assign weights1[26][512] = 16'b0000000000011000;
    assign weights1[26][513] = 16'b0000000000010001;
    assign weights1[26][514] = 16'b0000000000001100;
    assign weights1[26][515] = 16'b0000000000010110;
    assign weights1[26][516] = 16'b0000000000010111;
    assign weights1[26][517] = 16'b0000000000011001;
    assign weights1[26][518] = 16'b0000000000011011;
    assign weights1[26][519] = 16'b0000000000101010;
    assign weights1[26][520] = 16'b0000000001000110;
    assign weights1[26][521] = 16'b0000000000111111;
    assign weights1[26][522] = 16'b0000000000100101;
    assign weights1[26][523] = 16'b0000000000101101;
    assign weights1[26][524] = 16'b0000000000111100;
    assign weights1[26][525] = 16'b0000000000101001;
    assign weights1[26][526] = 16'b0000000000100110;
    assign weights1[26][527] = 16'b0000000001001101;
    assign weights1[26][528] = 16'b0000000001100001;
    assign weights1[26][529] = 16'b0000000001001000;
    assign weights1[26][530] = 16'b0000000001000011;
    assign weights1[26][531] = 16'b0000000000111100;
    assign weights1[26][532] = 16'b0000000000100001;
    assign weights1[26][533] = 16'b0000000000011101;
    assign weights1[26][534] = 16'b0000000000000111;
    assign weights1[26][535] = 16'b0000000000010011;
    assign weights1[26][536] = 16'b0000000000011100;
    assign weights1[26][537] = 16'b0000000000000111;
    assign weights1[26][538] = 16'b0000000000001101;
    assign weights1[26][539] = 16'b0000000000000011;
    assign weights1[26][540] = 16'b0000000000011000;
    assign weights1[26][541] = 16'b0000000000011010;
    assign weights1[26][542] = 16'b0000000000100000;
    assign weights1[26][543] = 16'b1111111111110111;
    assign weights1[26][544] = 16'b0000000000001011;
    assign weights1[26][545] = 16'b0000000000110011;
    assign weights1[26][546] = 16'b0000000000011010;
    assign weights1[26][547] = 16'b0000000000110011;
    assign weights1[26][548] = 16'b0000000000101111;
    assign weights1[26][549] = 16'b0000000001000101;
    assign weights1[26][550] = 16'b0000000000110111;
    assign weights1[26][551] = 16'b0000000001001001;
    assign weights1[26][552] = 16'b0000000000110000;
    assign weights1[26][553] = 16'b0000000001000011;
    assign weights1[26][554] = 16'b0000000000111111;
    assign weights1[26][555] = 16'b0000000000111000;
    assign weights1[26][556] = 16'b0000000001000100;
    assign weights1[26][557] = 16'b0000000001010110;
    assign weights1[26][558] = 16'b0000000001010100;
    assign weights1[26][559] = 16'b0000000001000000;
    assign weights1[26][560] = 16'b0000000000001001;
    assign weights1[26][561] = 16'b0000000000001100;
    assign weights1[26][562] = 16'b1111111111111101;
    assign weights1[26][563] = 16'b0000000000000010;
    assign weights1[26][564] = 16'b0000000000010010;
    assign weights1[26][565] = 16'b1111111111100000;
    assign weights1[26][566] = 16'b0000000000011000;
    assign weights1[26][567] = 16'b0000000000010000;
    assign weights1[26][568] = 16'b0000000000001011;
    assign weights1[26][569] = 16'b0000000000011011;
    assign weights1[26][570] = 16'b0000000000001000;
    assign weights1[26][571] = 16'b0000000000100001;
    assign weights1[26][572] = 16'b1111111111110101;
    assign weights1[26][573] = 16'b0000000000000100;
    assign weights1[26][574] = 16'b0000000000010000;
    assign weights1[26][575] = 16'b0000000000001010;
    assign weights1[26][576] = 16'b0000000000010101;
    assign weights1[26][577] = 16'b0000000000100000;
    assign weights1[26][578] = 16'b0000000000111101;
    assign weights1[26][579] = 16'b0000000001000001;
    assign weights1[26][580] = 16'b0000000001010110;
    assign weights1[26][581] = 16'b0000000001000000;
    assign weights1[26][582] = 16'b0000000000110001;
    assign weights1[26][583] = 16'b0000000000110111;
    assign weights1[26][584] = 16'b0000000001000110;
    assign weights1[26][585] = 16'b0000000000110110;
    assign weights1[26][586] = 16'b0000000001000100;
    assign weights1[26][587] = 16'b0000000000101000;
    assign weights1[26][588] = 16'b1111111111110100;
    assign weights1[26][589] = 16'b0000000000000111;
    assign weights1[26][590] = 16'b1111111111110001;
    assign weights1[26][591] = 16'b1111111111101011;
    assign weights1[26][592] = 16'b1111111111101110;
    assign weights1[26][593] = 16'b0000000000100101;
    assign weights1[26][594] = 16'b0000000000001110;
    assign weights1[26][595] = 16'b1111111111111011;
    assign weights1[26][596] = 16'b0000000000000101;
    assign weights1[26][597] = 16'b0000000000000111;
    assign weights1[26][598] = 16'b0000000000000110;
    assign weights1[26][599] = 16'b0000000000000010;
    assign weights1[26][600] = 16'b0000000000001000;
    assign weights1[26][601] = 16'b0000000000000011;
    assign weights1[26][602] = 16'b1111111111111011;
    assign weights1[26][603] = 16'b1111111111110011;
    assign weights1[26][604] = 16'b0000000000000010;
    assign weights1[26][605] = 16'b0000000000000001;
    assign weights1[26][606] = 16'b1111111111100000;
    assign weights1[26][607] = 16'b0000000000000110;
    assign weights1[26][608] = 16'b0000000000101100;
    assign weights1[26][609] = 16'b0000000000001101;
    assign weights1[26][610] = 16'b0000000000100011;
    assign weights1[26][611] = 16'b0000000000101001;
    assign weights1[26][612] = 16'b0000000000011101;
    assign weights1[26][613] = 16'b0000000000011010;
    assign weights1[26][614] = 16'b0000000000011010;
    assign weights1[26][615] = 16'b0000000000001001;
    assign weights1[26][616] = 16'b1111111111111000;
    assign weights1[26][617] = 16'b1111111111110111;
    assign weights1[26][618] = 16'b1111111111110001;
    assign weights1[26][619] = 16'b1111111111101110;
    assign weights1[26][620] = 16'b1111111111111101;
    assign weights1[26][621] = 16'b0000000000001011;
    assign weights1[26][622] = 16'b1111111111011111;
    assign weights1[26][623] = 16'b1111111111111010;
    assign weights1[26][624] = 16'b0000000000001000;
    assign weights1[26][625] = 16'b1111111111110000;
    assign weights1[26][626] = 16'b1111111111111101;
    assign weights1[26][627] = 16'b0000000000001011;
    assign weights1[26][628] = 16'b1111111111101101;
    assign weights1[26][629] = 16'b0000000000001010;
    assign weights1[26][630] = 16'b1111111111110010;
    assign weights1[26][631] = 16'b1111111111101100;
    assign weights1[26][632] = 16'b1111111111101000;
    assign weights1[26][633] = 16'b1111111111100110;
    assign weights1[26][634] = 16'b1111111111011010;
    assign weights1[26][635] = 16'b1111111111101011;
    assign weights1[26][636] = 16'b0000000000001000;
    assign weights1[26][637] = 16'b1111111111110110;
    assign weights1[26][638] = 16'b0000000000010001;
    assign weights1[26][639] = 16'b1111111111101111;
    assign weights1[26][640] = 16'b1111111111100110;
    assign weights1[26][641] = 16'b1111111111111000;
    assign weights1[26][642] = 16'b1111111111111000;
    assign weights1[26][643] = 16'b1111111111110111;
    assign weights1[26][644] = 16'b1111111111111001;
    assign weights1[26][645] = 16'b1111111111101010;
    assign weights1[26][646] = 16'b1111111111101110;
    assign weights1[26][647] = 16'b1111111111101011;
    assign weights1[26][648] = 16'b1111111111100011;
    assign weights1[26][649] = 16'b0000000000000000;
    assign weights1[26][650] = 16'b1111111111101110;
    assign weights1[26][651] = 16'b1111111111110001;
    assign weights1[26][652] = 16'b1111111111110110;
    assign weights1[26][653] = 16'b1111111111101010;
    assign weights1[26][654] = 16'b1111111111111001;
    assign weights1[26][655] = 16'b0000000000001001;
    assign weights1[26][656] = 16'b0000000000000000;
    assign weights1[26][657] = 16'b1111111111110100;
    assign weights1[26][658] = 16'b1111111111110011;
    assign weights1[26][659] = 16'b1111111111111000;
    assign weights1[26][660] = 16'b1111111111100100;
    assign weights1[26][661] = 16'b1111111111011110;
    assign weights1[26][662] = 16'b1111111111100101;
    assign weights1[26][663] = 16'b1111111111100101;
    assign weights1[26][664] = 16'b1111111111010110;
    assign weights1[26][665] = 16'b1111111111100111;
    assign weights1[26][666] = 16'b1111111111011100;
    assign weights1[26][667] = 16'b1111111111011101;
    assign weights1[26][668] = 16'b1111111111001111;
    assign weights1[26][669] = 16'b1111111111011101;
    assign weights1[26][670] = 16'b1111111111110001;
    assign weights1[26][671] = 16'b1111111111110100;
    assign weights1[26][672] = 16'b1111111111111001;
    assign weights1[26][673] = 16'b1111111111110001;
    assign weights1[26][674] = 16'b1111111111101110;
    assign weights1[26][675] = 16'b1111111111100100;
    assign weights1[26][676] = 16'b1111111111101110;
    assign weights1[26][677] = 16'b1111111111101101;
    assign weights1[26][678] = 16'b1111111111010001;
    assign weights1[26][679] = 16'b1111111111110010;
    assign weights1[26][680] = 16'b1111111111100111;
    assign weights1[26][681] = 16'b1111111111111010;
    assign weights1[26][682] = 16'b0000000000010010;
    assign weights1[26][683] = 16'b1111111111110000;
    assign weights1[26][684] = 16'b1111111111111011;
    assign weights1[26][685] = 16'b1111111111110001;
    assign weights1[26][686] = 16'b1111111111110000;
    assign weights1[26][687] = 16'b0000000000001111;
    assign weights1[26][688] = 16'b1111111111101110;
    assign weights1[26][689] = 16'b1111111111111011;
    assign weights1[26][690] = 16'b1111111111101110;
    assign weights1[26][691] = 16'b1111111111001100;
    assign weights1[26][692] = 16'b1111111111010110;
    assign weights1[26][693] = 16'b1111111111001001;
    assign weights1[26][694] = 16'b1111111111001010;
    assign weights1[26][695] = 16'b1111111111000101;
    assign weights1[26][696] = 16'b1111111111011011;
    assign weights1[26][697] = 16'b1111111111100010;
    assign weights1[26][698] = 16'b1111111111100110;
    assign weights1[26][699] = 16'b1111111111110011;
    assign weights1[26][700] = 16'b1111111111111101;
    assign weights1[26][701] = 16'b1111111111111000;
    assign weights1[26][702] = 16'b1111111111110011;
    assign weights1[26][703] = 16'b1111111111101101;
    assign weights1[26][704] = 16'b1111111111101000;
    assign weights1[26][705] = 16'b1111111111101001;
    assign weights1[26][706] = 16'b1111111111010100;
    assign weights1[26][707] = 16'b1111111111011010;
    assign weights1[26][708] = 16'b1111111111100011;
    assign weights1[26][709] = 16'b1111111111011011;
    assign weights1[26][710] = 16'b1111111111100101;
    assign weights1[26][711] = 16'b1111111111011011;
    assign weights1[26][712] = 16'b1111111111110111;
    assign weights1[26][713] = 16'b1111111111101010;
    assign weights1[26][714] = 16'b1111111111100010;
    assign weights1[26][715] = 16'b1111111111011010;
    assign weights1[26][716] = 16'b1111111111011111;
    assign weights1[26][717] = 16'b1111111111100110;
    assign weights1[26][718] = 16'b1111111111101101;
    assign weights1[26][719] = 16'b1111111111000001;
    assign weights1[26][720] = 16'b1111111111001100;
    assign weights1[26][721] = 16'b1111111111001010;
    assign weights1[26][722] = 16'b1111111111000110;
    assign weights1[26][723] = 16'b1111111111001011;
    assign weights1[26][724] = 16'b1111111111000110;
    assign weights1[26][725] = 16'b1111111111011100;
    assign weights1[26][726] = 16'b1111111111101010;
    assign weights1[26][727] = 16'b1111111111111000;
    assign weights1[26][728] = 16'b1111111111111100;
    assign weights1[26][729] = 16'b1111111111111011;
    assign weights1[26][730] = 16'b1111111111110101;
    assign weights1[26][731] = 16'b1111111111110010;
    assign weights1[26][732] = 16'b1111111111101011;
    assign weights1[26][733] = 16'b1111111111100110;
    assign weights1[26][734] = 16'b1111111111011001;
    assign weights1[26][735] = 16'b1111111111101001;
    assign weights1[26][736] = 16'b1111111111011101;
    assign weights1[26][737] = 16'b1111111111100111;
    assign weights1[26][738] = 16'b1111111111100101;
    assign weights1[26][739] = 16'b1111111111100110;
    assign weights1[26][740] = 16'b1111111111101010;
    assign weights1[26][741] = 16'b1111111111100000;
    assign weights1[26][742] = 16'b1111111111101100;
    assign weights1[26][743] = 16'b1111111111110001;
    assign weights1[26][744] = 16'b1111111111010110;
    assign weights1[26][745] = 16'b1111111111100111;
    assign weights1[26][746] = 16'b1111111111100100;
    assign weights1[26][747] = 16'b1111111111011100;
    assign weights1[26][748] = 16'b1111111111100001;
    assign weights1[26][749] = 16'b1111111111010010;
    assign weights1[26][750] = 16'b1111111111010101;
    assign weights1[26][751] = 16'b1111111111011100;
    assign weights1[26][752] = 16'b1111111111011101;
    assign weights1[26][753] = 16'b1111111111100101;
    assign weights1[26][754] = 16'b1111111111110000;
    assign weights1[26][755] = 16'b1111111111111000;
    assign weights1[26][756] = 16'b1111111111111111;
    assign weights1[26][757] = 16'b1111111111111110;
    assign weights1[26][758] = 16'b1111111111111001;
    assign weights1[26][759] = 16'b1111111111111101;
    assign weights1[26][760] = 16'b1111111111101111;
    assign weights1[26][761] = 16'b1111111111101000;
    assign weights1[26][762] = 16'b1111111111100110;
    assign weights1[26][763] = 16'b1111111111011011;
    assign weights1[26][764] = 16'b1111111111011100;
    assign weights1[26][765] = 16'b1111111111100001;
    assign weights1[26][766] = 16'b1111111111011010;
    assign weights1[26][767] = 16'b1111111111110000;
    assign weights1[26][768] = 16'b1111111111100011;
    assign weights1[26][769] = 16'b1111111111001100;
    assign weights1[26][770] = 16'b1111111111001111;
    assign weights1[26][771] = 16'b1111111111010010;
    assign weights1[26][772] = 16'b1111111111010111;
    assign weights1[26][773] = 16'b1111111111100100;
    assign weights1[26][774] = 16'b1111111111010101;
    assign weights1[26][775] = 16'b1111111111010000;
    assign weights1[26][776] = 16'b1111111111100000;
    assign weights1[26][777] = 16'b1111111111010001;
    assign weights1[26][778] = 16'b1111111111011101;
    assign weights1[26][779] = 16'b1111111111100110;
    assign weights1[26][780] = 16'b1111111111100111;
    assign weights1[26][781] = 16'b1111111111110001;
    assign weights1[26][782] = 16'b1111111111110111;
    assign weights1[26][783] = 16'b1111111111111101;
    assign weights1[27][0] = 16'b0000000000000000;
    assign weights1[27][1] = 16'b0000000000000000;
    assign weights1[27][2] = 16'b1111111111111101;
    assign weights1[27][3] = 16'b0000000000000000;
    assign weights1[27][4] = 16'b0000000000000001;
    assign weights1[27][5] = 16'b0000000000000000;
    assign weights1[27][6] = 16'b1111111111111110;
    assign weights1[27][7] = 16'b1111111111111011;
    assign weights1[27][8] = 16'b1111111111111010;
    assign weights1[27][9] = 16'b1111111111111100;
    assign weights1[27][10] = 16'b0000000000001000;
    assign weights1[27][11] = 16'b1111111111111011;
    assign weights1[27][12] = 16'b0000000000000110;
    assign weights1[27][13] = 16'b1111111111110110;
    assign weights1[27][14] = 16'b1111111111101011;
    assign weights1[27][15] = 16'b1111111111110110;
    assign weights1[27][16] = 16'b1111111111111011;
    assign weights1[27][17] = 16'b0000000000010010;
    assign weights1[27][18] = 16'b0000000000001001;
    assign weights1[27][19] = 16'b1111111111110111;
    assign weights1[27][20] = 16'b1111111111111000;
    assign weights1[27][21] = 16'b0000000000001001;
    assign weights1[27][22] = 16'b0000000000001100;
    assign weights1[27][23] = 16'b0000000000001010;
    assign weights1[27][24] = 16'b0000000000001111;
    assign weights1[27][25] = 16'b0000000000001001;
    assign weights1[27][26] = 16'b0000000000000001;
    assign weights1[27][27] = 16'b0000000000000010;
    assign weights1[27][28] = 16'b0000000000000001;
    assign weights1[27][29] = 16'b0000000000000000;
    assign weights1[27][30] = 16'b0000000000000001;
    assign weights1[27][31] = 16'b1111111111111110;
    assign weights1[27][32] = 16'b0000000000000011;
    assign weights1[27][33] = 16'b0000000000000011;
    assign weights1[27][34] = 16'b0000000000000001;
    assign weights1[27][35] = 16'b1111111111110100;
    assign weights1[27][36] = 16'b1111111111110011;
    assign weights1[27][37] = 16'b0000000000000110;
    assign weights1[27][38] = 16'b1111111111110011;
    assign weights1[27][39] = 16'b1111111111110001;
    assign weights1[27][40] = 16'b0000000000000000;
    assign weights1[27][41] = 16'b1111111111111100;
    assign weights1[27][42] = 16'b0000000000000001;
    assign weights1[27][43] = 16'b1111111111111110;
    assign weights1[27][44] = 16'b0000000000000011;
    assign weights1[27][45] = 16'b1111111111111111;
    assign weights1[27][46] = 16'b0000000000000011;
    assign weights1[27][47] = 16'b1111111111110111;
    assign weights1[27][48] = 16'b1111111111111011;
    assign weights1[27][49] = 16'b0000000000000010;
    assign weights1[27][50] = 16'b0000000000001100;
    assign weights1[27][51] = 16'b0000000000000011;
    assign weights1[27][52] = 16'b0000000000001000;
    assign weights1[27][53] = 16'b0000000000001010;
    assign weights1[27][54] = 16'b0000000000000001;
    assign weights1[27][55] = 16'b0000000000000100;
    assign weights1[27][56] = 16'b0000000000000000;
    assign weights1[27][57] = 16'b0000000000000010;
    assign weights1[27][58] = 16'b1111111111111110;
    assign weights1[27][59] = 16'b0000000000001010;
    assign weights1[27][60] = 16'b0000000000001011;
    assign weights1[27][61] = 16'b0000000000001111;
    assign weights1[27][62] = 16'b0000000000011101;
    assign weights1[27][63] = 16'b0000000000001001;
    assign weights1[27][64] = 16'b0000000000000001;
    assign weights1[27][65] = 16'b1111111111101101;
    assign weights1[27][66] = 16'b1111111111110101;
    assign weights1[27][67] = 16'b1111111111111001;
    assign weights1[27][68] = 16'b0000000000000011;
    assign weights1[27][69] = 16'b1111111111111001;
    assign weights1[27][70] = 16'b1111111111111100;
    assign weights1[27][71] = 16'b0000000000001100;
    assign weights1[27][72] = 16'b1111111111111000;
    assign weights1[27][73] = 16'b1111111111110110;
    assign weights1[27][74] = 16'b0000000000010000;
    assign weights1[27][75] = 16'b0000000000000110;
    assign weights1[27][76] = 16'b0000000000001101;
    assign weights1[27][77] = 16'b0000000000001100;
    assign weights1[27][78] = 16'b0000000000001000;
    assign weights1[27][79] = 16'b0000000000000111;
    assign weights1[27][80] = 16'b0000000000000011;
    assign weights1[27][81] = 16'b0000000000000110;
    assign weights1[27][82] = 16'b0000000000001011;
    assign weights1[27][83] = 16'b0000000000001000;
    assign weights1[27][84] = 16'b0000000000000010;
    assign weights1[27][85] = 16'b0000000000000011;
    assign weights1[27][86] = 16'b0000000000000111;
    assign weights1[27][87] = 16'b0000000000001111;
    assign weights1[27][88] = 16'b0000000000011111;
    assign weights1[27][89] = 16'b0000000000100111;
    assign weights1[27][90] = 16'b0000000000010111;
    assign weights1[27][91] = 16'b0000000000011011;
    assign weights1[27][92] = 16'b0000000000001000;
    assign weights1[27][93] = 16'b1111111111111111;
    assign weights1[27][94] = 16'b1111111111111100;
    assign weights1[27][95] = 16'b0000000000000011;
    assign weights1[27][96] = 16'b1111111111111100;
    assign weights1[27][97] = 16'b1111111111110011;
    assign weights1[27][98] = 16'b0000000000000010;
    assign weights1[27][99] = 16'b0000000000000111;
    assign weights1[27][100] = 16'b1111111111110101;
    assign weights1[27][101] = 16'b1111111111101111;
    assign weights1[27][102] = 16'b0000000000001011;
    assign weights1[27][103] = 16'b1111111111111010;
    assign weights1[27][104] = 16'b1111111111110101;
    assign weights1[27][105] = 16'b1111111111101000;
    assign weights1[27][106] = 16'b0000000000000001;
    assign weights1[27][107] = 16'b1111111111111110;
    assign weights1[27][108] = 16'b0000000000001011;
    assign weights1[27][109] = 16'b0000000000000001;
    assign weights1[27][110] = 16'b0000000000001010;
    assign weights1[27][111] = 16'b0000000000001010;
    assign weights1[27][112] = 16'b0000000000000001;
    assign weights1[27][113] = 16'b0000000000001000;
    assign weights1[27][114] = 16'b0000000000010001;
    assign weights1[27][115] = 16'b0000000000011101;
    assign weights1[27][116] = 16'b0000000000110010;
    assign weights1[27][117] = 16'b0000000000110011;
    assign weights1[27][118] = 16'b0000000000010101;
    assign weights1[27][119] = 16'b0000000000101100;
    assign weights1[27][120] = 16'b0000000000100111;
    assign weights1[27][121] = 16'b0000000000010000;
    assign weights1[27][122] = 16'b0000000000001010;
    assign weights1[27][123] = 16'b0000000000010100;
    assign weights1[27][124] = 16'b0000000000001101;
    assign weights1[27][125] = 16'b1111111111111101;
    assign weights1[27][126] = 16'b1111111111110101;
    assign weights1[27][127] = 16'b0000000000000001;
    assign weights1[27][128] = 16'b0000000000001110;
    assign weights1[27][129] = 16'b0000000000000010;
    assign weights1[27][130] = 16'b0000000000000001;
    assign weights1[27][131] = 16'b1111111111101000;
    assign weights1[27][132] = 16'b0000000000000011;
    assign weights1[27][133] = 16'b1111111111111101;
    assign weights1[27][134] = 16'b1111111111110001;
    assign weights1[27][135] = 16'b1111111111111100;
    assign weights1[27][136] = 16'b0000000000001010;
    assign weights1[27][137] = 16'b1111111111111000;
    assign weights1[27][138] = 16'b1111111111111101;
    assign weights1[27][139] = 16'b0000000000000001;
    assign weights1[27][140] = 16'b0000000000000101;
    assign weights1[27][141] = 16'b0000000000001111;
    assign weights1[27][142] = 16'b0000000000011011;
    assign weights1[27][143] = 16'b0000000000101001;
    assign weights1[27][144] = 16'b0000000000100010;
    assign weights1[27][145] = 16'b0000000000110011;
    assign weights1[27][146] = 16'b0000000000100000;
    assign weights1[27][147] = 16'b0000000000101000;
    assign weights1[27][148] = 16'b0000000000011001;
    assign weights1[27][149] = 16'b0000000000000110;
    assign weights1[27][150] = 16'b0000000000011011;
    assign weights1[27][151] = 16'b0000000000001000;
    assign weights1[27][152] = 16'b0000000000001001;
    assign weights1[27][153] = 16'b0000000000001000;
    assign weights1[27][154] = 16'b0000000000001100;
    assign weights1[27][155] = 16'b0000000000000101;
    assign weights1[27][156] = 16'b0000000000000100;
    assign weights1[27][157] = 16'b0000000000000100;
    assign weights1[27][158] = 16'b1111111111110011;
    assign weights1[27][159] = 16'b1111111111111110;
    assign weights1[27][160] = 16'b0000000000000111;
    assign weights1[27][161] = 16'b1111111111110001;
    assign weights1[27][162] = 16'b1111111111110101;
    assign weights1[27][163] = 16'b0000000000000010;
    assign weights1[27][164] = 16'b1111111111110110;
    assign weights1[27][165] = 16'b1111111111101111;
    assign weights1[27][166] = 16'b0000000000000000;
    assign weights1[27][167] = 16'b1111111111111101;
    assign weights1[27][168] = 16'b0000000000001011;
    assign weights1[27][169] = 16'b0000000000011100;
    assign weights1[27][170] = 16'b0000000000011000;
    assign weights1[27][171] = 16'b0000000000011111;
    assign weights1[27][172] = 16'b0000000000110000;
    assign weights1[27][173] = 16'b0000000000101110;
    assign weights1[27][174] = 16'b0000000000011110;
    assign weights1[27][175] = 16'b0000000000001011;
    assign weights1[27][176] = 16'b0000000000100111;
    assign weights1[27][177] = 16'b0000000000101101;
    assign weights1[27][178] = 16'b0000000000101100;
    assign weights1[27][179] = 16'b0000000000011100;
    assign weights1[27][180] = 16'b0000000000011110;
    assign weights1[27][181] = 16'b0000000000010011;
    assign weights1[27][182] = 16'b0000000000010010;
    assign weights1[27][183] = 16'b1111111111111011;
    assign weights1[27][184] = 16'b1111111111111100;
    assign weights1[27][185] = 16'b1111111111111101;
    assign weights1[27][186] = 16'b0000000000001001;
    assign weights1[27][187] = 16'b0000000000000110;
    assign weights1[27][188] = 16'b1111111111101101;
    assign weights1[27][189] = 16'b0000000000001001;
    assign weights1[27][190] = 16'b0000000000000010;
    assign weights1[27][191] = 16'b1111111111111110;
    assign weights1[27][192] = 16'b0000000000001000;
    assign weights1[27][193] = 16'b0000000000001101;
    assign weights1[27][194] = 16'b0000000000001010;
    assign weights1[27][195] = 16'b1111111111111000;
    assign weights1[27][196] = 16'b0000000000010011;
    assign weights1[27][197] = 16'b0000000000001111;
    assign weights1[27][198] = 16'b0000000000010000;
    assign weights1[27][199] = 16'b0000000000011010;
    assign weights1[27][200] = 16'b0000000000100100;
    assign weights1[27][201] = 16'b0000000000100011;
    assign weights1[27][202] = 16'b0000000000100110;
    assign weights1[27][203] = 16'b0000000000110010;
    assign weights1[27][204] = 16'b0000000000110011;
    assign weights1[27][205] = 16'b0000000000110000;
    assign weights1[27][206] = 16'b1111111111111100;
    assign weights1[27][207] = 16'b0000000000001111;
    assign weights1[27][208] = 16'b0000000000001001;
    assign weights1[27][209] = 16'b1111111111111001;
    assign weights1[27][210] = 16'b1111111111111101;
    assign weights1[27][211] = 16'b0000000000001011;
    assign weights1[27][212] = 16'b1111111111111010;
    assign weights1[27][213] = 16'b1111111111111011;
    assign weights1[27][214] = 16'b0000000000001111;
    assign weights1[27][215] = 16'b1111111111111011;
    assign weights1[27][216] = 16'b1111111111111101;
    assign weights1[27][217] = 16'b1111111111111000;
    assign weights1[27][218] = 16'b0000000000000011;
    assign weights1[27][219] = 16'b1111111111111100;
    assign weights1[27][220] = 16'b0000000000000010;
    assign weights1[27][221] = 16'b1111111111111001;
    assign weights1[27][222] = 16'b1111111111111000;
    assign weights1[27][223] = 16'b1111111111111110;
    assign weights1[27][224] = 16'b0000000000001110;
    assign weights1[27][225] = 16'b0000000000001001;
    assign weights1[27][226] = 16'b1111111111110000;
    assign weights1[27][227] = 16'b1111111111111011;
    assign weights1[27][228] = 16'b0000000000000011;
    assign weights1[27][229] = 16'b1111111111001111;
    assign weights1[27][230] = 16'b0000000000000111;
    assign weights1[27][231] = 16'b1111111111110110;
    assign weights1[27][232] = 16'b1111111111001111;
    assign weights1[27][233] = 16'b1111111111010011;
    assign weights1[27][234] = 16'b1111111111111111;
    assign weights1[27][235] = 16'b1111111111100001;
    assign weights1[27][236] = 16'b0000000000001010;
    assign weights1[27][237] = 16'b1111111111110011;
    assign weights1[27][238] = 16'b1111111111111011;
    assign weights1[27][239] = 16'b1111111111111000;
    assign weights1[27][240] = 16'b1111111111111001;
    assign weights1[27][241] = 16'b1111111111111000;
    assign weights1[27][242] = 16'b1111111111110001;
    assign weights1[27][243] = 16'b1111111111111001;
    assign weights1[27][244] = 16'b1111111111111111;
    assign weights1[27][245] = 16'b1111111111111111;
    assign weights1[27][246] = 16'b0000000000001000;
    assign weights1[27][247] = 16'b1111111111111101;
    assign weights1[27][248] = 16'b0000000000010011;
    assign weights1[27][249] = 16'b1111111111111011;
    assign weights1[27][250] = 16'b1111111111111110;
    assign weights1[27][251] = 16'b1111111111111110;
    assign weights1[27][252] = 16'b0000000000001001;
    assign weights1[27][253] = 16'b1111111111101010;
    assign weights1[27][254] = 16'b1111111111010010;
    assign weights1[27][255] = 16'b1111111111001110;
    assign weights1[27][256] = 16'b1111111111000111;
    assign weights1[27][257] = 16'b1111111110110010;
    assign weights1[27][258] = 16'b1111111110010101;
    assign weights1[27][259] = 16'b1111111110010111;
    assign weights1[27][260] = 16'b1111111110100101;
    assign weights1[27][261] = 16'b1111111110101001;
    assign weights1[27][262] = 16'b1111111111000100;
    assign weights1[27][263] = 16'b1111111111101100;
    assign weights1[27][264] = 16'b1111111111100111;
    assign weights1[27][265] = 16'b1111111111110100;
    assign weights1[27][266] = 16'b1111111111110001;
    assign weights1[27][267] = 16'b0000000000000100;
    assign weights1[27][268] = 16'b1111111111111101;
    assign weights1[27][269] = 16'b0000000000000110;
    assign weights1[27][270] = 16'b0000000000000000;
    assign weights1[27][271] = 16'b0000000000010011;
    assign weights1[27][272] = 16'b0000000000010010;
    assign weights1[27][273] = 16'b0000000000000101;
    assign weights1[27][274] = 16'b1111111111110110;
    assign weights1[27][275] = 16'b1111111111111010;
    assign weights1[27][276] = 16'b1111111111111011;
    assign weights1[27][277] = 16'b1111111111100101;
    assign weights1[27][278] = 16'b1111111111110100;
    assign weights1[27][279] = 16'b1111111111101011;
    assign weights1[27][280] = 16'b1111111111110010;
    assign weights1[27][281] = 16'b1111111111011011;
    assign weights1[27][282] = 16'b1111111111000010;
    assign weights1[27][283] = 16'b1111111110101111;
    assign weights1[27][284] = 16'b1111111110011000;
    assign weights1[27][285] = 16'b1111111110010100;
    assign weights1[27][286] = 16'b1111111110110010;
    assign weights1[27][287] = 16'b1111111111001010;
    assign weights1[27][288] = 16'b1111111111010010;
    assign weights1[27][289] = 16'b1111111111111110;
    assign weights1[27][290] = 16'b1111111111110010;
    assign weights1[27][291] = 16'b1111111111111000;
    assign weights1[27][292] = 16'b0000000000001010;
    assign weights1[27][293] = 16'b1111111111111100;
    assign weights1[27][294] = 16'b0000000000000101;
    assign weights1[27][295] = 16'b0000000000000001;
    assign weights1[27][296] = 16'b0000000000001101;
    assign weights1[27][297] = 16'b0000000000000110;
    assign weights1[27][298] = 16'b1111111111111011;
    assign weights1[27][299] = 16'b1111111111111111;
    assign weights1[27][300] = 16'b1111111111110000;
    assign weights1[27][301] = 16'b1111111111111011;
    assign weights1[27][302] = 16'b1111111111110101;
    assign weights1[27][303] = 16'b0000000000001100;
    assign weights1[27][304] = 16'b1111111111111010;
    assign weights1[27][305] = 16'b0000000000000010;
    assign weights1[27][306] = 16'b1111111111111111;
    assign weights1[27][307] = 16'b1111111111100111;
    assign weights1[27][308] = 16'b1111111111100111;
    assign weights1[27][309] = 16'b1111111111010111;
    assign weights1[27][310] = 16'b1111111111001110;
    assign weights1[27][311] = 16'b1111111111000000;
    assign weights1[27][312] = 16'b1111111111001101;
    assign weights1[27][313] = 16'b1111111111011100;
    assign weights1[27][314] = 16'b1111111111111011;
    assign weights1[27][315] = 16'b0000000000011000;
    assign weights1[27][316] = 16'b1111111111111011;
    assign weights1[27][317] = 16'b0000000000001100;
    assign weights1[27][318] = 16'b0000000000011000;
    assign weights1[27][319] = 16'b0000000000010010;
    assign weights1[27][320] = 16'b0000000000011101;
    assign weights1[27][321] = 16'b0000000000100010;
    assign weights1[27][322] = 16'b0000000000001011;
    assign weights1[27][323] = 16'b0000000000010101;
    assign weights1[27][324] = 16'b1111111111110000;
    assign weights1[27][325] = 16'b1111111111111011;
    assign weights1[27][326] = 16'b1111111111110100;
    assign weights1[27][327] = 16'b0000000000000001;
    assign weights1[27][328] = 16'b1111111111110011;
    assign weights1[27][329] = 16'b1111111111110100;
    assign weights1[27][330] = 16'b1111111111111100;
    assign weights1[27][331] = 16'b1111111111110000;
    assign weights1[27][332] = 16'b1111111111110100;
    assign weights1[27][333] = 16'b1111111111101010;
    assign weights1[27][334] = 16'b0000000000000010;
    assign weights1[27][335] = 16'b1111111111101000;
    assign weights1[27][336] = 16'b1111111111100100;
    assign weights1[27][337] = 16'b1111111111010010;
    assign weights1[27][338] = 16'b1111111111100101;
    assign weights1[27][339] = 16'b1111111111110101;
    assign weights1[27][340] = 16'b0000000000000100;
    assign weights1[27][341] = 16'b0000000000101010;
    assign weights1[27][342] = 16'b0000000000001001;
    assign weights1[27][343] = 16'b0000000000101100;
    assign weights1[27][344] = 16'b0000000000111100;
    assign weights1[27][345] = 16'b0000000000110000;
    assign weights1[27][346] = 16'b0000000000100100;
    assign weights1[27][347] = 16'b0000000000011011;
    assign weights1[27][348] = 16'b0000000000100011;
    assign weights1[27][349] = 16'b0000000000010101;
    assign weights1[27][350] = 16'b0000000000010010;
    assign weights1[27][351] = 16'b1111111111111000;
    assign weights1[27][352] = 16'b0000000000001010;
    assign weights1[27][353] = 16'b1111111111111001;
    assign weights1[27][354] = 16'b1111111111110010;
    assign weights1[27][355] = 16'b1111111111110001;
    assign weights1[27][356] = 16'b1111111111101111;
    assign weights1[27][357] = 16'b1111111111111100;
    assign weights1[27][358] = 16'b1111111111111000;
    assign weights1[27][359] = 16'b1111111111110000;
    assign weights1[27][360] = 16'b0000000000001100;
    assign weights1[27][361] = 16'b1111111111100111;
    assign weights1[27][362] = 16'b1111111111111000;
    assign weights1[27][363] = 16'b1111111111101011;
    assign weights1[27][364] = 16'b1111111111011100;
    assign weights1[27][365] = 16'b1111111111011001;
    assign weights1[27][366] = 16'b1111111111101100;
    assign weights1[27][367] = 16'b1111111111110110;
    assign weights1[27][368] = 16'b0000000000011101;
    assign weights1[27][369] = 16'b0000000000110110;
    assign weights1[27][370] = 16'b0000000000010100;
    assign weights1[27][371] = 16'b0000000000111011;
    assign weights1[27][372] = 16'b0000000000101010;
    assign weights1[27][373] = 16'b0000000000001001;
    assign weights1[27][374] = 16'b0000000000100100;
    assign weights1[27][375] = 16'b0000000000100010;
    assign weights1[27][376] = 16'b0000000000100000;
    assign weights1[27][377] = 16'b0000000000001100;
    assign weights1[27][378] = 16'b0000000000000101;
    assign weights1[27][379] = 16'b1111111111101010;
    assign weights1[27][380] = 16'b1111111111011011;
    assign weights1[27][381] = 16'b1111111111110111;
    assign weights1[27][382] = 16'b0000000000000000;
    assign weights1[27][383] = 16'b1111111111110110;
    assign weights1[27][384] = 16'b1111111111110101;
    assign weights1[27][385] = 16'b1111111111101111;
    assign weights1[27][386] = 16'b1111111111110001;
    assign weights1[27][387] = 16'b0000000000000101;
    assign weights1[27][388] = 16'b1111111111101100;
    assign weights1[27][389] = 16'b1111111111101001;
    assign weights1[27][390] = 16'b0000000000000000;
    assign weights1[27][391] = 16'b1111111111110001;
    assign weights1[27][392] = 16'b1111111111011011;
    assign weights1[27][393] = 16'b1111111111010101;
    assign weights1[27][394] = 16'b1111111111010011;
    assign weights1[27][395] = 16'b1111111111011111;
    assign weights1[27][396] = 16'b1111111111010111;
    assign weights1[27][397] = 16'b1111111111101110;
    assign weights1[27][398] = 16'b0000000000001101;
    assign weights1[27][399] = 16'b0000000000010100;
    assign weights1[27][400] = 16'b0000000000000001;
    assign weights1[27][401] = 16'b0000000000100100;
    assign weights1[27][402] = 16'b0000000000001101;
    assign weights1[27][403] = 16'b0000000000001100;
    assign weights1[27][404] = 16'b1111111111111000;
    assign weights1[27][405] = 16'b1111111111101110;
    assign weights1[27][406] = 16'b1111111111101000;
    assign weights1[27][407] = 16'b1111111111101110;
    assign weights1[27][408] = 16'b1111111111011111;
    assign weights1[27][409] = 16'b1111111111110101;
    assign weights1[27][410] = 16'b1111111111110011;
    assign weights1[27][411] = 16'b1111111111111010;
    assign weights1[27][412] = 16'b1111111111110101;
    assign weights1[27][413] = 16'b0000000000001101;
    assign weights1[27][414] = 16'b0000000000001101;
    assign weights1[27][415] = 16'b0000000000001001;
    assign weights1[27][416] = 16'b0000000000010000;
    assign weights1[27][417] = 16'b1111111111111101;
    assign weights1[27][418] = 16'b1111111111110001;
    assign weights1[27][419] = 16'b1111111111110010;
    assign weights1[27][420] = 16'b1111111111011100;
    assign weights1[27][421] = 16'b1111111110111011;
    assign weights1[27][422] = 16'b1111111110110110;
    assign weights1[27][423] = 16'b1111111110010100;
    assign weights1[27][424] = 16'b1111111110010000;
    assign weights1[27][425] = 16'b1111111101101110;
    assign weights1[27][426] = 16'b1111111110100010;
    assign weights1[27][427] = 16'b1111111111010011;
    assign weights1[27][428] = 16'b1111111111101111;
    assign weights1[27][429] = 16'b0000000000000110;
    assign weights1[27][430] = 16'b0000000000011100;
    assign weights1[27][431] = 16'b1111111111101001;
    assign weights1[27][432] = 16'b1111111111100100;
    assign weights1[27][433] = 16'b1111111111001110;
    assign weights1[27][434] = 16'b1111111111001011;
    assign weights1[27][435] = 16'b1111111111011010;
    assign weights1[27][436] = 16'b1111111111110010;
    assign weights1[27][437] = 16'b1111111111101010;
    assign weights1[27][438] = 16'b1111111111110000;
    assign weights1[27][439] = 16'b0000000000001010;
    assign weights1[27][440] = 16'b1111111111110100;
    assign weights1[27][441] = 16'b1111111111111000;
    assign weights1[27][442] = 16'b1111111111110111;
    assign weights1[27][443] = 16'b1111111111100110;
    assign weights1[27][444] = 16'b0000000000001011;
    assign weights1[27][445] = 16'b1111111111111110;
    assign weights1[27][446] = 16'b1111111111111100;
    assign weights1[27][447] = 16'b1111111111110111;
    assign weights1[27][448] = 16'b1111111111010000;
    assign weights1[27][449] = 16'b1111111110110111;
    assign weights1[27][450] = 16'b1111111110010110;
    assign weights1[27][451] = 16'b1111111101110010;
    assign weights1[27][452] = 16'b1111111101001101;
    assign weights1[27][453] = 16'b1111111100100101;
    assign weights1[27][454] = 16'b1111111100100001;
    assign weights1[27][455] = 16'b1111111100011100;
    assign weights1[27][456] = 16'b1111111100001101;
    assign weights1[27][457] = 16'b1111111101010111;
    assign weights1[27][458] = 16'b1111111101010101;
    assign weights1[27][459] = 16'b1111111101111101;
    assign weights1[27][460] = 16'b1111111110010101;
    assign weights1[27][461] = 16'b1111111110101011;
    assign weights1[27][462] = 16'b1111111111000110;
    assign weights1[27][463] = 16'b1111111111100111;
    assign weights1[27][464] = 16'b1111111111100111;
    assign weights1[27][465] = 16'b1111111111101010;
    assign weights1[27][466] = 16'b1111111111100110;
    assign weights1[27][467] = 16'b0000000000001001;
    assign weights1[27][468] = 16'b1111111111111101;
    assign weights1[27][469] = 16'b0000000000001010;
    assign weights1[27][470] = 16'b1111111111110100;
    assign weights1[27][471] = 16'b0000000000000001;
    assign weights1[27][472] = 16'b0000000000000010;
    assign weights1[27][473] = 16'b0000000000001001;
    assign weights1[27][474] = 16'b1111111111111100;
    assign weights1[27][475] = 16'b1111111111111001;
    assign weights1[27][476] = 16'b1111111111011100;
    assign weights1[27][477] = 16'b1111111110111000;
    assign weights1[27][478] = 16'b1111111110101011;
    assign weights1[27][479] = 16'b1111111110100111;
    assign weights1[27][480] = 16'b1111111101111101;
    assign weights1[27][481] = 16'b1111111101011111;
    assign weights1[27][482] = 16'b1111111101100100;
    assign weights1[27][483] = 16'b1111111100110000;
    assign weights1[27][484] = 16'b1111111100101100;
    assign weights1[27][485] = 16'b1111111100011111;
    assign weights1[27][486] = 16'b1111111101011110;
    assign weights1[27][487] = 16'b1111111110000100;
    assign weights1[27][488] = 16'b1111111110110010;
    assign weights1[27][489] = 16'b1111111111001110;
    assign weights1[27][490] = 16'b1111111111100101;
    assign weights1[27][491] = 16'b1111111111101010;
    assign weights1[27][492] = 16'b1111111111110100;
    assign weights1[27][493] = 16'b0000000000001001;
    assign weights1[27][494] = 16'b1111111111111010;
    assign weights1[27][495] = 16'b0000000000000110;
    assign weights1[27][496] = 16'b1111111111111000;
    assign weights1[27][497] = 16'b0000000000001011;
    assign weights1[27][498] = 16'b0000000000000110;
    assign weights1[27][499] = 16'b0000000000000100;
    assign weights1[27][500] = 16'b1111111111110100;
    assign weights1[27][501] = 16'b0000000000000011;
    assign weights1[27][502] = 16'b0000000000001001;
    assign weights1[27][503] = 16'b1111111111110111;
    assign weights1[27][504] = 16'b1111111111110011;
    assign weights1[27][505] = 16'b1111111111011001;
    assign weights1[27][506] = 16'b1111111111011111;
    assign weights1[27][507] = 16'b1111111111100110;
    assign weights1[27][508] = 16'b1111111111100000;
    assign weights1[27][509] = 16'b1111111111100000;
    assign weights1[27][510] = 16'b1111111111100010;
    assign weights1[27][511] = 16'b1111111111000101;
    assign weights1[27][512] = 16'b1111111111100100;
    assign weights1[27][513] = 16'b0000000000010001;
    assign weights1[27][514] = 16'b0000000000001111;
    assign weights1[27][515] = 16'b1111111111111111;
    assign weights1[27][516] = 16'b0000000000011001;
    assign weights1[27][517] = 16'b0000000000010001;
    assign weights1[27][518] = 16'b1111111111111111;
    assign weights1[27][519] = 16'b0000000000001100;
    assign weights1[27][520] = 16'b0000000000001100;
    assign weights1[27][521] = 16'b1111111111111110;
    assign weights1[27][522] = 16'b0000000000000111;
    assign weights1[27][523] = 16'b0000000000010010;
    assign weights1[27][524] = 16'b0000000000001110;
    assign weights1[27][525] = 16'b0000000000010111;
    assign weights1[27][526] = 16'b0000000000001100;
    assign weights1[27][527] = 16'b0000000000001111;
    assign weights1[27][528] = 16'b0000000000000100;
    assign weights1[27][529] = 16'b1111111111110111;
    assign weights1[27][530] = 16'b1111111111111011;
    assign weights1[27][531] = 16'b0000000000000101;
    assign weights1[27][532] = 16'b0000000000000010;
    assign weights1[27][533] = 16'b1111111111111010;
    assign weights1[27][534] = 16'b0000000000000011;
    assign weights1[27][535] = 16'b0000000000101000;
    assign weights1[27][536] = 16'b0000000000010100;
    assign weights1[27][537] = 16'b0000000000110101;
    assign weights1[27][538] = 16'b0000000000110101;
    assign weights1[27][539] = 16'b0000000001000111;
    assign weights1[27][540] = 16'b0000000001001110;
    assign weights1[27][541] = 16'b0000000000111111;
    assign weights1[27][542] = 16'b0000000000101010;
    assign weights1[27][543] = 16'b0000000000101011;
    assign weights1[27][544] = 16'b0000000000110001;
    assign weights1[27][545] = 16'b0000000000011011;
    assign weights1[27][546] = 16'b0000000000011001;
    assign weights1[27][547] = 16'b0000000000000010;
    assign weights1[27][548] = 16'b0000000000000011;
    assign weights1[27][549] = 16'b0000000000010101;
    assign weights1[27][550] = 16'b0000000000001100;
    assign weights1[27][551] = 16'b0000000000000010;
    assign weights1[27][552] = 16'b0000000000001010;
    assign weights1[27][553] = 16'b0000000000010000;
    assign weights1[27][554] = 16'b0000000000010000;
    assign weights1[27][555] = 16'b0000000000000100;
    assign weights1[27][556] = 16'b1111111111111111;
    assign weights1[27][557] = 16'b0000000000000111;
    assign weights1[27][558] = 16'b0000000000001001;
    assign weights1[27][559] = 16'b0000000000000101;
    assign weights1[27][560] = 16'b0000000000010010;
    assign weights1[27][561] = 16'b0000000000010100;
    assign weights1[27][562] = 16'b0000000000000111;
    assign weights1[27][563] = 16'b0000000001000101;
    assign weights1[27][564] = 16'b0000000001000011;
    assign weights1[27][565] = 16'b0000000000110101;
    assign weights1[27][566] = 16'b0000000000101101;
    assign weights1[27][567] = 16'b0000000000111011;
    assign weights1[27][568] = 16'b0000000001001000;
    assign weights1[27][569] = 16'b0000000000100101;
    assign weights1[27][570] = 16'b0000000000001101;
    assign weights1[27][571] = 16'b0000000000100000;
    assign weights1[27][572] = 16'b0000000000001111;
    assign weights1[27][573] = 16'b0000000000001010;
    assign weights1[27][574] = 16'b0000000000010100;
    assign weights1[27][575] = 16'b0000000000010011;
    assign weights1[27][576] = 16'b1111111111111101;
    assign weights1[27][577] = 16'b0000000000001101;
    assign weights1[27][578] = 16'b1111111111110001;
    assign weights1[27][579] = 16'b1111111111111100;
    assign weights1[27][580] = 16'b0000000000011001;
    assign weights1[27][581] = 16'b1111111111111010;
    assign weights1[27][582] = 16'b1111111111111110;
    assign weights1[27][583] = 16'b1111111111111110;
    assign weights1[27][584] = 16'b0000000000001000;
    assign weights1[27][585] = 16'b0000000000001110;
    assign weights1[27][586] = 16'b0000000000001101;
    assign weights1[27][587] = 16'b0000000000001110;
    assign weights1[27][588] = 16'b0000000000010100;
    assign weights1[27][589] = 16'b0000000000011011;
    assign weights1[27][590] = 16'b0000000000100011;
    assign weights1[27][591] = 16'b0000000000100011;
    assign weights1[27][592] = 16'b0000000000110001;
    assign weights1[27][593] = 16'b0000000000100010;
    assign weights1[27][594] = 16'b0000000000001111;
    assign weights1[27][595] = 16'b0000000000100110;
    assign weights1[27][596] = 16'b0000000000001001;
    assign weights1[27][597] = 16'b0000000000010010;
    assign weights1[27][598] = 16'b0000000000010001;
    assign weights1[27][599] = 16'b0000000000010001;
    assign weights1[27][600] = 16'b1111111111110100;
    assign weights1[27][601] = 16'b0000000000011100;
    assign weights1[27][602] = 16'b0000000000000011;
    assign weights1[27][603] = 16'b0000000000000011;
    assign weights1[27][604] = 16'b0000000000010001;
    assign weights1[27][605] = 16'b1111111111110111;
    assign weights1[27][606] = 16'b0000000000001111;
    assign weights1[27][607] = 16'b1111111111111100;
    assign weights1[27][608] = 16'b0000000000000101;
    assign weights1[27][609] = 16'b1111111111111010;
    assign weights1[27][610] = 16'b0000000000010111;
    assign weights1[27][611] = 16'b1111111111111111;
    assign weights1[27][612] = 16'b0000000000011101;
    assign weights1[27][613] = 16'b0000000000001101;
    assign weights1[27][614] = 16'b0000000000010110;
    assign weights1[27][615] = 16'b0000000000010100;
    assign weights1[27][616] = 16'b0000000000000110;
    assign weights1[27][617] = 16'b0000000000010000;
    assign weights1[27][618] = 16'b0000000000010010;
    assign weights1[27][619] = 16'b0000000000011011;
    assign weights1[27][620] = 16'b0000000000100011;
    assign weights1[27][621] = 16'b1111111111111101;
    assign weights1[27][622] = 16'b0000000000010011;
    assign weights1[27][623] = 16'b0000000000010101;
    assign weights1[27][624] = 16'b0000000000010111;
    assign weights1[27][625] = 16'b0000000000010101;
    assign weights1[27][626] = 16'b0000000000000101;
    assign weights1[27][627] = 16'b0000000000001010;
    assign weights1[27][628] = 16'b0000000000010111;
    assign weights1[27][629] = 16'b1111111111111101;
    assign weights1[27][630] = 16'b1111111111111100;
    assign weights1[27][631] = 16'b1111111111111110;
    assign weights1[27][632] = 16'b0000000000001100;
    assign weights1[27][633] = 16'b0000000000001101;
    assign weights1[27][634] = 16'b0000000000000000;
    assign weights1[27][635] = 16'b0000000000101010;
    assign weights1[27][636] = 16'b0000000000000111;
    assign weights1[27][637] = 16'b1111111111111000;
    assign weights1[27][638] = 16'b1111111111111110;
    assign weights1[27][639] = 16'b0000000000010011;
    assign weights1[27][640] = 16'b1111111111110010;
    assign weights1[27][641] = 16'b0000000000001010;
    assign weights1[27][642] = 16'b0000000000010100;
    assign weights1[27][643] = 16'b0000000000001101;
    assign weights1[27][644] = 16'b0000000000000101;
    assign weights1[27][645] = 16'b0000000000000111;
    assign weights1[27][646] = 16'b0000000000010010;
    assign weights1[27][647] = 16'b0000000000011000;
    assign weights1[27][648] = 16'b0000000000001011;
    assign weights1[27][649] = 16'b0000000000100101;
    assign weights1[27][650] = 16'b0000000000000101;
    assign weights1[27][651] = 16'b0000000000010111;
    assign weights1[27][652] = 16'b1111111111111101;
    assign weights1[27][653] = 16'b0000000000100100;
    assign weights1[27][654] = 16'b0000000000001000;
    assign weights1[27][655] = 16'b0000000000000111;
    assign weights1[27][656] = 16'b0000000000001011;
    assign weights1[27][657] = 16'b0000000000000110;
    assign weights1[27][658] = 16'b0000000000001100;
    assign weights1[27][659] = 16'b0000000000001100;
    assign weights1[27][660] = 16'b0000000000000100;
    assign weights1[27][661] = 16'b1111111111111101;
    assign weights1[27][662] = 16'b1111111111110110;
    assign weights1[27][663] = 16'b1111111111110101;
    assign weights1[27][664] = 16'b0000000000000001;
    assign weights1[27][665] = 16'b0000000000000011;
    assign weights1[27][666] = 16'b1111111111110111;
    assign weights1[27][667] = 16'b1111111111111111;
    assign weights1[27][668] = 16'b0000000000001000;
    assign weights1[27][669] = 16'b0000000000001110;
    assign weights1[27][670] = 16'b0000000000011010;
    assign weights1[27][671] = 16'b0000000000001111;
    assign weights1[27][672] = 16'b0000000000000011;
    assign weights1[27][673] = 16'b0000000000000010;
    assign weights1[27][674] = 16'b1111111111111101;
    assign weights1[27][675] = 16'b0000000000010011;
    assign weights1[27][676] = 16'b0000000000001010;
    assign weights1[27][677] = 16'b1111111111111101;
    assign weights1[27][678] = 16'b0000000000010111;
    assign weights1[27][679] = 16'b1111111111101010;
    assign weights1[27][680] = 16'b1111111111111010;
    assign weights1[27][681] = 16'b1111111111101111;
    assign weights1[27][682] = 16'b1111111111111000;
    assign weights1[27][683] = 16'b0000000000000011;
    assign weights1[27][684] = 16'b1111111111111010;
    assign weights1[27][685] = 16'b0000000000010000;
    assign weights1[27][686] = 16'b1111111111111000;
    assign weights1[27][687] = 16'b1111111111101011;
    assign weights1[27][688] = 16'b1111111111110100;
    assign weights1[27][689] = 16'b1111111111110001;
    assign weights1[27][690] = 16'b1111111111110110;
    assign weights1[27][691] = 16'b0000000000000110;
    assign weights1[27][692] = 16'b0000000000000101;
    assign weights1[27][693] = 16'b1111111111111001;
    assign weights1[27][694] = 16'b0000000000001101;
    assign weights1[27][695] = 16'b0000000000001110;
    assign weights1[27][696] = 16'b1111111111111101;
    assign weights1[27][697] = 16'b0000000000001001;
    assign weights1[27][698] = 16'b0000000000010110;
    assign weights1[27][699] = 16'b0000000000001000;
    assign weights1[27][700] = 16'b0000000000000100;
    assign weights1[27][701] = 16'b0000000000001010;
    assign weights1[27][702] = 16'b1111111111111100;
    assign weights1[27][703] = 16'b1111111111110110;
    assign weights1[27][704] = 16'b1111111111111011;
    assign weights1[27][705] = 16'b1111111111101110;
    assign weights1[27][706] = 16'b1111111111111000;
    assign weights1[27][707] = 16'b1111111111110110;
    assign weights1[27][708] = 16'b1111111111111010;
    assign weights1[27][709] = 16'b1111111111101001;
    assign weights1[27][710] = 16'b0000000000010010;
    assign weights1[27][711] = 16'b0000000000010011;
    assign weights1[27][712] = 16'b1111111111110111;
    assign weights1[27][713] = 16'b1111111111101011;
    assign weights1[27][714] = 16'b0000000000000101;
    assign weights1[27][715] = 16'b1111111111111101;
    assign weights1[27][716] = 16'b0000000000000011;
    assign weights1[27][717] = 16'b1111111111111110;
    assign weights1[27][718] = 16'b0000000000001110;
    assign weights1[27][719] = 16'b0000000000000011;
    assign weights1[27][720] = 16'b1111111111111101;
    assign weights1[27][721] = 16'b0000000000001010;
    assign weights1[27][722] = 16'b1111111111110100;
    assign weights1[27][723] = 16'b1111111111111000;
    assign weights1[27][724] = 16'b0000000000001011;
    assign weights1[27][725] = 16'b0000000000001000;
    assign weights1[27][726] = 16'b0000000000000000;
    assign weights1[27][727] = 16'b0000000000000111;
    assign weights1[27][728] = 16'b0000000000000111;
    assign weights1[27][729] = 16'b0000000000001001;
    assign weights1[27][730] = 16'b0000000000000011;
    assign weights1[27][731] = 16'b1111111111111010;
    assign weights1[27][732] = 16'b1111111111111000;
    assign weights1[27][733] = 16'b1111111111100101;
    assign weights1[27][734] = 16'b1111111111110100;
    assign weights1[27][735] = 16'b1111111111101001;
    assign weights1[27][736] = 16'b1111111111111100;
    assign weights1[27][737] = 16'b1111111111110011;
    assign weights1[27][738] = 16'b1111111111110000;
    assign weights1[27][739] = 16'b1111111111111101;
    assign weights1[27][740] = 16'b1111111111101101;
    assign weights1[27][741] = 16'b0000000000001100;
    assign weights1[27][742] = 16'b1111111111111110;
    assign weights1[27][743] = 16'b0000000000001001;
    assign weights1[27][744] = 16'b1111111111111110;
    assign weights1[27][745] = 16'b0000000000000110;
    assign weights1[27][746] = 16'b0000000000000111;
    assign weights1[27][747] = 16'b0000000000000110;
    assign weights1[27][748] = 16'b0000000000001010;
    assign weights1[27][749] = 16'b0000000000011000;
    assign weights1[27][750] = 16'b0000000000001111;
    assign weights1[27][751] = 16'b1111111111111001;
    assign weights1[27][752] = 16'b0000000000000101;
    assign weights1[27][753] = 16'b0000000000001000;
    assign weights1[27][754] = 16'b0000000000000100;
    assign weights1[27][755] = 16'b0000000000000001;
    assign weights1[27][756] = 16'b0000000000000010;
    assign weights1[27][757] = 16'b0000000000001010;
    assign weights1[27][758] = 16'b0000000000001011;
    assign weights1[27][759] = 16'b0000000000001000;
    assign weights1[27][760] = 16'b0000000000000111;
    assign weights1[27][761] = 16'b1111111111111111;
    assign weights1[27][762] = 16'b0000000000001101;
    assign weights1[27][763] = 16'b1111111111111111;
    assign weights1[27][764] = 16'b0000000000000110;
    assign weights1[27][765] = 16'b0000000000000100;
    assign weights1[27][766] = 16'b0000000000000111;
    assign weights1[27][767] = 16'b0000000000001110;
    assign weights1[27][768] = 16'b0000000000010010;
    assign weights1[27][769] = 16'b0000000000100011;
    assign weights1[27][770] = 16'b0000000000011001;
    assign weights1[27][771] = 16'b0000000000011000;
    assign weights1[27][772] = 16'b0000000000001101;
    assign weights1[27][773] = 16'b0000000000010100;
    assign weights1[27][774] = 16'b0000000000000011;
    assign weights1[27][775] = 16'b0000000000001101;
    assign weights1[27][776] = 16'b0000000000001110;
    assign weights1[27][777] = 16'b0000000000010001;
    assign weights1[27][778] = 16'b1111111111111110;
    assign weights1[27][779] = 16'b0000000000000000;
    assign weights1[27][780] = 16'b1111111111111001;
    assign weights1[27][781] = 16'b0000000000000011;
    assign weights1[27][782] = 16'b0000000000000101;
    assign weights1[27][783] = 16'b0000000000000000;
    assign weights1[28][0] = 16'b0000000000000000;
    assign weights1[28][1] = 16'b0000000000000000;
    assign weights1[28][2] = 16'b0000000000000000;
    assign weights1[28][3] = 16'b0000000000000000;
    assign weights1[28][4] = 16'b0000000000000000;
    assign weights1[28][5] = 16'b0000000000000000;
    assign weights1[28][6] = 16'b1111111111111011;
    assign weights1[28][7] = 16'b1111111111111100;
    assign weights1[28][8] = 16'b1111111111111010;
    assign weights1[28][9] = 16'b1111111111111010;
    assign weights1[28][10] = 16'b1111111111111100;
    assign weights1[28][11] = 16'b1111111111110101;
    assign weights1[28][12] = 16'b1111111111110000;
    assign weights1[28][13] = 16'b1111111111101111;
    assign weights1[28][14] = 16'b1111111111101100;
    assign weights1[28][15] = 16'b1111111111110101;
    assign weights1[28][16] = 16'b1111111111101000;
    assign weights1[28][17] = 16'b1111111111101010;
    assign weights1[28][18] = 16'b1111111111110110;
    assign weights1[28][19] = 16'b1111111111111010;
    assign weights1[28][20] = 16'b1111111111111001;
    assign weights1[28][21] = 16'b1111111111111000;
    assign weights1[28][22] = 16'b0000000000000000;
    assign weights1[28][23] = 16'b0000000000000011;
    assign weights1[28][24] = 16'b0000000000000100;
    assign weights1[28][25] = 16'b0000000000000110;
    assign weights1[28][26] = 16'b0000000000000001;
    assign weights1[28][27] = 16'b1111111111111111;
    assign weights1[28][28] = 16'b0000000000000000;
    assign weights1[28][29] = 16'b0000000000000000;
    assign weights1[28][30] = 16'b0000000000000001;
    assign weights1[28][31] = 16'b0000000000000001;
    assign weights1[28][32] = 16'b1111111111111100;
    assign weights1[28][33] = 16'b0000000000000010;
    assign weights1[28][34] = 16'b0000000000000000;
    assign weights1[28][35] = 16'b0000000000000001;
    assign weights1[28][36] = 16'b0000000000000000;
    assign weights1[28][37] = 16'b1111111111111111;
    assign weights1[28][38] = 16'b1111111111111011;
    assign weights1[28][39] = 16'b1111111111101111;
    assign weights1[28][40] = 16'b1111111111101100;
    assign weights1[28][41] = 16'b1111111111101100;
    assign weights1[28][42] = 16'b1111111111100011;
    assign weights1[28][43] = 16'b1111111111100110;
    assign weights1[28][44] = 16'b1111111111100100;
    assign weights1[28][45] = 16'b1111111111010101;
    assign weights1[28][46] = 16'b1111111111100101;
    assign weights1[28][47] = 16'b1111111111100011;
    assign weights1[28][48] = 16'b1111111111101001;
    assign weights1[28][49] = 16'b1111111111101111;
    assign weights1[28][50] = 16'b1111111111111000;
    assign weights1[28][51] = 16'b1111111111111010;
    assign weights1[28][52] = 16'b1111111111111100;
    assign weights1[28][53] = 16'b0000000000000000;
    assign weights1[28][54] = 16'b0000000000000011;
    assign weights1[28][55] = 16'b0000000000000011;
    assign weights1[28][56] = 16'b0000000000000000;
    assign weights1[28][57] = 16'b0000000000000000;
    assign weights1[28][58] = 16'b0000000000000000;
    assign weights1[28][59] = 16'b1111111111111101;
    assign weights1[28][60] = 16'b1111111111111011;
    assign weights1[28][61] = 16'b1111111111111101;
    assign weights1[28][62] = 16'b1111111111111011;
    assign weights1[28][63] = 16'b0000000000000100;
    assign weights1[28][64] = 16'b1111111111111111;
    assign weights1[28][65] = 16'b0000000000000001;
    assign weights1[28][66] = 16'b1111111111110101;
    assign weights1[28][67] = 16'b1111111111101101;
    assign weights1[28][68] = 16'b1111111111010010;
    assign weights1[28][69] = 16'b1111111111011011;
    assign weights1[28][70] = 16'b1111111111110011;
    assign weights1[28][71] = 16'b1111111111101001;
    assign weights1[28][72] = 16'b1111111111101010;
    assign weights1[28][73] = 16'b1111111111100011;
    assign weights1[28][74] = 16'b0000000000000011;
    assign weights1[28][75] = 16'b0000000000000010;
    assign weights1[28][76] = 16'b1111111111101100;
    assign weights1[28][77] = 16'b1111111111111111;
    assign weights1[28][78] = 16'b1111111111101100;
    assign weights1[28][79] = 16'b1111111111111100;
    assign weights1[28][80] = 16'b1111111111110100;
    assign weights1[28][81] = 16'b0000000000000110;
    assign weights1[28][82] = 16'b0000000000000011;
    assign weights1[28][83] = 16'b0000000000000101;
    assign weights1[28][84] = 16'b0000000000000000;
    assign weights1[28][85] = 16'b0000000000000000;
    assign weights1[28][86] = 16'b1111111111111101;
    assign weights1[28][87] = 16'b1111111111111101;
    assign weights1[28][88] = 16'b1111111111111010;
    assign weights1[28][89] = 16'b1111111111110111;
    assign weights1[28][90] = 16'b1111111111111101;
    assign weights1[28][91] = 16'b1111111111110111;
    assign weights1[28][92] = 16'b1111111111110001;
    assign weights1[28][93] = 16'b1111111111101011;
    assign weights1[28][94] = 16'b1111111111011000;
    assign weights1[28][95] = 16'b1111111111011110;
    assign weights1[28][96] = 16'b1111111111001011;
    assign weights1[28][97] = 16'b1111111111110010;
    assign weights1[28][98] = 16'b1111111111010101;
    assign weights1[28][99] = 16'b1111111111100010;
    assign weights1[28][100] = 16'b1111111111101111;
    assign weights1[28][101] = 16'b0000000000001001;
    assign weights1[28][102] = 16'b0000000000000110;
    assign weights1[28][103] = 16'b1111111111111110;
    assign weights1[28][104] = 16'b1111111111110100;
    assign weights1[28][105] = 16'b1111111111111110;
    assign weights1[28][106] = 16'b0000000000000110;
    assign weights1[28][107] = 16'b1111111111111110;
    assign weights1[28][108] = 16'b1111111111111000;
    assign weights1[28][109] = 16'b1111111111110011;
    assign weights1[28][110] = 16'b1111111111110101;
    assign weights1[28][111] = 16'b0000000000000001;
    assign weights1[28][112] = 16'b1111111111111110;
    assign weights1[28][113] = 16'b0000000000000000;
    assign weights1[28][114] = 16'b1111111111111110;
    assign weights1[28][115] = 16'b1111111111111101;
    assign weights1[28][116] = 16'b1111111111111101;
    assign weights1[28][117] = 16'b1111111111110100;
    assign weights1[28][118] = 16'b1111111111100000;
    assign weights1[28][119] = 16'b1111111111011111;
    assign weights1[28][120] = 16'b1111111111011111;
    assign weights1[28][121] = 16'b1111111111111011;
    assign weights1[28][122] = 16'b1111111111110111;
    assign weights1[28][123] = 16'b1111111111111101;
    assign weights1[28][124] = 16'b1111111111110000;
    assign weights1[28][125] = 16'b0000000000000100;
    assign weights1[28][126] = 16'b1111111111101110;
    assign weights1[28][127] = 16'b1111111111101000;
    assign weights1[28][128] = 16'b1111111111110110;
    assign weights1[28][129] = 16'b1111111111111001;
    assign weights1[28][130] = 16'b1111111111101111;
    assign weights1[28][131] = 16'b1111111111111000;
    assign weights1[28][132] = 16'b1111111111100010;
    assign weights1[28][133] = 16'b0000000000000111;
    assign weights1[28][134] = 16'b1111111111110000;
    assign weights1[28][135] = 16'b0000000000000000;
    assign weights1[28][136] = 16'b1111111111111000;
    assign weights1[28][137] = 16'b0000000000001010;
    assign weights1[28][138] = 16'b1111111111111001;
    assign weights1[28][139] = 16'b1111111111111100;
    assign weights1[28][140] = 16'b1111111111111110;
    assign weights1[28][141] = 16'b1111111111111100;
    assign weights1[28][142] = 16'b1111111111111100;
    assign weights1[28][143] = 16'b1111111111111000;
    assign weights1[28][144] = 16'b1111111111111111;
    assign weights1[28][145] = 16'b0000000000010010;
    assign weights1[28][146] = 16'b1111111111110110;
    assign weights1[28][147] = 16'b1111111111011011;
    assign weights1[28][148] = 16'b1111111111100111;
    assign weights1[28][149] = 16'b0000000000000110;
    assign weights1[28][150] = 16'b1111111111110001;
    assign weights1[28][151] = 16'b0000000000001001;
    assign weights1[28][152] = 16'b1111111111110001;
    assign weights1[28][153] = 16'b1111111111101011;
    assign weights1[28][154] = 16'b1111111111111000;
    assign weights1[28][155] = 16'b0000000000000011;
    assign weights1[28][156] = 16'b0000000000000010;
    assign weights1[28][157] = 16'b0000000000001100;
    assign weights1[28][158] = 16'b1111111111101111;
    assign weights1[28][159] = 16'b0000000000001010;
    assign weights1[28][160] = 16'b0000000000000001;
    assign weights1[28][161] = 16'b1111111111111110;
    assign weights1[28][162] = 16'b1111111111111111;
    assign weights1[28][163] = 16'b1111111111111010;
    assign weights1[28][164] = 16'b0000000000000110;
    assign weights1[28][165] = 16'b0000000000000011;
    assign weights1[28][166] = 16'b0000000000001001;
    assign weights1[28][167] = 16'b0000000000000011;
    assign weights1[28][168] = 16'b1111111111111100;
    assign weights1[28][169] = 16'b1111111111110110;
    assign weights1[28][170] = 16'b1111111111101111;
    assign weights1[28][171] = 16'b1111111111110111;
    assign weights1[28][172] = 16'b0000000000000000;
    assign weights1[28][173] = 16'b0000000000001101;
    assign weights1[28][174] = 16'b1111111111110110;
    assign weights1[28][175] = 16'b1111111111101101;
    assign weights1[28][176] = 16'b1111111111100011;
    assign weights1[28][177] = 16'b1111111111100100;
    assign weights1[28][178] = 16'b1111111111110111;
    assign weights1[28][179] = 16'b0000000000000001;
    assign weights1[28][180] = 16'b0000000000000101;
    assign weights1[28][181] = 16'b1111111111110011;
    assign weights1[28][182] = 16'b0000000000000000;
    assign weights1[28][183] = 16'b1111111111110111;
    assign weights1[28][184] = 16'b1111111111111110;
    assign weights1[28][185] = 16'b0000000000000111;
    assign weights1[28][186] = 16'b0000000000001101;
    assign weights1[28][187] = 16'b0000000000010000;
    assign weights1[28][188] = 16'b0000000000011100;
    assign weights1[28][189] = 16'b0000000000001110;
    assign weights1[28][190] = 16'b0000000000000111;
    assign weights1[28][191] = 16'b0000000000000100;
    assign weights1[28][192] = 16'b0000000000101111;
    assign weights1[28][193] = 16'b0000000000010111;
    assign weights1[28][194] = 16'b0000000000010101;
    assign weights1[28][195] = 16'b0000000000010001;
    assign weights1[28][196] = 16'b1111111111111100;
    assign weights1[28][197] = 16'b1111111111110111;
    assign weights1[28][198] = 16'b1111111111101111;
    assign weights1[28][199] = 16'b1111111111110110;
    assign weights1[28][200] = 16'b1111111111111001;
    assign weights1[28][201] = 16'b1111111111100011;
    assign weights1[28][202] = 16'b0000000000000011;
    assign weights1[28][203] = 16'b1111111111101101;
    assign weights1[28][204] = 16'b1111111111111100;
    assign weights1[28][205] = 16'b1111111111111011;
    assign weights1[28][206] = 16'b1111111111110110;
    assign weights1[28][207] = 16'b1111111111111000;
    assign weights1[28][208] = 16'b1111111111111110;
    assign weights1[28][209] = 16'b0000000000010000;
    assign weights1[28][210] = 16'b1111111111110010;
    assign weights1[28][211] = 16'b0000000000001000;
    assign weights1[28][212] = 16'b1111111111110100;
    assign weights1[28][213] = 16'b0000000000001110;
    assign weights1[28][214] = 16'b0000000000000010;
    assign weights1[28][215] = 16'b1111111111110011;
    assign weights1[28][216] = 16'b0000000000001101;
    assign weights1[28][217] = 16'b0000000000100101;
    assign weights1[28][218] = 16'b0000000000101110;
    assign weights1[28][219] = 16'b0000000000011011;
    assign weights1[28][220] = 16'b1111111111111100;
    assign weights1[28][221] = 16'b0000000000011001;
    assign weights1[28][222] = 16'b0000000000011000;
    assign weights1[28][223] = 16'b0000000000011110;
    assign weights1[28][224] = 16'b1111111111111010;
    assign weights1[28][225] = 16'b1111111111110101;
    assign weights1[28][226] = 16'b1111111111110101;
    assign weights1[28][227] = 16'b1111111111111000;
    assign weights1[28][228] = 16'b1111111111110010;
    assign weights1[28][229] = 16'b1111111111101011;
    assign weights1[28][230] = 16'b0000000000000001;
    assign weights1[28][231] = 16'b1111111111011101;
    assign weights1[28][232] = 16'b0000000000000010;
    assign weights1[28][233] = 16'b1111111111110001;
    assign weights1[28][234] = 16'b0000000000001001;
    assign weights1[28][235] = 16'b1111111111111110;
    assign weights1[28][236] = 16'b1111111111111001;
    assign weights1[28][237] = 16'b1111111111110101;
    assign weights1[28][238] = 16'b0000000000001000;
    assign weights1[28][239] = 16'b0000000000010101;
    assign weights1[28][240] = 16'b0000000000011011;
    assign weights1[28][241] = 16'b0000000000000001;
    assign weights1[28][242] = 16'b0000000000010010;
    assign weights1[28][243] = 16'b0000000000000100;
    assign weights1[28][244] = 16'b0000000000010010;
    assign weights1[28][245] = 16'b0000000000011110;
    assign weights1[28][246] = 16'b0000000000010111;
    assign weights1[28][247] = 16'b0000000000010110;
    assign weights1[28][248] = 16'b0000000000110110;
    assign weights1[28][249] = 16'b0000000000101010;
    assign weights1[28][250] = 16'b0000000000011110;
    assign weights1[28][251] = 16'b0000000000110101;
    assign weights1[28][252] = 16'b1111111111110101;
    assign weights1[28][253] = 16'b1111111111111101;
    assign weights1[28][254] = 16'b1111111111111001;
    assign weights1[28][255] = 16'b1111111111110100;
    assign weights1[28][256] = 16'b1111111111111111;
    assign weights1[28][257] = 16'b1111111111110101;
    assign weights1[28][258] = 16'b1111111111101110;
    assign weights1[28][259] = 16'b1111111111011111;
    assign weights1[28][260] = 16'b0000000000000011;
    assign weights1[28][261] = 16'b1111111111110010;
    assign weights1[28][262] = 16'b1111111111101110;
    assign weights1[28][263] = 16'b1111111111111010;
    assign weights1[28][264] = 16'b1111111111111111;
    assign weights1[28][265] = 16'b0000000000001000;
    assign weights1[28][266] = 16'b0000000000000101;
    assign weights1[28][267] = 16'b0000000000010100;
    assign weights1[28][268] = 16'b0000000000010000;
    assign weights1[28][269] = 16'b0000000000100010;
    assign weights1[28][270] = 16'b0000000000100110;
    assign weights1[28][271] = 16'b0000000000111001;
    assign weights1[28][272] = 16'b0000000000101100;
    assign weights1[28][273] = 16'b0000000000100100;
    assign weights1[28][274] = 16'b0000000000101110;
    assign weights1[28][275] = 16'b0000000000111000;
    assign weights1[28][276] = 16'b0000000001000001;
    assign weights1[28][277] = 16'b0000000000110101;
    assign weights1[28][278] = 16'b0000000000000101;
    assign weights1[28][279] = 16'b0000000000101100;
    assign weights1[28][280] = 16'b1111111111110010;
    assign weights1[28][281] = 16'b1111111111111100;
    assign weights1[28][282] = 16'b0000000000010101;
    assign weights1[28][283] = 16'b1111111111110100;
    assign weights1[28][284] = 16'b1111111111100110;
    assign weights1[28][285] = 16'b1111111111101110;
    assign weights1[28][286] = 16'b1111111111111000;
    assign weights1[28][287] = 16'b1111111111110101;
    assign weights1[28][288] = 16'b1111111111110101;
    assign weights1[28][289] = 16'b1111111111101000;
    assign weights1[28][290] = 16'b0000000000000000;
    assign weights1[28][291] = 16'b1111111111110100;
    assign weights1[28][292] = 16'b1111111111111000;
    assign weights1[28][293] = 16'b0000000000001000;
    assign weights1[28][294] = 16'b1111111111110110;
    assign weights1[28][295] = 16'b1111111111111011;
    assign weights1[28][296] = 16'b0000000000010010;
    assign weights1[28][297] = 16'b0000000000011100;
    assign weights1[28][298] = 16'b0000000000100111;
    assign weights1[28][299] = 16'b0000000000011000;
    assign weights1[28][300] = 16'b0000000000110011;
    assign weights1[28][301] = 16'b0000000000110000;
    assign weights1[28][302] = 16'b0000000000111000;
    assign weights1[28][303] = 16'b0000000001001111;
    assign weights1[28][304] = 16'b0000000000100110;
    assign weights1[28][305] = 16'b0000000001000011;
    assign weights1[28][306] = 16'b0000000000001101;
    assign weights1[28][307] = 16'b1111111111111100;
    assign weights1[28][308] = 16'b1111111111110001;
    assign weights1[28][309] = 16'b1111111111110000;
    assign weights1[28][310] = 16'b0000000000000011;
    assign weights1[28][311] = 16'b1111111111101110;
    assign weights1[28][312] = 16'b1111111111111110;
    assign weights1[28][313] = 16'b1111111111110111;
    assign weights1[28][314] = 16'b1111111111110011;
    assign weights1[28][315] = 16'b0000000000000101;
    assign weights1[28][316] = 16'b1111111111110110;
    assign weights1[28][317] = 16'b0000000000000111;
    assign weights1[28][318] = 16'b1111111111110100;
    assign weights1[28][319] = 16'b1111111111100111;
    assign weights1[28][320] = 16'b1111111111110100;
    assign weights1[28][321] = 16'b1111111111011100;
    assign weights1[28][322] = 16'b1111111111010001;
    assign weights1[28][323] = 16'b1111111111000011;
    assign weights1[28][324] = 16'b1111111110110111;
    assign weights1[28][325] = 16'b1111111111001100;
    assign weights1[28][326] = 16'b1111111111001001;
    assign weights1[28][327] = 16'b1111111111100001;
    assign weights1[28][328] = 16'b1111111111100110;
    assign weights1[28][329] = 16'b0000000000011111;
    assign weights1[28][330] = 16'b0000000000010100;
    assign weights1[28][331] = 16'b0000000000000010;
    assign weights1[28][332] = 16'b1111111111110110;
    assign weights1[28][333] = 16'b1111111111111100;
    assign weights1[28][334] = 16'b1111111111101001;
    assign weights1[28][335] = 16'b1111111111101100;
    assign weights1[28][336] = 16'b1111111111111100;
    assign weights1[28][337] = 16'b1111111111110001;
    assign weights1[28][338] = 16'b0000000000001000;
    assign weights1[28][339] = 16'b1111111111111101;
    assign weights1[28][340] = 16'b1111111111110001;
    assign weights1[28][341] = 16'b0000000000000010;
    assign weights1[28][342] = 16'b1111111111111101;
    assign weights1[28][343] = 16'b1111111111101010;
    assign weights1[28][344] = 16'b1111111111111001;
    assign weights1[28][345] = 16'b1111111111100000;
    assign weights1[28][346] = 16'b1111111111111000;
    assign weights1[28][347] = 16'b1111111111101110;
    assign weights1[28][348] = 16'b1111111111011100;
    assign weights1[28][349] = 16'b1111111111101100;
    assign weights1[28][350] = 16'b1111111111010001;
    assign weights1[28][351] = 16'b1111111110111101;
    assign weights1[28][352] = 16'b1111111101110101;
    assign weights1[28][353] = 16'b1111111101000110;
    assign weights1[28][354] = 16'b1111111100011110;
    assign weights1[28][355] = 16'b1111111100100010;
    assign weights1[28][356] = 16'b1111111100010110;
    assign weights1[28][357] = 16'b1111111101000010;
    assign weights1[28][358] = 16'b1111111101010010;
    assign weights1[28][359] = 16'b1111111101100001;
    assign weights1[28][360] = 16'b1111111110001110;
    assign weights1[28][361] = 16'b1111111110011010;
    assign weights1[28][362] = 16'b1111111110101111;
    assign weights1[28][363] = 16'b1111111110110010;
    assign weights1[28][364] = 16'b0000000000001000;
    assign weights1[28][365] = 16'b1111111111111010;
    assign weights1[28][366] = 16'b0000000000010000;
    assign weights1[28][367] = 16'b0000000000001101;
    assign weights1[28][368] = 16'b1111111111111101;
    assign weights1[28][369] = 16'b1111111111111110;
    assign weights1[28][370] = 16'b1111111111110000;
    assign weights1[28][371] = 16'b1111111111110111;
    assign weights1[28][372] = 16'b0000000000000100;
    assign weights1[28][373] = 16'b1111111111110010;
    assign weights1[28][374] = 16'b1111111111101101;
    assign weights1[28][375] = 16'b1111111111111010;
    assign weights1[28][376] = 16'b0000000000001111;
    assign weights1[28][377] = 16'b1111111111111100;
    assign weights1[28][378] = 16'b1111111111111101;
    assign weights1[28][379] = 16'b1111111111101011;
    assign weights1[28][380] = 16'b1111111111101011;
    assign weights1[28][381] = 16'b1111111111001111;
    assign weights1[28][382] = 16'b1111111110001001;
    assign weights1[28][383] = 16'b1111111100010000;
    assign weights1[28][384] = 16'b1111111100001111;
    assign weights1[28][385] = 16'b1111111100011001;
    assign weights1[28][386] = 16'b1111111100111000;
    assign weights1[28][387] = 16'b1111111101000000;
    assign weights1[28][388] = 16'b1111111101011101;
    assign weights1[28][389] = 16'b1111111110000100;
    assign weights1[28][390] = 16'b1111111110101100;
    assign weights1[28][391] = 16'b1111111110110001;
    assign weights1[28][392] = 16'b0000000000000101;
    assign weights1[28][393] = 16'b1111111111111110;
    assign weights1[28][394] = 16'b1111111111111111;
    assign weights1[28][395] = 16'b0000000000010001;
    assign weights1[28][396] = 16'b0000000000010010;
    assign weights1[28][397] = 16'b1111111111111001;
    assign weights1[28][398] = 16'b0000000000001000;
    assign weights1[28][399] = 16'b1111111111110101;
    assign weights1[28][400] = 16'b0000000000000011;
    assign weights1[28][401] = 16'b0000000000001100;
    assign weights1[28][402] = 16'b0000000000000010;
    assign weights1[28][403] = 16'b1111111111111110;
    assign weights1[28][404] = 16'b1111111111110011;
    assign weights1[28][405] = 16'b1111111111110101;
    assign weights1[28][406] = 16'b0000000000010010;
    assign weights1[28][407] = 16'b0000000000001010;
    assign weights1[28][408] = 16'b0000000000011101;
    assign weights1[28][409] = 16'b0000000000000111;
    assign weights1[28][410] = 16'b0000000000001010;
    assign weights1[28][411] = 16'b1111111111011111;
    assign weights1[28][412] = 16'b1111111110100110;
    assign weights1[28][413] = 16'b1111111101010111;
    assign weights1[28][414] = 16'b1111111101010010;
    assign weights1[28][415] = 16'b1111111101100101;
    assign weights1[28][416] = 16'b1111111101110100;
    assign weights1[28][417] = 16'b1111111110001101;
    assign weights1[28][418] = 16'b1111111110101001;
    assign weights1[28][419] = 16'b1111111110101000;
    assign weights1[28][420] = 16'b0000000000000101;
    assign weights1[28][421] = 16'b0000000000000011;
    assign weights1[28][422] = 16'b0000000000001001;
    assign weights1[28][423] = 16'b0000000000000010;
    assign weights1[28][424] = 16'b1111111111111001;
    assign weights1[28][425] = 16'b0000000000001011;
    assign weights1[28][426] = 16'b0000000000010111;
    assign weights1[28][427] = 16'b1111111111111110;
    assign weights1[28][428] = 16'b0000000000001011;
    assign weights1[28][429] = 16'b0000000000001010;
    assign weights1[28][430] = 16'b1111111111110100;
    assign weights1[28][431] = 16'b0000000000000001;
    assign weights1[28][432] = 16'b1111111111111011;
    assign weights1[28][433] = 16'b1111111111111001;
    assign weights1[28][434] = 16'b1111111111111111;
    assign weights1[28][435] = 16'b0000000000000001;
    assign weights1[28][436] = 16'b0000000000000100;
    assign weights1[28][437] = 16'b0000000000011110;
    assign weights1[28][438] = 16'b0000000000101100;
    assign weights1[28][439] = 16'b0000000000001000;
    assign weights1[28][440] = 16'b0000000000010010;
    assign weights1[28][441] = 16'b1111111111011111;
    assign weights1[28][442] = 16'b1111111110101000;
    assign weights1[28][443] = 16'b1111111110010101;
    assign weights1[28][444] = 16'b1111111101110010;
    assign weights1[28][445] = 16'b1111111110011001;
    assign weights1[28][446] = 16'b1111111110111100;
    assign weights1[28][447] = 16'b1111111110011101;
    assign weights1[28][448] = 16'b0000000000010000;
    assign weights1[28][449] = 16'b0000000000010110;
    assign weights1[28][450] = 16'b1111111111101111;
    assign weights1[28][451] = 16'b1111111111111001;
    assign weights1[28][452] = 16'b1111111111110111;
    assign weights1[28][453] = 16'b0000000000010000;
    assign weights1[28][454] = 16'b1111111111111111;
    assign weights1[28][455] = 16'b0000000000001001;
    assign weights1[28][456] = 16'b1111111111111011;
    assign weights1[28][457] = 16'b0000000000001100;
    assign weights1[28][458] = 16'b1111111111110111;
    assign weights1[28][459] = 16'b0000000000000000;
    assign weights1[28][460] = 16'b0000000000001000;
    assign weights1[28][461] = 16'b1111111111111011;
    assign weights1[28][462] = 16'b1111111111110110;
    assign weights1[28][463] = 16'b1111111111111101;
    assign weights1[28][464] = 16'b0000000000010000;
    assign weights1[28][465] = 16'b0000000000000010;
    assign weights1[28][466] = 16'b0000000000001100;
    assign weights1[28][467] = 16'b0000000000001111;
    assign weights1[28][468] = 16'b0000000000010100;
    assign weights1[28][469] = 16'b0000000000011100;
    assign weights1[28][470] = 16'b0000000000011110;
    assign weights1[28][471] = 16'b1111111111101011;
    assign weights1[28][472] = 16'b1111111110110100;
    assign weights1[28][473] = 16'b1111111110100111;
    assign weights1[28][474] = 16'b1111111110111110;
    assign weights1[28][475] = 16'b1111111110111011;
    assign weights1[28][476] = 16'b0000000000001101;
    assign weights1[28][477] = 16'b0000000000000101;
    assign weights1[28][478] = 16'b1111111111101111;
    assign weights1[28][479] = 16'b1111111111111000;
    assign weights1[28][480] = 16'b0000000000001001;
    assign weights1[28][481] = 16'b0000000000000100;
    assign weights1[28][482] = 16'b0000000000000001;
    assign weights1[28][483] = 16'b0000000000010001;
    assign weights1[28][484] = 16'b1111111111111110;
    assign weights1[28][485] = 16'b1111111111111000;
    assign weights1[28][486] = 16'b0000000000000111;
    assign weights1[28][487] = 16'b1111111111101001;
    assign weights1[28][488] = 16'b1111111111111111;
    assign weights1[28][489] = 16'b1111111111111100;
    assign weights1[28][490] = 16'b1111111111111101;
    assign weights1[28][491] = 16'b0000000000001101;
    assign weights1[28][492] = 16'b0000000000000111;
    assign weights1[28][493] = 16'b0000000000001010;
    assign weights1[28][494] = 16'b0000000000001000;
    assign weights1[28][495] = 16'b0000000000010111;
    assign weights1[28][496] = 16'b0000000000011110;
    assign weights1[28][497] = 16'b1111111111111000;
    assign weights1[28][498] = 16'b0000000000011100;
    assign weights1[28][499] = 16'b0000000000011011;
    assign weights1[28][500] = 16'b1111111111110110;
    assign weights1[28][501] = 16'b1111111111100111;
    assign weights1[28][502] = 16'b1111111111001110;
    assign weights1[28][503] = 16'b1111111111001010;
    assign weights1[28][504] = 16'b0000000000000001;
    assign weights1[28][505] = 16'b0000000000000101;
    assign weights1[28][506] = 16'b0000000000001100;
    assign weights1[28][507] = 16'b0000000000000110;
    assign weights1[28][508] = 16'b0000000000000010;
    assign weights1[28][509] = 16'b0000000000000101;
    assign weights1[28][510] = 16'b1111111111111111;
    assign weights1[28][511] = 16'b0000000000001111;
    assign weights1[28][512] = 16'b0000000000000000;
    assign weights1[28][513] = 16'b1111111111111011;
    assign weights1[28][514] = 16'b0000000000000111;
    assign weights1[28][515] = 16'b0000000000000011;
    assign weights1[28][516] = 16'b0000000000000000;
    assign weights1[28][517] = 16'b1111111111111001;
    assign weights1[28][518] = 16'b0000000000001000;
    assign weights1[28][519] = 16'b1111111111111110;
    assign weights1[28][520] = 16'b0000000000001100;
    assign weights1[28][521] = 16'b0000000000001000;
    assign weights1[28][522] = 16'b0000000000010011;
    assign weights1[28][523] = 16'b1111111111111111;
    assign weights1[28][524] = 16'b0000000000011110;
    assign weights1[28][525] = 16'b1111111111111110;
    assign weights1[28][526] = 16'b0000000000001000;
    assign weights1[28][527] = 16'b0000000000001000;
    assign weights1[28][528] = 16'b1111111111110101;
    assign weights1[28][529] = 16'b1111111111101001;
    assign weights1[28][530] = 16'b1111111111011011;
    assign weights1[28][531] = 16'b1111111111010001;
    assign weights1[28][532] = 16'b1111111111111101;
    assign weights1[28][533] = 16'b0000000000001010;
    assign weights1[28][534] = 16'b1111111111111111;
    assign weights1[28][535] = 16'b0000000000001001;
    assign weights1[28][536] = 16'b1111111111110100;
    assign weights1[28][537] = 16'b1111111111111011;
    assign weights1[28][538] = 16'b0000000000000111;
    assign weights1[28][539] = 16'b0000000000001111;
    assign weights1[28][540] = 16'b0000000000000101;
    assign weights1[28][541] = 16'b0000000000000011;
    assign weights1[28][542] = 16'b1111111111110101;
    assign weights1[28][543] = 16'b0000000000001110;
    assign weights1[28][544] = 16'b0000000000000011;
    assign weights1[28][545] = 16'b1111111111111100;
    assign weights1[28][546] = 16'b0000000000000001;
    assign weights1[28][547] = 16'b0000000000001011;
    assign weights1[28][548] = 16'b0000000000001100;
    assign weights1[28][549] = 16'b0000000000000101;
    assign weights1[28][550] = 16'b0000000000000010;
    assign weights1[28][551] = 16'b0000000000000101;
    assign weights1[28][552] = 16'b0000000000010110;
    assign weights1[28][553] = 16'b0000000000000101;
    assign weights1[28][554] = 16'b0000000000100000;
    assign weights1[28][555] = 16'b0000000000011000;
    assign weights1[28][556] = 16'b0000000000001110;
    assign weights1[28][557] = 16'b1111111111110100;
    assign weights1[28][558] = 16'b1111111111100101;
    assign weights1[28][559] = 16'b1111111111011111;
    assign weights1[28][560] = 16'b1111111111111010;
    assign weights1[28][561] = 16'b1111111111111001;
    assign weights1[28][562] = 16'b0000000000010010;
    assign weights1[28][563] = 16'b1111111111111101;
    assign weights1[28][564] = 16'b1111111111111110;
    assign weights1[28][565] = 16'b0000000000001010;
    assign weights1[28][566] = 16'b0000000000000000;
    assign weights1[28][567] = 16'b1111111111110111;
    assign weights1[28][568] = 16'b0000000000001010;
    assign weights1[28][569] = 16'b1111111111111000;
    assign weights1[28][570] = 16'b0000000000000110;
    assign weights1[28][571] = 16'b0000000000000101;
    assign weights1[28][572] = 16'b0000000000000101;
    assign weights1[28][573] = 16'b1111111111111010;
    assign weights1[28][574] = 16'b0000000000000100;
    assign weights1[28][575] = 16'b0000000000000110;
    assign weights1[28][576] = 16'b0000000000000101;
    assign weights1[28][577] = 16'b1111111111111011;
    assign weights1[28][578] = 16'b0000000000011101;
    assign weights1[28][579] = 16'b1111111111110110;
    assign weights1[28][580] = 16'b0000000000011000;
    assign weights1[28][581] = 16'b0000000000000111;
    assign weights1[28][582] = 16'b0000000000000001;
    assign weights1[28][583] = 16'b0000000000010010;
    assign weights1[28][584] = 16'b0000000000000100;
    assign weights1[28][585] = 16'b0000000000000111;
    assign weights1[28][586] = 16'b1111111111111001;
    assign weights1[28][587] = 16'b1111111111101101;
    assign weights1[28][588] = 16'b0000000000000010;
    assign weights1[28][589] = 16'b1111111111110100;
    assign weights1[28][590] = 16'b0000000000001000;
    assign weights1[28][591] = 16'b0000000000000010;
    assign weights1[28][592] = 16'b1111111111111001;
    assign weights1[28][593] = 16'b1111111111111001;
    assign weights1[28][594] = 16'b1111111111101000;
    assign weights1[28][595] = 16'b0000000000000111;
    assign weights1[28][596] = 16'b0000000000001010;
    assign weights1[28][597] = 16'b0000000000000100;
    assign weights1[28][598] = 16'b0000000000001100;
    assign weights1[28][599] = 16'b1111111111110100;
    assign weights1[28][600] = 16'b0000000000010010;
    assign weights1[28][601] = 16'b0000000000000111;
    assign weights1[28][602] = 16'b0000000000001010;
    assign weights1[28][603] = 16'b0000000000000101;
    assign weights1[28][604] = 16'b0000000000001001;
    assign weights1[28][605] = 16'b0000000000001100;
    assign weights1[28][606] = 16'b0000000000001110;
    assign weights1[28][607] = 16'b0000000000000110;
    assign weights1[28][608] = 16'b0000000000001110;
    assign weights1[28][609] = 16'b0000000000010011;
    assign weights1[28][610] = 16'b0000000000001110;
    assign weights1[28][611] = 16'b0000000000001110;
    assign weights1[28][612] = 16'b0000000000000001;
    assign weights1[28][613] = 16'b0000000000010000;
    assign weights1[28][614] = 16'b0000000000000111;
    assign weights1[28][615] = 16'b1111111111111001;
    assign weights1[28][616] = 16'b1111111111111100;
    assign weights1[28][617] = 16'b0000000000000110;
    assign weights1[28][618] = 16'b0000000000001101;
    assign weights1[28][619] = 16'b0000000000000101;
    assign weights1[28][620] = 16'b1111111111110110;
    assign weights1[28][621] = 16'b0000000000000001;
    assign weights1[28][622] = 16'b1111111111111010;
    assign weights1[28][623] = 16'b1111111111111001;
    assign weights1[28][624] = 16'b1111111111101010;
    assign weights1[28][625] = 16'b0000000000010001;
    assign weights1[28][626] = 16'b0000000000000001;
    assign weights1[28][627] = 16'b0000000000001100;
    assign weights1[28][628] = 16'b0000000000010001;
    assign weights1[28][629] = 16'b0000000000000101;
    assign weights1[28][630] = 16'b0000000000001000;
    assign weights1[28][631] = 16'b0000000000010010;
    assign weights1[28][632] = 16'b0000000000001011;
    assign weights1[28][633] = 16'b0000000000001010;
    assign weights1[28][634] = 16'b0000000000010010;
    assign weights1[28][635] = 16'b1111111111111010;
    assign weights1[28][636] = 16'b0000000000010100;
    assign weights1[28][637] = 16'b0000000000011001;
    assign weights1[28][638] = 16'b0000000000000110;
    assign weights1[28][639] = 16'b0000000000000100;
    assign weights1[28][640] = 16'b0000000000100100;
    assign weights1[28][641] = 16'b0000000000010100;
    assign weights1[28][642] = 16'b0000000000001100;
    assign weights1[28][643] = 16'b0000000000000010;
    assign weights1[28][644] = 16'b0000000000000000;
    assign weights1[28][645] = 16'b0000000000001100;
    assign weights1[28][646] = 16'b0000000000000101;
    assign weights1[28][647] = 16'b0000000000001101;
    assign weights1[28][648] = 16'b0000000000000011;
    assign weights1[28][649] = 16'b1111111111111111;
    assign weights1[28][650] = 16'b0000000000010001;
    assign weights1[28][651] = 16'b1111111111111100;
    assign weights1[28][652] = 16'b1111111111111001;
    assign weights1[28][653] = 16'b1111111111111001;
    assign weights1[28][654] = 16'b0000000000000110;
    assign weights1[28][655] = 16'b0000000000000110;
    assign weights1[28][656] = 16'b1111111111111111;
    assign weights1[28][657] = 16'b1111111111111111;
    assign weights1[28][658] = 16'b0000000000001000;
    assign weights1[28][659] = 16'b1111111111111101;
    assign weights1[28][660] = 16'b0000000000000001;
    assign weights1[28][661] = 16'b1111111111110111;
    assign weights1[28][662] = 16'b0000000000001001;
    assign weights1[28][663] = 16'b1111111111110010;
    assign weights1[28][664] = 16'b0000000000001101;
    assign weights1[28][665] = 16'b0000000000010001;
    assign weights1[28][666] = 16'b0000000000000111;
    assign weights1[28][667] = 16'b0000000000010110;
    assign weights1[28][668] = 16'b0000000000100100;
    assign weights1[28][669] = 16'b0000000000011101;
    assign weights1[28][670] = 16'b0000000000011011;
    assign weights1[28][671] = 16'b0000000000000001;
    assign weights1[28][672] = 16'b0000000000000000;
    assign weights1[28][673] = 16'b0000000000000010;
    assign weights1[28][674] = 16'b0000000000001110;
    assign weights1[28][675] = 16'b1111111111111101;
    assign weights1[28][676] = 16'b1111111111111000;
    assign weights1[28][677] = 16'b0000000000000010;
    assign weights1[28][678] = 16'b0000000000000011;
    assign weights1[28][679] = 16'b0000000000000100;
    assign weights1[28][680] = 16'b0000000000001000;
    assign weights1[28][681] = 16'b0000000000001000;
    assign weights1[28][682] = 16'b0000000000000100;
    assign weights1[28][683] = 16'b1111111111111101;
    assign weights1[28][684] = 16'b0000000000000011;
    assign weights1[28][685] = 16'b0000000000000100;
    assign weights1[28][686] = 16'b0000000000000000;
    assign weights1[28][687] = 16'b0000000000010001;
    assign weights1[28][688] = 16'b0000000000000101;
    assign weights1[28][689] = 16'b0000000000011010;
    assign weights1[28][690] = 16'b0000000000001101;
    assign weights1[28][691] = 16'b0000000000000001;
    assign weights1[28][692] = 16'b0000000000000101;
    assign weights1[28][693] = 16'b0000000000010011;
    assign weights1[28][694] = 16'b1111111111111110;
    assign weights1[28][695] = 16'b1111111111110100;
    assign weights1[28][696] = 16'b0000000000001011;
    assign weights1[28][697] = 16'b1111111111110111;
    assign weights1[28][698] = 16'b0000000000000011;
    assign weights1[28][699] = 16'b1111111111111111;
    assign weights1[28][700] = 16'b0000000000000000;
    assign weights1[28][701] = 16'b0000000000000110;
    assign weights1[28][702] = 16'b1111111111111100;
    assign weights1[28][703] = 16'b0000000000000011;
    assign weights1[28][704] = 16'b0000000000000100;
    assign weights1[28][705] = 16'b0000000000000000;
    assign weights1[28][706] = 16'b0000000000000010;
    assign weights1[28][707] = 16'b0000000000000110;
    assign weights1[28][708] = 16'b0000000000010101;
    assign weights1[28][709] = 16'b1111111111111011;
    assign weights1[28][710] = 16'b0000000000010001;
    assign weights1[28][711] = 16'b0000000000000001;
    assign weights1[28][712] = 16'b0000000000011001;
    assign weights1[28][713] = 16'b0000000000001000;
    assign weights1[28][714] = 16'b0000000000001001;
    assign weights1[28][715] = 16'b1111111111110111;
    assign weights1[28][716] = 16'b1111111111111001;
    assign weights1[28][717] = 16'b0000000000000000;
    assign weights1[28][718] = 16'b1111111111111101;
    assign weights1[28][719] = 16'b0000000000000001;
    assign weights1[28][720] = 16'b0000000000010000;
    assign weights1[28][721] = 16'b0000000000001100;
    assign weights1[28][722] = 16'b1111111111111111;
    assign weights1[28][723] = 16'b0000000000000010;
    assign weights1[28][724] = 16'b0000000000010011;
    assign weights1[28][725] = 16'b0000000000000011;
    assign weights1[28][726] = 16'b0000000000000010;
    assign weights1[28][727] = 16'b1111111111111100;
    assign weights1[28][728] = 16'b1111111111111111;
    assign weights1[28][729] = 16'b1111111111110110;
    assign weights1[28][730] = 16'b1111111111110110;
    assign weights1[28][731] = 16'b0000000000000011;
    assign weights1[28][732] = 16'b0000000000001001;
    assign weights1[28][733] = 16'b1111111111111111;
    assign weights1[28][734] = 16'b0000000000000001;
    assign weights1[28][735] = 16'b0000000000000001;
    assign weights1[28][736] = 16'b0000000000000001;
    assign weights1[28][737] = 16'b0000000000000000;
    assign weights1[28][738] = 16'b1111111111110011;
    assign weights1[28][739] = 16'b1111111111111111;
    assign weights1[28][740] = 16'b0000000000000001;
    assign weights1[28][741] = 16'b0000000000000100;
    assign weights1[28][742] = 16'b1111111111110101;
    assign weights1[28][743] = 16'b0000000000000110;
    assign weights1[28][744] = 16'b0000000000010011;
    assign weights1[28][745] = 16'b0000000000000100;
    assign weights1[28][746] = 16'b0000000000010011;
    assign weights1[28][747] = 16'b1111111111111010;
    assign weights1[28][748] = 16'b0000000000001010;
    assign weights1[28][749] = 16'b0000000000010111;
    assign weights1[28][750] = 16'b1111111111111000;
    assign weights1[28][751] = 16'b0000000000000100;
    assign weights1[28][752] = 16'b0000000000001110;
    assign weights1[28][753] = 16'b0000000000001001;
    assign weights1[28][754] = 16'b0000000000000010;
    assign weights1[28][755] = 16'b0000000000000000;
    assign weights1[28][756] = 16'b1111111111111110;
    assign weights1[28][757] = 16'b1111111111111100;
    assign weights1[28][758] = 16'b1111111111111101;
    assign weights1[28][759] = 16'b1111111111110111;
    assign weights1[28][760] = 16'b1111111111111000;
    assign weights1[28][761] = 16'b0000000000001100;
    assign weights1[28][762] = 16'b0000000000001001;
    assign weights1[28][763] = 16'b0000000000001100;
    assign weights1[28][764] = 16'b0000000000001000;
    assign weights1[28][765] = 16'b0000000000001110;
    assign weights1[28][766] = 16'b0000000000001010;
    assign weights1[28][767] = 16'b0000000000010111;
    assign weights1[28][768] = 16'b0000000000010001;
    assign weights1[28][769] = 16'b0000000000000000;
    assign weights1[28][770] = 16'b0000000000011000;
    assign weights1[28][771] = 16'b0000000000001010;
    assign weights1[28][772] = 16'b1111111111111000;
    assign weights1[28][773] = 16'b0000000000000000;
    assign weights1[28][774] = 16'b0000000000010010;
    assign weights1[28][775] = 16'b0000000000000111;
    assign weights1[28][776] = 16'b0000000000011010;
    assign weights1[28][777] = 16'b0000000000010000;
    assign weights1[28][778] = 16'b0000000000000110;
    assign weights1[28][779] = 16'b0000000000000100;
    assign weights1[28][780] = 16'b0000000000000101;
    assign weights1[28][781] = 16'b0000000000001001;
    assign weights1[28][782] = 16'b1111111111111111;
    assign weights1[28][783] = 16'b1111111111111111;
    assign weights1[29][0] = 16'b0000000000000000;
    assign weights1[29][1] = 16'b0000000000000000;
    assign weights1[29][2] = 16'b1111111111111110;
    assign weights1[29][3] = 16'b1111111111110011;
    assign weights1[29][4] = 16'b1111111111101011;
    assign weights1[29][5] = 16'b1111111111100011;
    assign weights1[29][6] = 16'b1111111111110000;
    assign weights1[29][7] = 16'b0000000000000001;
    assign weights1[29][8] = 16'b0000000000011001;
    assign weights1[29][9] = 16'b0000000000111011;
    assign weights1[29][10] = 16'b0000000001010000;
    assign weights1[29][11] = 16'b0000000001010111;
    assign weights1[29][12] = 16'b0000000001000101;
    assign weights1[29][13] = 16'b0000000000101000;
    assign weights1[29][14] = 16'b0000000000100010;
    assign weights1[29][15] = 16'b0000000000010001;
    assign weights1[29][16] = 16'b0000000000001100;
    assign weights1[29][17] = 16'b1111111111110011;
    assign weights1[29][18] = 16'b1111111111101010;
    assign weights1[29][19] = 16'b1111111111101110;
    assign weights1[29][20] = 16'b1111111111100101;
    assign weights1[29][21] = 16'b1111111111100111;
    assign weights1[29][22] = 16'b1111111111101100;
    assign weights1[29][23] = 16'b1111111111111110;
    assign weights1[29][24] = 16'b1111111111111011;
    assign weights1[29][25] = 16'b0000000000000001;
    assign weights1[29][26] = 16'b0000000000000010;
    assign weights1[29][27] = 16'b0000000000000001;
    assign weights1[29][28] = 16'b0000000000000000;
    assign weights1[29][29] = 16'b1111111111111110;
    assign weights1[29][30] = 16'b1111111111110111;
    assign weights1[29][31] = 16'b1111111111100111;
    assign weights1[29][32] = 16'b1111111111011110;
    assign weights1[29][33] = 16'b1111111111011101;
    assign weights1[29][34] = 16'b1111111111100011;
    assign weights1[29][35] = 16'b0000000000001110;
    assign weights1[29][36] = 16'b0000000000010110;
    assign weights1[29][37] = 16'b0000000000110010;
    assign weights1[29][38] = 16'b0000000001000101;
    assign weights1[29][39] = 16'b0000000000111110;
    assign weights1[29][40] = 16'b0000000000100111;
    assign weights1[29][41] = 16'b0000000000010010;
    assign weights1[29][42] = 16'b1111111111111010;
    assign weights1[29][43] = 16'b1111111111111110;
    assign weights1[29][44] = 16'b1111111111111111;
    assign weights1[29][45] = 16'b1111111111101001;
    assign weights1[29][46] = 16'b1111111111010010;
    assign weights1[29][47] = 16'b1111111111000100;
    assign weights1[29][48] = 16'b1111111110111111;
    assign weights1[29][49] = 16'b1111111111011001;
    assign weights1[29][50] = 16'b1111111111100011;
    assign weights1[29][51] = 16'b1111111111110010;
    assign weights1[29][52] = 16'b1111111111111001;
    assign weights1[29][53] = 16'b0000000000000100;
    assign weights1[29][54] = 16'b0000000000001010;
    assign weights1[29][55] = 16'b0000000000000000;
    assign weights1[29][56] = 16'b1111111111111100;
    assign weights1[29][57] = 16'b1111111111111000;
    assign weights1[29][58] = 16'b1111111111110000;
    assign weights1[29][59] = 16'b1111111111011101;
    assign weights1[29][60] = 16'b1111111111001011;
    assign weights1[29][61] = 16'b1111111111001111;
    assign weights1[29][62] = 16'b1111111111101110;
    assign weights1[29][63] = 16'b0000000000101111;
    assign weights1[29][64] = 16'b0000000000111010;
    assign weights1[29][65] = 16'b0000000001001010;
    assign weights1[29][66] = 16'b0000000000101110;
    assign weights1[29][67] = 16'b0000000000011111;
    assign weights1[29][68] = 16'b0000000000101110;
    assign weights1[29][69] = 16'b0000000000011101;
    assign weights1[29][70] = 16'b0000000000000111;
    assign weights1[29][71] = 16'b1111111111110011;
    assign weights1[29][72] = 16'b1111111111011100;
    assign weights1[29][73] = 16'b1111111110111001;
    assign weights1[29][74] = 16'b1111111110100011;
    assign weights1[29][75] = 16'b1111111110011110;
    assign weights1[29][76] = 16'b1111111110101100;
    assign weights1[29][77] = 16'b1111111111010101;
    assign weights1[29][78] = 16'b1111111111101100;
    assign weights1[29][79] = 16'b1111111111111010;
    assign weights1[29][80] = 16'b1111111111111010;
    assign weights1[29][81] = 16'b0000000000000001;
    assign weights1[29][82] = 16'b0000000000000110;
    assign weights1[29][83] = 16'b1111111111111101;
    assign weights1[29][84] = 16'b1111111111110110;
    assign weights1[29][85] = 16'b1111111111101111;
    assign weights1[29][86] = 16'b1111111111011110;
    assign weights1[29][87] = 16'b1111111111000111;
    assign weights1[29][88] = 16'b1111111111000001;
    assign weights1[29][89] = 16'b1111111111011110;
    assign weights1[29][90] = 16'b1111111111110101;
    assign weights1[29][91] = 16'b0000000000011111;
    assign weights1[29][92] = 16'b0000000000111110;
    assign weights1[29][93] = 16'b0000000001001001;
    assign weights1[29][94] = 16'b0000000000110011;
    assign weights1[29][95] = 16'b0000000000101101;
    assign weights1[29][96] = 16'b0000000000100110;
    assign weights1[29][97] = 16'b0000000000000111;
    assign weights1[29][98] = 16'b1111111111100101;
    assign weights1[29][99] = 16'b1111111111000001;
    assign weights1[29][100] = 16'b1111111110010111;
    assign weights1[29][101] = 16'b1111111101110110;
    assign weights1[29][102] = 16'b1111111110000100;
    assign weights1[29][103] = 16'b1111111110011001;
    assign weights1[29][104] = 16'b1111111111000010;
    assign weights1[29][105] = 16'b1111111111100101;
    assign weights1[29][106] = 16'b0000000000000010;
    assign weights1[29][107] = 16'b0000000000000010;
    assign weights1[29][108] = 16'b1111111111111101;
    assign weights1[29][109] = 16'b0000000000000100;
    assign weights1[29][110] = 16'b0000000000001110;
    assign weights1[29][111] = 16'b0000000000001000;
    assign weights1[29][112] = 16'b1111111111110101;
    assign weights1[29][113] = 16'b1111111111100111;
    assign weights1[29][114] = 16'b1111111111010100;
    assign weights1[29][115] = 16'b1111111110111010;
    assign weights1[29][116] = 16'b1111111111001100;
    assign weights1[29][117] = 16'b1111111111111100;
    assign weights1[29][118] = 16'b0000000000000011;
    assign weights1[29][119] = 16'b0000000000110100;
    assign weights1[29][120] = 16'b0000000001000111;
    assign weights1[29][121] = 16'b0000000000111001;
    assign weights1[29][122] = 16'b0000000000100101;
    assign weights1[29][123] = 16'b0000000000110101;
    assign weights1[29][124] = 16'b0000000000001001;
    assign weights1[29][125] = 16'b1111111111011110;
    assign weights1[29][126] = 16'b1111111110100100;
    assign weights1[29][127] = 16'b1111111101111110;
    assign weights1[29][128] = 16'b1111111101010111;
    assign weights1[29][129] = 16'b1111111101100010;
    assign weights1[29][130] = 16'b1111111110000111;
    assign weights1[29][131] = 16'b1111111111000111;
    assign weights1[29][132] = 16'b1111111111101000;
    assign weights1[29][133] = 16'b1111111111101010;
    assign weights1[29][134] = 16'b1111111111111111;
    assign weights1[29][135] = 16'b1111111111111111;
    assign weights1[29][136] = 16'b1111111111111011;
    assign weights1[29][137] = 16'b1111111111111010;
    assign weights1[29][138] = 16'b1111111111111110;
    assign weights1[29][139] = 16'b0000000000001001;
    assign weights1[29][140] = 16'b1111111111110100;
    assign weights1[29][141] = 16'b1111111111100110;
    assign weights1[29][142] = 16'b1111111111001100;
    assign weights1[29][143] = 16'b1111111110111110;
    assign weights1[29][144] = 16'b1111111111100000;
    assign weights1[29][145] = 16'b0000000000001100;
    assign weights1[29][146] = 16'b0000000000001010;
    assign weights1[29][147] = 16'b0000000000011001;
    assign weights1[29][148] = 16'b0000000000001000;
    assign weights1[29][149] = 16'b0000000000100000;
    assign weights1[29][150] = 16'b0000000000111110;
    assign weights1[29][151] = 16'b0000000000011100;
    assign weights1[29][152] = 16'b1111111111001100;
    assign weights1[29][153] = 16'b1111111110010011;
    assign weights1[29][154] = 16'b1111111110001010;
    assign weights1[29][155] = 16'b1111111101100010;
    assign weights1[29][156] = 16'b1111111110001000;
    assign weights1[29][157] = 16'b1111111111000111;
    assign weights1[29][158] = 16'b1111111111010100;
    assign weights1[29][159] = 16'b1111111111101111;
    assign weights1[29][160] = 16'b1111111111111111;
    assign weights1[29][161] = 16'b0000000000000101;
    assign weights1[29][162] = 16'b1111111111111100;
    assign weights1[29][163] = 16'b1111111111100111;
    assign weights1[29][164] = 16'b1111111111111000;
    assign weights1[29][165] = 16'b0000000000000001;
    assign weights1[29][166] = 16'b0000000000011100;
    assign weights1[29][167] = 16'b0000000000010001;
    assign weights1[29][168] = 16'b1111111111110110;
    assign weights1[29][169] = 16'b1111111111100000;
    assign weights1[29][170] = 16'b1111111111001010;
    assign weights1[29][171] = 16'b1111111111000011;
    assign weights1[29][172] = 16'b1111111111110010;
    assign weights1[29][173] = 16'b0000000000010010;
    assign weights1[29][174] = 16'b0000000000011000;
    assign weights1[29][175] = 16'b0000000000001100;
    assign weights1[29][176] = 16'b0000000000010100;
    assign weights1[29][177] = 16'b0000000000110111;
    assign weights1[29][178] = 16'b0000000000111011;
    assign weights1[29][179] = 16'b0000000000000111;
    assign weights1[29][180] = 16'b1111111110101000;
    assign weights1[29][181] = 16'b1111111110010000;
    assign weights1[29][182] = 16'b1111111101110001;
    assign weights1[29][183] = 16'b1111111101111011;
    assign weights1[29][184] = 16'b1111111110101011;
    assign weights1[29][185] = 16'b1111111111101111;
    assign weights1[29][186] = 16'b1111111111111000;
    assign weights1[29][187] = 16'b0000000000000111;
    assign weights1[29][188] = 16'b0000000000000111;
    assign weights1[29][189] = 16'b0000000000001101;
    assign weights1[29][190] = 16'b1111111111110111;
    assign weights1[29][191] = 16'b0000000000010101;
    assign weights1[29][192] = 16'b1111111111111011;
    assign weights1[29][193] = 16'b0000000000001101;
    assign weights1[29][194] = 16'b0000000000010101;
    assign weights1[29][195] = 16'b0000000000010000;
    assign weights1[29][196] = 16'b1111111111101110;
    assign weights1[29][197] = 16'b1111111111011100;
    assign weights1[29][198] = 16'b1111111111001001;
    assign weights1[29][199] = 16'b1111111111010110;
    assign weights1[29][200] = 16'b1111111111110111;
    assign weights1[29][201] = 16'b0000000000011100;
    assign weights1[29][202] = 16'b0000000000010110;
    assign weights1[29][203] = 16'b0000000000101100;
    assign weights1[29][204] = 16'b0000000000010011;
    assign weights1[29][205] = 16'b0000000000010110;
    assign weights1[29][206] = 16'b0000000000100111;
    assign weights1[29][207] = 16'b1111111111101011;
    assign weights1[29][208] = 16'b1111111101111011;
    assign weights1[29][209] = 16'b1111111110001001;
    assign weights1[29][210] = 16'b1111111110100111;
    assign weights1[29][211] = 16'b1111111110111000;
    assign weights1[29][212] = 16'b1111111111101110;
    assign weights1[29][213] = 16'b1111111111111010;
    assign weights1[29][214] = 16'b1111111111010011;
    assign weights1[29][215] = 16'b0000000000000010;
    assign weights1[29][216] = 16'b0000000000010000;
    assign weights1[29][217] = 16'b0000000000011110;
    assign weights1[29][218] = 16'b1111111111111101;
    assign weights1[29][219] = 16'b0000000000010111;
    assign weights1[29][220] = 16'b0000000000000110;
    assign weights1[29][221] = 16'b1111111111111101;
    assign weights1[29][222] = 16'b0000000000010000;
    assign weights1[29][223] = 16'b0000000000001110;
    assign weights1[29][224] = 16'b1111111111110100;
    assign weights1[29][225] = 16'b1111111111100010;
    assign weights1[29][226] = 16'b1111111111011001;
    assign weights1[29][227] = 16'b1111111111010100;
    assign weights1[29][228] = 16'b1111111111111100;
    assign weights1[29][229] = 16'b0000000000010001;
    assign weights1[29][230] = 16'b0000000000000000;
    assign weights1[29][231] = 16'b0000000000011110;
    assign weights1[29][232] = 16'b0000000000010111;
    assign weights1[29][233] = 16'b0000000000100001;
    assign weights1[29][234] = 16'b0000000000110001;
    assign weights1[29][235] = 16'b1111111111010000;
    assign weights1[29][236] = 16'b1111111110010000;
    assign weights1[29][237] = 16'b1111111111000010;
    assign weights1[29][238] = 16'b1111111111000100;
    assign weights1[29][239] = 16'b1111111111100100;
    assign weights1[29][240] = 16'b1111111111110111;
    assign weights1[29][241] = 16'b0000000000011011;
    assign weights1[29][242] = 16'b0000000000011011;
    assign weights1[29][243] = 16'b0000000000011101;
    assign weights1[29][244] = 16'b0000000000001010;
    assign weights1[29][245] = 16'b0000000000011001;
    assign weights1[29][246] = 16'b0000000000001110;
    assign weights1[29][247] = 16'b0000000000100100;
    assign weights1[29][248] = 16'b0000000000001110;
    assign weights1[29][249] = 16'b0000000000011010;
    assign weights1[29][250] = 16'b0000000000001001;
    assign weights1[29][251] = 16'b0000000000000101;
    assign weights1[29][252] = 16'b1111111111111000;
    assign weights1[29][253] = 16'b1111111111101110;
    assign weights1[29][254] = 16'b1111111111101010;
    assign weights1[29][255] = 16'b1111111111010111;
    assign weights1[29][256] = 16'b1111111111110011;
    assign weights1[29][257] = 16'b1111111111111100;
    assign weights1[29][258] = 16'b0000000000001000;
    assign weights1[29][259] = 16'b0000000000001011;
    assign weights1[29][260] = 16'b0000000000010000;
    assign weights1[29][261] = 16'b0000000000001100;
    assign weights1[29][262] = 16'b0000000000010100;
    assign weights1[29][263] = 16'b1111111111001111;
    assign weights1[29][264] = 16'b1111111110011100;
    assign weights1[29][265] = 16'b1111111111000001;
    assign weights1[29][266] = 16'b1111111111001101;
    assign weights1[29][267] = 16'b1111111111111010;
    assign weights1[29][268] = 16'b0000000000010101;
    assign weights1[29][269] = 16'b0000000000001011;
    assign weights1[29][270] = 16'b0000000000011011;
    assign weights1[29][271] = 16'b0000000000001100;
    assign weights1[29][272] = 16'b0000000000001000;
    assign weights1[29][273] = 16'b0000000000011110;
    assign weights1[29][274] = 16'b0000000000001011;
    assign weights1[29][275] = 16'b0000000000000111;
    assign weights1[29][276] = 16'b1111111111111110;
    assign weights1[29][277] = 16'b0000000000001101;
    assign weights1[29][278] = 16'b0000000000010011;
    assign weights1[29][279] = 16'b0000000000001011;
    assign weights1[29][280] = 16'b1111111111110111;
    assign weights1[29][281] = 16'b1111111111110101;
    assign weights1[29][282] = 16'b1111111111100001;
    assign weights1[29][283] = 16'b1111111111011110;
    assign weights1[29][284] = 16'b0000000000000000;
    assign weights1[29][285] = 16'b1111111111110011;
    assign weights1[29][286] = 16'b1111111111110010;
    assign weights1[29][287] = 16'b0000000000001010;
    assign weights1[29][288] = 16'b0000000000001111;
    assign weights1[29][289] = 16'b0000000000001101;
    assign weights1[29][290] = 16'b0000000000001001;
    assign weights1[29][291] = 16'b1111111110110011;
    assign weights1[29][292] = 16'b1111111110110010;
    assign weights1[29][293] = 16'b1111111111100100;
    assign weights1[29][294] = 16'b0000000000000110;
    assign weights1[29][295] = 16'b1111111111111110;
    assign weights1[29][296] = 16'b0000000000011110;
    assign weights1[29][297] = 16'b0000000000011111;
    assign weights1[29][298] = 16'b0000000000010001;
    assign weights1[29][299] = 16'b0000000000011011;
    assign weights1[29][300] = 16'b0000000000010011;
    assign weights1[29][301] = 16'b0000000000010001;
    assign weights1[29][302] = 16'b1111111111111011;
    assign weights1[29][303] = 16'b0000000000000010;
    assign weights1[29][304] = 16'b0000000000011010;
    assign weights1[29][305] = 16'b0000000000001010;
    assign weights1[29][306] = 16'b0000000000011101;
    assign weights1[29][307] = 16'b0000000000001100;
    assign weights1[29][308] = 16'b0000000000000001;
    assign weights1[29][309] = 16'b1111111111111001;
    assign weights1[29][310] = 16'b1111111111100000;
    assign weights1[29][311] = 16'b1111111111101101;
    assign weights1[29][312] = 16'b1111111111110000;
    assign weights1[29][313] = 16'b1111111111110010;
    assign weights1[29][314] = 16'b1111111111111101;
    assign weights1[29][315] = 16'b0000000000010000;
    assign weights1[29][316] = 16'b0000000000010000;
    assign weights1[29][317] = 16'b0000000000100000;
    assign weights1[29][318] = 16'b1111111111101000;
    assign weights1[29][319] = 16'b1111111111010000;
    assign weights1[29][320] = 16'b1111111111001010;
    assign weights1[29][321] = 16'b1111111111110001;
    assign weights1[29][322] = 16'b0000000000000000;
    assign weights1[29][323] = 16'b0000000000001000;
    assign weights1[29][324] = 16'b0000000000100000;
    assign weights1[29][325] = 16'b0000000000001111;
    assign weights1[29][326] = 16'b0000000000101001;
    assign weights1[29][327] = 16'b0000000000000100;
    assign weights1[29][328] = 16'b0000000000010010;
    assign weights1[29][329] = 16'b0000000000001100;
    assign weights1[29][330] = 16'b0000000000001000;
    assign weights1[29][331] = 16'b0000000000010011;
    assign weights1[29][332] = 16'b0000000000000011;
    assign weights1[29][333] = 16'b1111111111110100;
    assign weights1[29][334] = 16'b0000000000000011;
    assign weights1[29][335] = 16'b0000000000010101;
    assign weights1[29][336] = 16'b1111111111111111;
    assign weights1[29][337] = 16'b1111111111110111;
    assign weights1[29][338] = 16'b1111111111101111;
    assign weights1[29][339] = 16'b1111111111100100;
    assign weights1[29][340] = 16'b0000000000000011;
    assign weights1[29][341] = 16'b0000000000001001;
    assign weights1[29][342] = 16'b0000000000000011;
    assign weights1[29][343] = 16'b0000000000001110;
    assign weights1[29][344] = 16'b1111111111110100;
    assign weights1[29][345] = 16'b0000000000010000;
    assign weights1[29][346] = 16'b1111111111101001;
    assign weights1[29][347] = 16'b1111111111001000;
    assign weights1[29][348] = 16'b1111111111010001;
    assign weights1[29][349] = 16'b1111111111110000;
    assign weights1[29][350] = 16'b0000000000000110;
    assign weights1[29][351] = 16'b0000000000001101;
    assign weights1[29][352] = 16'b0000000000001110;
    assign weights1[29][353] = 16'b0000000000000101;
    assign weights1[29][354] = 16'b0000000000010000;
    assign weights1[29][355] = 16'b0000000000010011;
    assign weights1[29][356] = 16'b1111111111111000;
    assign weights1[29][357] = 16'b1111111111010101;
    assign weights1[29][358] = 16'b1111111111000110;
    assign weights1[29][359] = 16'b1111111111000001;
    assign weights1[29][360] = 16'b1111111111001111;
    assign weights1[29][361] = 16'b1111111111000010;
    assign weights1[29][362] = 16'b1111111111011100;
    assign weights1[29][363] = 16'b1111111111101000;
    assign weights1[29][364] = 16'b1111111111111010;
    assign weights1[29][365] = 16'b0000000000000000;
    assign weights1[29][366] = 16'b0000000000000010;
    assign weights1[29][367] = 16'b1111111111111111;
    assign weights1[29][368] = 16'b1111111111111100;
    assign weights1[29][369] = 16'b1111111111111000;
    assign weights1[29][370] = 16'b1111111111111100;
    assign weights1[29][371] = 16'b1111111111111000;
    assign weights1[29][372] = 16'b0000000000001110;
    assign weights1[29][373] = 16'b0000000000010001;
    assign weights1[29][374] = 16'b0000000000001000;
    assign weights1[29][375] = 16'b1111111111100101;
    assign weights1[29][376] = 16'b1111111111110001;
    assign weights1[29][377] = 16'b1111111111110101;
    assign weights1[29][378] = 16'b0000000000001010;
    assign weights1[29][379] = 16'b0000000000000010;
    assign weights1[29][380] = 16'b0000000000001111;
    assign weights1[29][381] = 16'b1111111111111110;
    assign weights1[29][382] = 16'b0000000000000011;
    assign weights1[29][383] = 16'b1111111111101001;
    assign weights1[29][384] = 16'b1111111111011011;
    assign weights1[29][385] = 16'b1111111111001110;
    assign weights1[29][386] = 16'b1111111111001110;
    assign weights1[29][387] = 16'b1111111111000000;
    assign weights1[29][388] = 16'b1111111111000111;
    assign weights1[29][389] = 16'b1111111111000000;
    assign weights1[29][390] = 16'b1111111111001001;
    assign weights1[29][391] = 16'b1111111111011100;
    assign weights1[29][392] = 16'b1111111111111000;
    assign weights1[29][393] = 16'b1111111111111111;
    assign weights1[29][394] = 16'b1111111111111110;
    assign weights1[29][395] = 16'b0000000000000111;
    assign weights1[29][396] = 16'b0000000000000011;
    assign weights1[29][397] = 16'b1111111111111100;
    assign weights1[29][398] = 16'b0000000000010011;
    assign weights1[29][399] = 16'b1111111111111100;
    assign weights1[29][400] = 16'b0000000000000100;
    assign weights1[29][401] = 16'b1111111111110111;
    assign weights1[29][402] = 16'b0000000000010101;
    assign weights1[29][403] = 16'b1111111111111110;
    assign weights1[29][404] = 16'b1111111111101001;
    assign weights1[29][405] = 16'b1111111111111110;
    assign weights1[29][406] = 16'b1111111111111110;
    assign weights1[29][407] = 16'b0000000000010011;
    assign weights1[29][408] = 16'b0000000000000011;
    assign weights1[29][409] = 16'b1111111111111110;
    assign weights1[29][410] = 16'b1111111111110000;
    assign weights1[29][411] = 16'b1111111111101100;
    assign weights1[29][412] = 16'b1111111111110110;
    assign weights1[29][413] = 16'b1111111111110010;
    assign weights1[29][414] = 16'b0000000000000100;
    assign weights1[29][415] = 16'b1111111111110100;
    assign weights1[29][416] = 16'b1111111111100100;
    assign weights1[29][417] = 16'b1111111111010110;
    assign weights1[29][418] = 16'b1111111111011001;
    assign weights1[29][419] = 16'b1111111111100100;
    assign weights1[29][420] = 16'b1111111111111011;
    assign weights1[29][421] = 16'b1111111111111000;
    assign weights1[29][422] = 16'b1111111111111100;
    assign weights1[29][423] = 16'b1111111111110111;
    assign weights1[29][424] = 16'b1111111111110100;
    assign weights1[29][425] = 16'b0000000000000010;
    assign weights1[29][426] = 16'b1111111111111110;
    assign weights1[29][427] = 16'b0000000000010000;
    assign weights1[29][428] = 16'b1111111111111001;
    assign weights1[29][429] = 16'b0000000000011101;
    assign weights1[29][430] = 16'b0000000000000101;
    assign weights1[29][431] = 16'b0000000000000010;
    assign weights1[29][432] = 16'b1111111111111001;
    assign weights1[29][433] = 16'b0000000000000000;
    assign weights1[29][434] = 16'b1111111111110100;
    assign weights1[29][435] = 16'b0000000000000101;
    assign weights1[29][436] = 16'b0000000000000101;
    assign weights1[29][437] = 16'b1111111111101000;
    assign weights1[29][438] = 16'b1111111111101100;
    assign weights1[29][439] = 16'b1111111111101100;
    assign weights1[29][440] = 16'b0000000000000000;
    assign weights1[29][441] = 16'b0000000000000100;
    assign weights1[29][442] = 16'b1111111111111110;
    assign weights1[29][443] = 16'b0000000000001000;
    assign weights1[29][444] = 16'b1111111111111101;
    assign weights1[29][445] = 16'b1111111111110111;
    assign weights1[29][446] = 16'b1111111111110000;
    assign weights1[29][447] = 16'b1111111111101001;
    assign weights1[29][448] = 16'b1111111111110011;
    assign weights1[29][449] = 16'b1111111111111101;
    assign weights1[29][450] = 16'b0000000000000001;
    assign weights1[29][451] = 16'b0000000000000111;
    assign weights1[29][452] = 16'b0000000000000001;
    assign weights1[29][453] = 16'b0000000000001100;
    assign weights1[29][454] = 16'b0000000000010111;
    assign weights1[29][455] = 16'b0000000000001001;
    assign weights1[29][456] = 16'b0000000000001111;
    assign weights1[29][457] = 16'b0000000000010010;
    assign weights1[29][458] = 16'b1111111111111110;
    assign weights1[29][459] = 16'b0000000000001100;
    assign weights1[29][460] = 16'b1111111111111000;
    assign weights1[29][461] = 16'b0000000000001100;
    assign weights1[29][462] = 16'b1111111111101101;
    assign weights1[29][463] = 16'b1111111111111100;
    assign weights1[29][464] = 16'b1111111111111100;
    assign weights1[29][465] = 16'b0000000000000000;
    assign weights1[29][466] = 16'b1111111111101010;
    assign weights1[29][467] = 16'b1111111111110111;
    assign weights1[29][468] = 16'b1111111111011101;
    assign weights1[29][469] = 16'b1111111111101111;
    assign weights1[29][470] = 16'b1111111111110011;
    assign weights1[29][471] = 16'b0000000000001100;
    assign weights1[29][472] = 16'b0000000000001010;
    assign weights1[29][473] = 16'b0000000000001111;
    assign weights1[29][474] = 16'b0000000000001001;
    assign weights1[29][475] = 16'b1111111111111001;
    assign weights1[29][476] = 16'b1111111111110100;
    assign weights1[29][477] = 16'b0000000000001010;
    assign weights1[29][478] = 16'b0000000000001100;
    assign weights1[29][479] = 16'b1111111111111011;
    assign weights1[29][480] = 16'b1111111111110110;
    assign weights1[29][481] = 16'b0000000000001110;
    assign weights1[29][482] = 16'b0000000000000101;
    assign weights1[29][483] = 16'b0000000000000010;
    assign weights1[29][484] = 16'b1111111111111100;
    assign weights1[29][485] = 16'b0000000000001101;
    assign weights1[29][486] = 16'b1111111111111100;
    assign weights1[29][487] = 16'b0000000000010000;
    assign weights1[29][488] = 16'b0000000000000000;
    assign weights1[29][489] = 16'b0000000000000101;
    assign weights1[29][490] = 16'b1111111111101100;
    assign weights1[29][491] = 16'b1111111111111011;
    assign weights1[29][492] = 16'b1111111111111001;
    assign weights1[29][493] = 16'b1111111111110111;
    assign weights1[29][494] = 16'b0000000000001000;
    assign weights1[29][495] = 16'b1111111111101101;
    assign weights1[29][496] = 16'b1111111111111110;
    assign weights1[29][497] = 16'b1111111111111110;
    assign weights1[29][498] = 16'b0000000000010001;
    assign weights1[29][499] = 16'b1111111111111101;
    assign weights1[29][500] = 16'b0000000000000010;
    assign weights1[29][501] = 16'b0000000000001101;
    assign weights1[29][502] = 16'b0000000000000100;
    assign weights1[29][503] = 16'b1111111111111010;
    assign weights1[29][504] = 16'b1111111111110111;
    assign weights1[29][505] = 16'b0000000000010001;
    assign weights1[29][506] = 16'b0000000000001010;
    assign weights1[29][507] = 16'b1111111111111010;
    assign weights1[29][508] = 16'b1111111111010111;
    assign weights1[29][509] = 16'b0000000000000011;
    assign weights1[29][510] = 16'b1111111111110100;
    assign weights1[29][511] = 16'b0000000000001001;
    assign weights1[29][512] = 16'b1111111111111000;
    assign weights1[29][513] = 16'b0000000000000001;
    assign weights1[29][514] = 16'b0000000000000011;
    assign weights1[29][515] = 16'b0000000000001010;
    assign weights1[29][516] = 16'b0000000000001001;
    assign weights1[29][517] = 16'b1111111111101110;
    assign weights1[29][518] = 16'b1111111111111101;
    assign weights1[29][519] = 16'b1111111111110001;
    assign weights1[29][520] = 16'b1111111111110101;
    assign weights1[29][521] = 16'b1111111111110101;
    assign weights1[29][522] = 16'b1111111111111101;
    assign weights1[29][523] = 16'b1111111111111011;
    assign weights1[29][524] = 16'b1111111111110011;
    assign weights1[29][525] = 16'b1111111111110111;
    assign weights1[29][526] = 16'b0000000000001010;
    assign weights1[29][527] = 16'b0000000000011010;
    assign weights1[29][528] = 16'b0000000000000000;
    assign weights1[29][529] = 16'b0000000000000001;
    assign weights1[29][530] = 16'b0000000000001001;
    assign weights1[29][531] = 16'b1111111111110011;
    assign weights1[29][532] = 16'b1111111111111000;
    assign weights1[29][533] = 16'b0000000000001011;
    assign weights1[29][534] = 16'b0000000000010011;
    assign weights1[29][535] = 16'b0000000000001100;
    assign weights1[29][536] = 16'b1111111111110000;
    assign weights1[29][537] = 16'b1111111111111110;
    assign weights1[29][538] = 16'b0000000000011000;
    assign weights1[29][539] = 16'b1111111111111111;
    assign weights1[29][540] = 16'b1111111111110011;
    assign weights1[29][541] = 16'b0000000000010101;
    assign weights1[29][542] = 16'b0000000000000001;
    assign weights1[29][543] = 16'b0000000000001011;
    assign weights1[29][544] = 16'b0000000000000000;
    assign weights1[29][545] = 16'b0000000000001101;
    assign weights1[29][546] = 16'b0000000000001001;
    assign weights1[29][547] = 16'b1111111111111110;
    assign weights1[29][548] = 16'b1111111111111010;
    assign weights1[29][549] = 16'b1111111111111001;
    assign weights1[29][550] = 16'b1111111111111011;
    assign weights1[29][551] = 16'b1111111111100011;
    assign weights1[29][552] = 16'b0000000000001101;
    assign weights1[29][553] = 16'b0000000000000011;
    assign weights1[29][554] = 16'b0000000000010011;
    assign weights1[29][555] = 16'b0000000000000000;
    assign weights1[29][556] = 16'b1111111111111100;
    assign weights1[29][557] = 16'b0000000000000000;
    assign weights1[29][558] = 16'b0000000000000001;
    assign weights1[29][559] = 16'b0000000000000100;
    assign weights1[29][560] = 16'b0000000000000001;
    assign weights1[29][561] = 16'b1111111111111001;
    assign weights1[29][562] = 16'b0000000000001001;
    assign weights1[29][563] = 16'b0000000000001000;
    assign weights1[29][564] = 16'b0000000000001101;
    assign weights1[29][565] = 16'b1111111111110110;
    assign weights1[29][566] = 16'b0000000000000101;
    assign weights1[29][567] = 16'b1111111111111100;
    assign weights1[29][568] = 16'b0000000000000000;
    assign weights1[29][569] = 16'b0000000000001110;
    assign weights1[29][570] = 16'b0000000000010010;
    assign weights1[29][571] = 16'b1111111111111011;
    assign weights1[29][572] = 16'b0000000000010110;
    assign weights1[29][573] = 16'b0000000000000000;
    assign weights1[29][574] = 16'b0000000000000011;
    assign weights1[29][575] = 16'b1111111111111001;
    assign weights1[29][576] = 16'b1111111111110011;
    assign weights1[29][577] = 16'b1111111111111101;
    assign weights1[29][578] = 16'b1111111111110101;
    assign weights1[29][579] = 16'b0000000000000001;
    assign weights1[29][580] = 16'b1111111111111000;
    assign weights1[29][581] = 16'b1111111111111101;
    assign weights1[29][582] = 16'b1111111111111000;
    assign weights1[29][583] = 16'b1111111111111001;
    assign weights1[29][584] = 16'b0000000000010010;
    assign weights1[29][585] = 16'b1111111111111110;
    assign weights1[29][586] = 16'b0000000000000110;
    assign weights1[29][587] = 16'b0000000000000101;
    assign weights1[29][588] = 16'b0000000000000010;
    assign weights1[29][589] = 16'b1111111111111011;
    assign weights1[29][590] = 16'b1111111111111111;
    assign weights1[29][591] = 16'b0000000000000001;
    assign weights1[29][592] = 16'b0000000000010110;
    assign weights1[29][593] = 16'b0000000000001101;
    assign weights1[29][594] = 16'b0000000000000111;
    assign weights1[29][595] = 16'b1111111111111100;
    assign weights1[29][596] = 16'b0000000000010101;
    assign weights1[29][597] = 16'b1111111111110000;
    assign weights1[29][598] = 16'b1111111111111110;
    assign weights1[29][599] = 16'b1111111111111001;
    assign weights1[29][600] = 16'b1111111111111101;
    assign weights1[29][601] = 16'b1111111111110011;
    assign weights1[29][602] = 16'b1111111111111101;
    assign weights1[29][603] = 16'b0000000000001100;
    assign weights1[29][604] = 16'b1111111111111110;
    assign weights1[29][605] = 16'b1111111111110001;
    assign weights1[29][606] = 16'b1111111111110111;
    assign weights1[29][607] = 16'b1111111111110001;
    assign weights1[29][608] = 16'b0000000000000101;
    assign weights1[29][609] = 16'b0000000000010000;
    assign weights1[29][610] = 16'b1111111111111001;
    assign weights1[29][611] = 16'b0000000000000110;
    assign weights1[29][612] = 16'b0000000000010110;
    assign weights1[29][613] = 16'b1111111111110010;
    assign weights1[29][614] = 16'b0000000000000000;
    assign weights1[29][615] = 16'b1111111111110101;
    assign weights1[29][616] = 16'b0000000000000001;
    assign weights1[29][617] = 16'b1111111111111101;
    assign weights1[29][618] = 16'b1111111111111111;
    assign weights1[29][619] = 16'b1111111111110100;
    assign weights1[29][620] = 16'b0000000000001010;
    assign weights1[29][621] = 16'b0000000000000100;
    assign weights1[29][622] = 16'b0000000000001101;
    assign weights1[29][623] = 16'b1111111111101111;
    assign weights1[29][624] = 16'b1111111111111001;
    assign weights1[29][625] = 16'b0000000000000110;
    assign weights1[29][626] = 16'b0000000000010100;
    assign weights1[29][627] = 16'b0000000000000011;
    assign weights1[29][628] = 16'b0000000000001000;
    assign weights1[29][629] = 16'b0000000000000011;
    assign weights1[29][630] = 16'b1111111111111001;
    assign weights1[29][631] = 16'b1111111111111010;
    assign weights1[29][632] = 16'b1111111111111000;
    assign weights1[29][633] = 16'b1111111111110110;
    assign weights1[29][634] = 16'b0000000000001001;
    assign weights1[29][635] = 16'b1111111111111100;
    assign weights1[29][636] = 16'b1111111111111101;
    assign weights1[29][637] = 16'b1111111111101111;
    assign weights1[29][638] = 16'b0000000000000010;
    assign weights1[29][639] = 16'b0000000000001010;
    assign weights1[29][640] = 16'b0000000000010100;
    assign weights1[29][641] = 16'b1111111111111101;
    assign weights1[29][642] = 16'b1111111111111111;
    assign weights1[29][643] = 16'b1111111111111101;
    assign weights1[29][644] = 16'b1111111111111001;
    assign weights1[29][645] = 16'b1111111111111101;
    assign weights1[29][646] = 16'b1111111111111011;
    assign weights1[29][647] = 16'b0000000000000000;
    assign weights1[29][648] = 16'b1111111111111000;
    assign weights1[29][649] = 16'b0000000000000100;
    assign weights1[29][650] = 16'b0000000000000111;
    assign weights1[29][651] = 16'b1111111111111101;
    assign weights1[29][652] = 16'b0000000000000001;
    assign weights1[29][653] = 16'b0000000000000000;
    assign weights1[29][654] = 16'b0000000000001110;
    assign weights1[29][655] = 16'b0000000000000101;
    assign weights1[29][656] = 16'b0000000000001111;
    assign weights1[29][657] = 16'b0000000000000011;
    assign weights1[29][658] = 16'b0000000000001010;
    assign weights1[29][659] = 16'b0000000000010010;
    assign weights1[29][660] = 16'b0000000000000011;
    assign weights1[29][661] = 16'b0000000000000010;
    assign weights1[29][662] = 16'b0000000000000001;
    assign weights1[29][663] = 16'b1111111111110001;
    assign weights1[29][664] = 16'b0000000000000001;
    assign weights1[29][665] = 16'b0000000000001100;
    assign weights1[29][666] = 16'b0000000000010110;
    assign weights1[29][667] = 16'b1111111111111100;
    assign weights1[29][668] = 16'b1111111111110111;
    assign weights1[29][669] = 16'b0000000000000000;
    assign weights1[29][670] = 16'b0000000000000000;
    assign weights1[29][671] = 16'b1111111111110011;
    assign weights1[29][672] = 16'b1111111111111000;
    assign weights1[29][673] = 16'b1111111111111101;
    assign weights1[29][674] = 16'b0000000000000000;
    assign weights1[29][675] = 16'b1111111111101010;
    assign weights1[29][676] = 16'b1111111111111101;
    assign weights1[29][677] = 16'b0000000000000010;
    assign weights1[29][678] = 16'b1111111111110010;
    assign weights1[29][679] = 16'b1111111111110100;
    assign weights1[29][680] = 16'b1111111111110001;
    assign weights1[29][681] = 16'b1111111111111011;
    assign weights1[29][682] = 16'b1111111111110000;
    assign weights1[29][683] = 16'b0000000000000001;
    assign weights1[29][684] = 16'b0000000000000010;
    assign weights1[29][685] = 16'b1111111111111110;
    assign weights1[29][686] = 16'b0000000000000100;
    assign weights1[29][687] = 16'b1111111111111011;
    assign weights1[29][688] = 16'b1111111111111111;
    assign weights1[29][689] = 16'b0000000000001110;
    assign weights1[29][690] = 16'b0000000000000100;
    assign weights1[29][691] = 16'b0000000000001010;
    assign weights1[29][692] = 16'b0000000000001101;
    assign weights1[29][693] = 16'b0000000000001100;
    assign weights1[29][694] = 16'b0000000000000111;
    assign weights1[29][695] = 16'b0000000000000010;
    assign weights1[29][696] = 16'b1111111111111010;
    assign weights1[29][697] = 16'b1111111111111001;
    assign weights1[29][698] = 16'b1111111111111000;
    assign weights1[29][699] = 16'b1111111111110100;
    assign weights1[29][700] = 16'b1111111111111111;
    assign weights1[29][701] = 16'b1111111111110110;
    assign weights1[29][702] = 16'b1111111111110100;
    assign weights1[29][703] = 16'b1111111111111010;
    assign weights1[29][704] = 16'b1111111111111010;
    assign weights1[29][705] = 16'b0000000000001010;
    assign weights1[29][706] = 16'b1111111111110111;
    assign weights1[29][707] = 16'b1111111111111001;
    assign weights1[29][708] = 16'b0000000000001010;
    assign weights1[29][709] = 16'b1111111111111101;
    assign weights1[29][710] = 16'b1111111111111100;
    assign weights1[29][711] = 16'b0000000000001010;
    assign weights1[29][712] = 16'b1111111111101111;
    assign weights1[29][713] = 16'b1111111111111110;
    assign weights1[29][714] = 16'b1111111111111101;
    assign weights1[29][715] = 16'b0000000000000011;
    assign weights1[29][716] = 16'b0000000000010010;
    assign weights1[29][717] = 16'b1111111111111101;
    assign weights1[29][718] = 16'b0000000000010000;
    assign weights1[29][719] = 16'b1111111111110010;
    assign weights1[29][720] = 16'b1111111111110001;
    assign weights1[29][721] = 16'b0000000000001001;
    assign weights1[29][722] = 16'b0000000000001101;
    assign weights1[29][723] = 16'b0000000000000011;
    assign weights1[29][724] = 16'b1111111111100100;
    assign weights1[29][725] = 16'b1111111111111010;
    assign weights1[29][726] = 16'b0000000000000100;
    assign weights1[29][727] = 16'b1111111111111001;
    assign weights1[29][728] = 16'b1111111111111111;
    assign weights1[29][729] = 16'b1111111111111111;
    assign weights1[29][730] = 16'b1111111111110111;
    assign weights1[29][731] = 16'b1111111111111100;
    assign weights1[29][732] = 16'b0000000000000111;
    assign weights1[29][733] = 16'b1111111111110000;
    assign weights1[29][734] = 16'b1111111111110011;
    assign weights1[29][735] = 16'b1111111111110100;
    assign weights1[29][736] = 16'b1111111111110001;
    assign weights1[29][737] = 16'b1111111111111100;
    assign weights1[29][738] = 16'b0000000000001011;
    assign weights1[29][739] = 16'b1111111111110100;
    assign weights1[29][740] = 16'b1111111111111010;
    assign weights1[29][741] = 16'b1111111111110110;
    assign weights1[29][742] = 16'b1111111111111100;
    assign weights1[29][743] = 16'b1111111111101010;
    assign weights1[29][744] = 16'b1111111111110001;
    assign weights1[29][745] = 16'b1111111111110100;
    assign weights1[29][746] = 16'b1111111111111001;
    assign weights1[29][747] = 16'b1111111111101100;
    assign weights1[29][748] = 16'b0000000000001001;
    assign weights1[29][749] = 16'b1111111111011100;
    assign weights1[29][750] = 16'b1111111111111011;
    assign weights1[29][751] = 16'b1111111111111000;
    assign weights1[29][752] = 16'b1111111111101111;
    assign weights1[29][753] = 16'b1111111111111001;
    assign weights1[29][754] = 16'b1111111111110110;
    assign weights1[29][755] = 16'b1111111111111010;
    assign weights1[29][756] = 16'b0000000000000000;
    assign weights1[29][757] = 16'b0000000000000111;
    assign weights1[29][758] = 16'b0000000000000001;
    assign weights1[29][759] = 16'b1111111111111111;
    assign weights1[29][760] = 16'b0000000000000010;
    assign weights1[29][761] = 16'b1111111111110110;
    assign weights1[29][762] = 16'b1111111111101001;
    assign weights1[29][763] = 16'b1111111111111011;
    assign weights1[29][764] = 16'b0000000000000010;
    assign weights1[29][765] = 16'b1111111111111000;
    assign weights1[29][766] = 16'b1111111111110000;
    assign weights1[29][767] = 16'b1111111111110010;
    assign weights1[29][768] = 16'b1111111111111010;
    assign weights1[29][769] = 16'b1111111111110111;
    assign weights1[29][770] = 16'b1111111111110111;
    assign weights1[29][771] = 16'b1111111111110010;
    assign weights1[29][772] = 16'b1111111111111110;
    assign weights1[29][773] = 16'b1111111111111011;
    assign weights1[29][774] = 16'b0000000000000000;
    assign weights1[29][775] = 16'b1111111111111011;
    assign weights1[29][776] = 16'b1111111111111010;
    assign weights1[29][777] = 16'b1111111111100110;
    assign weights1[29][778] = 16'b1111111111111000;
    assign weights1[29][779] = 16'b1111111111101010;
    assign weights1[29][780] = 16'b1111111111101101;
    assign weights1[29][781] = 16'b1111111111111000;
    assign weights1[29][782] = 16'b1111111111111010;
    assign weights1[29][783] = 16'b1111111111111110;
    assign weights1[30][0] = 16'b0000000000000000;
    assign weights1[30][1] = 16'b0000000000000000;
    assign weights1[30][2] = 16'b0000000000000001;
    assign weights1[30][3] = 16'b0000000000000010;
    assign weights1[30][4] = 16'b0000000000000001;
    assign weights1[30][5] = 16'b0000000000000010;
    assign weights1[30][6] = 16'b1111111111111100;
    assign weights1[30][7] = 16'b0000000000000011;
    assign weights1[30][8] = 16'b1111111111111000;
    assign weights1[30][9] = 16'b1111111111111111;
    assign weights1[30][10] = 16'b1111111111111100;
    assign weights1[30][11] = 16'b0000000000000100;
    assign weights1[30][12] = 16'b0000000000010001;
    assign weights1[30][13] = 16'b0000000000010000;
    assign weights1[30][14] = 16'b0000000000011100;
    assign weights1[30][15] = 16'b0000000000001110;
    assign weights1[30][16] = 16'b0000000000000001;
    assign weights1[30][17] = 16'b1111111111110110;
    assign weights1[30][18] = 16'b1111111111110100;
    assign weights1[30][19] = 16'b1111111111111001;
    assign weights1[30][20] = 16'b1111111111110110;
    assign weights1[30][21] = 16'b1111111111110100;
    assign weights1[30][22] = 16'b1111111111111010;
    assign weights1[30][23] = 16'b1111111111111001;
    assign weights1[30][24] = 16'b1111111111111100;
    assign weights1[30][25] = 16'b1111111111111111;
    assign weights1[30][26] = 16'b0000000000000000;
    assign weights1[30][27] = 16'b0000000000000000;
    assign weights1[30][28] = 16'b0000000000000000;
    assign weights1[30][29] = 16'b0000000000000000;
    assign weights1[30][30] = 16'b0000000000000001;
    assign weights1[30][31] = 16'b0000000000000001;
    assign weights1[30][32] = 16'b0000000000000000;
    assign weights1[30][33] = 16'b1111111111111111;
    assign weights1[30][34] = 16'b1111111111111000;
    assign weights1[30][35] = 16'b1111111111101111;
    assign weights1[30][36] = 16'b1111111111101101;
    assign weights1[30][37] = 16'b1111111111110111;
    assign weights1[30][38] = 16'b0000000000000010;
    assign weights1[30][39] = 16'b0000000000000011;
    assign weights1[30][40] = 16'b1111111111111111;
    assign weights1[30][41] = 16'b1111111111111110;
    assign weights1[30][42] = 16'b0000000000010010;
    assign weights1[30][43] = 16'b0000000000010111;
    assign weights1[30][44] = 16'b1111111111111101;
    assign weights1[30][45] = 16'b0000000000000110;
    assign weights1[30][46] = 16'b0000000000001001;
    assign weights1[30][47] = 16'b1111111111111111;
    assign weights1[30][48] = 16'b1111111111101100;
    assign weights1[30][49] = 16'b1111111111110011;
    assign weights1[30][50] = 16'b1111111111110101;
    assign weights1[30][51] = 16'b1111111111101100;
    assign weights1[30][52] = 16'b1111111111111100;
    assign weights1[30][53] = 16'b0000000000000000;
    assign weights1[30][54] = 16'b0000000000000001;
    assign weights1[30][55] = 16'b0000000000000000;
    assign weights1[30][56] = 16'b0000000000000000;
    assign weights1[30][57] = 16'b0000000000000000;
    assign weights1[30][58] = 16'b0000000000000000;
    assign weights1[30][59] = 16'b0000000000000001;
    assign weights1[30][60] = 16'b1111111111110111;
    assign weights1[30][61] = 16'b1111111111110101;
    assign weights1[30][62] = 16'b1111111111110010;
    assign weights1[30][63] = 16'b1111111111100101;
    assign weights1[30][64] = 16'b1111111111011011;
    assign weights1[30][65] = 16'b1111111111100011;
    assign weights1[30][66] = 16'b1111111111011101;
    assign weights1[30][67] = 16'b1111111111100011;
    assign weights1[30][68] = 16'b1111111111100001;
    assign weights1[30][69] = 16'b1111111111111011;
    assign weights1[30][70] = 16'b0000000000000001;
    assign weights1[30][71] = 16'b1111111111111111;
    assign weights1[30][72] = 16'b1111111111110110;
    assign weights1[30][73] = 16'b1111111111110110;
    assign weights1[30][74] = 16'b1111111111111111;
    assign weights1[30][75] = 16'b0000000000000110;
    assign weights1[30][76] = 16'b1111111111101111;
    assign weights1[30][77] = 16'b1111111111110100;
    assign weights1[30][78] = 16'b1111111111101010;
    assign weights1[30][79] = 16'b1111111111101110;
    assign weights1[30][80] = 16'b1111111111110111;
    assign weights1[30][81] = 16'b1111111111111111;
    assign weights1[30][82] = 16'b0000000000000000;
    assign weights1[30][83] = 16'b0000000000000000;
    assign weights1[30][84] = 16'b0000000000000001;
    assign weights1[30][85] = 16'b0000000000000001;
    assign weights1[30][86] = 16'b0000000000000001;
    assign weights1[30][87] = 16'b1111111111111111;
    assign weights1[30][88] = 16'b1111111111110110;
    assign weights1[30][89] = 16'b1111111111110000;
    assign weights1[30][90] = 16'b1111111111101100;
    assign weights1[30][91] = 16'b1111111111011011;
    assign weights1[30][92] = 16'b1111111111000101;
    assign weights1[30][93] = 16'b1111111111000111;
    assign weights1[30][94] = 16'b1111111111001101;
    assign weights1[30][95] = 16'b1111111111100111;
    assign weights1[30][96] = 16'b1111111111101111;
    assign weights1[30][97] = 16'b1111111111111000;
    assign weights1[30][98] = 16'b1111111111111000;
    assign weights1[30][99] = 16'b1111111111110011;
    assign weights1[30][100] = 16'b1111111111110001;
    assign weights1[30][101] = 16'b1111111111110000;
    assign weights1[30][102] = 16'b1111111111110111;
    assign weights1[30][103] = 16'b1111111111110000;
    assign weights1[30][104] = 16'b1111111111100100;
    assign weights1[30][105] = 16'b1111111111100111;
    assign weights1[30][106] = 16'b1111111111111000;
    assign weights1[30][107] = 16'b1111111111110101;
    assign weights1[30][108] = 16'b1111111111110100;
    assign weights1[30][109] = 16'b1111111111111000;
    assign weights1[30][110] = 16'b1111111111111111;
    assign weights1[30][111] = 16'b0000000000000000;
    assign weights1[30][112] = 16'b1111111111111111;
    assign weights1[30][113] = 16'b0000000000000000;
    assign weights1[30][114] = 16'b0000000000000000;
    assign weights1[30][115] = 16'b1111111111110101;
    assign weights1[30][116] = 16'b1111111111111011;
    assign weights1[30][117] = 16'b1111111111110111;
    assign weights1[30][118] = 16'b1111111111101110;
    assign weights1[30][119] = 16'b1111111111010110;
    assign weights1[30][120] = 16'b1111111111101010;
    assign weights1[30][121] = 16'b1111111111101101;
    assign weights1[30][122] = 16'b1111111111111011;
    assign weights1[30][123] = 16'b0000000000000000;
    assign weights1[30][124] = 16'b1111111111101111;
    assign weights1[30][125] = 16'b0000000000010110;
    assign weights1[30][126] = 16'b1111111111111010;
    assign weights1[30][127] = 16'b0000000000001111;
    assign weights1[30][128] = 16'b0000000000001000;
    assign weights1[30][129] = 16'b0000000000001100;
    assign weights1[30][130] = 16'b0000000000010011;
    assign weights1[30][131] = 16'b1111111111111000;
    assign weights1[30][132] = 16'b1111111111111010;
    assign weights1[30][133] = 16'b1111111111110100;
    assign weights1[30][134] = 16'b1111111111010010;
    assign weights1[30][135] = 16'b1111111111100010;
    assign weights1[30][136] = 16'b1111111111110001;
    assign weights1[30][137] = 16'b1111111111110110;
    assign weights1[30][138] = 16'b1111111111111110;
    assign weights1[30][139] = 16'b1111111111111111;
    assign weights1[30][140] = 16'b1111111111111101;
    assign weights1[30][141] = 16'b0000000000000011;
    assign weights1[30][142] = 16'b1111111111111110;
    assign weights1[30][143] = 16'b1111111111111111;
    assign weights1[30][144] = 16'b0000000000000000;
    assign weights1[30][145] = 16'b1111111111111111;
    assign weights1[30][146] = 16'b0000000000000100;
    assign weights1[30][147] = 16'b0000000000000101;
    assign weights1[30][148] = 16'b1111111111110111;
    assign weights1[30][149] = 16'b0000000000010001;
    assign weights1[30][150] = 16'b1111111111111000;
    assign weights1[30][151] = 16'b1111111111111011;
    assign weights1[30][152] = 16'b0000000000000000;
    assign weights1[30][153] = 16'b0000000000100011;
    assign weights1[30][154] = 16'b0000000000000011;
    assign weights1[30][155] = 16'b0000000000001001;
    assign weights1[30][156] = 16'b0000000000010101;
    assign weights1[30][157] = 16'b1111111111111011;
    assign weights1[30][158] = 16'b0000000000000001;
    assign weights1[30][159] = 16'b0000000000001010;
    assign weights1[30][160] = 16'b1111111111111010;
    assign weights1[30][161] = 16'b1111111111010011;
    assign weights1[30][162] = 16'b1111111111000111;
    assign weights1[30][163] = 16'b1111111111000000;
    assign weights1[30][164] = 16'b1111111111101011;
    assign weights1[30][165] = 16'b1111111111110010;
    assign weights1[30][166] = 16'b1111111111111100;
    assign weights1[30][167] = 16'b0000000000000010;
    assign weights1[30][168] = 16'b1111111111111111;
    assign weights1[30][169] = 16'b0000000000000001;
    assign weights1[30][170] = 16'b1111111111111100;
    assign weights1[30][171] = 16'b0000000000000110;
    assign weights1[30][172] = 16'b0000000000001001;
    assign weights1[30][173] = 16'b0000000000010101;
    assign weights1[30][174] = 16'b0000000000010001;
    assign weights1[30][175] = 16'b0000000000011110;
    assign weights1[30][176] = 16'b0000000000011001;
    assign weights1[30][177] = 16'b0000000000011110;
    assign weights1[30][178] = 16'b0000000000011000;
    assign weights1[30][179] = 16'b0000000000000001;
    assign weights1[30][180] = 16'b1111111111111111;
    assign weights1[30][181] = 16'b0000000000011111;
    assign weights1[30][182] = 16'b0000000000010001;
    assign weights1[30][183] = 16'b0000000000001001;
    assign weights1[30][184] = 16'b0000000000000101;
    assign weights1[30][185] = 16'b0000000000000100;
    assign weights1[30][186] = 16'b0000000000000100;
    assign weights1[30][187] = 16'b1111111111111011;
    assign weights1[30][188] = 16'b0000000000010110;
    assign weights1[30][189] = 16'b1111111111001011;
    assign weights1[30][190] = 16'b1111111111010111;
    assign weights1[30][191] = 16'b1111111111001010;
    assign weights1[30][192] = 16'b1111111111101110;
    assign weights1[30][193] = 16'b1111111111110101;
    assign weights1[30][194] = 16'b1111111111111010;
    assign weights1[30][195] = 16'b1111111111111101;
    assign weights1[30][196] = 16'b0000000000000000;
    assign weights1[30][197] = 16'b0000000000000011;
    assign weights1[30][198] = 16'b0000000000001000;
    assign weights1[30][199] = 16'b0000000000001011;
    assign weights1[30][200] = 16'b0000000000010011;
    assign weights1[30][201] = 16'b0000000000001011;
    assign weights1[30][202] = 16'b0000000000100101;
    assign weights1[30][203] = 16'b0000000000111000;
    assign weights1[30][204] = 16'b0000000000100001;
    assign weights1[30][205] = 16'b0000000000100011;
    assign weights1[30][206] = 16'b0000000000101101;
    assign weights1[30][207] = 16'b0000000000010001;
    assign weights1[30][208] = 16'b0000000000110100;
    assign weights1[30][209] = 16'b0000000000011100;
    assign weights1[30][210] = 16'b0000000000101011;
    assign weights1[30][211] = 16'b0000000000001100;
    assign weights1[30][212] = 16'b0000000000000101;
    assign weights1[30][213] = 16'b0000000000101011;
    assign weights1[30][214] = 16'b0000000000000010;
    assign weights1[30][215] = 16'b1111111111110110;
    assign weights1[30][216] = 16'b0000000000001000;
    assign weights1[30][217] = 16'b1111111111110010;
    assign weights1[30][218] = 16'b1111111111101001;
    assign weights1[30][219] = 16'b1111111111010011;
    assign weights1[30][220] = 16'b1111111111100101;
    assign weights1[30][221] = 16'b1111111111110011;
    assign weights1[30][222] = 16'b1111111111111010;
    assign weights1[30][223] = 16'b1111111111111101;
    assign weights1[30][224] = 16'b0000000000000010;
    assign weights1[30][225] = 16'b0000000000001001;
    assign weights1[30][226] = 16'b0000000000001001;
    assign weights1[30][227] = 16'b0000000000001100;
    assign weights1[30][228] = 16'b0000000000011000;
    assign weights1[30][229] = 16'b0000000000011001;
    assign weights1[30][230] = 16'b0000000000010110;
    assign weights1[30][231] = 16'b0000000000100101;
    assign weights1[30][232] = 16'b0000000000011111;
    assign weights1[30][233] = 16'b0000000000111010;
    assign weights1[30][234] = 16'b0000000000111101;
    assign weights1[30][235] = 16'b0000000000011100;
    assign weights1[30][236] = 16'b1111111111111000;
    assign weights1[30][237] = 16'b0000000000010010;
    assign weights1[30][238] = 16'b0000000000001101;
    assign weights1[30][239] = 16'b0000000000100000;
    assign weights1[30][240] = 16'b0000000000010100;
    assign weights1[30][241] = 16'b0000000000010100;
    assign weights1[30][242] = 16'b0000000000001010;
    assign weights1[30][243] = 16'b0000000000000111;
    assign weights1[30][244] = 16'b1111111111100100;
    assign weights1[30][245] = 16'b1111111111110011;
    assign weights1[30][246] = 16'b1111111111011100;
    assign weights1[30][247] = 16'b1111111111000101;
    assign weights1[30][248] = 16'b1111111111001000;
    assign weights1[30][249] = 16'b1111111111101011;
    assign weights1[30][250] = 16'b1111111111110110;
    assign weights1[30][251] = 16'b1111111111111011;
    assign weights1[30][252] = 16'b0000000000000011;
    assign weights1[30][253] = 16'b0000000000001101;
    assign weights1[30][254] = 16'b1111111111111100;
    assign weights1[30][255] = 16'b0000000000000110;
    assign weights1[30][256] = 16'b0000000000101001;
    assign weights1[30][257] = 16'b0000000000001000;
    assign weights1[30][258] = 16'b0000000000101001;
    assign weights1[30][259] = 16'b0000000001000111;
    assign weights1[30][260] = 16'b0000000000111111;
    assign weights1[30][261] = 16'b0000000000111010;
    assign weights1[30][262] = 16'b1111111111111011;
    assign weights1[30][263] = 16'b1111111111011000;
    assign weights1[30][264] = 16'b1111111110000110;
    assign weights1[30][265] = 16'b1111111110111010;
    assign weights1[30][266] = 16'b1111111111110111;
    assign weights1[30][267] = 16'b0000000000000110;
    assign weights1[30][268] = 16'b0000000000001110;
    assign weights1[30][269] = 16'b0000000000001111;
    assign weights1[30][270] = 16'b1111111111111110;
    assign weights1[30][271] = 16'b0000000000001000;
    assign weights1[30][272] = 16'b1111111111101000;
    assign weights1[30][273] = 16'b1111111111111111;
    assign weights1[30][274] = 16'b1111111111011100;
    assign weights1[30][275] = 16'b1111111111011001;
    assign weights1[30][276] = 16'b1111111111100111;
    assign weights1[30][277] = 16'b1111111111110010;
    assign weights1[30][278] = 16'b1111111111110011;
    assign weights1[30][279] = 16'b1111111111111010;
    assign weights1[30][280] = 16'b0000000000000110;
    assign weights1[30][281] = 16'b0000000000000100;
    assign weights1[30][282] = 16'b1111111111110101;
    assign weights1[30][283] = 16'b1111111111111110;
    assign weights1[30][284] = 16'b0000000000010111;
    assign weights1[30][285] = 16'b0000000000011101;
    assign weights1[30][286] = 16'b0000000000001100;
    assign weights1[30][287] = 16'b1111111111110000;
    assign weights1[30][288] = 16'b1111111111000100;
    assign weights1[30][289] = 16'b1111111101110010;
    assign weights1[30][290] = 16'b1111111100011001;
    assign weights1[30][291] = 16'b1111111011111010;
    assign weights1[30][292] = 16'b1111111110100000;
    assign weights1[30][293] = 16'b1111111111011001;
    assign weights1[30][294] = 16'b1111111111111100;
    assign weights1[30][295] = 16'b0000000000001111;
    assign weights1[30][296] = 16'b0000000000010100;
    assign weights1[30][297] = 16'b0000000000011101;
    assign weights1[30][298] = 16'b0000000000000001;
    assign weights1[30][299] = 16'b1111111111101111;
    assign weights1[30][300] = 16'b1111111111100111;
    assign weights1[30][301] = 16'b1111111111011110;
    assign weights1[30][302] = 16'b1111111111011001;
    assign weights1[30][303] = 16'b1111111111100010;
    assign weights1[30][304] = 16'b1111111111110001;
    assign weights1[30][305] = 16'b1111111111110000;
    assign weights1[30][306] = 16'b1111111111111010;
    assign weights1[30][307] = 16'b1111111111110110;
    assign weights1[30][308] = 16'b1111111111111110;
    assign weights1[30][309] = 16'b1111111111110011;
    assign weights1[30][310] = 16'b1111111111101100;
    assign weights1[30][311] = 16'b1111111111100111;
    assign weights1[30][312] = 16'b1111111111111100;
    assign weights1[30][313] = 16'b1111111111100011;
    assign weights1[30][314] = 16'b1111111110111001;
    assign weights1[30][315] = 16'b1111111101100111;
    assign weights1[30][316] = 16'b1111111100011001;
    assign weights1[30][317] = 16'b1111111011011001;
    assign weights1[30][318] = 16'b1111111101011100;
    assign weights1[30][319] = 16'b1111111111100101;
    assign weights1[30][320] = 16'b1111111111101100;
    assign weights1[30][321] = 16'b0000000000000111;
    assign weights1[30][322] = 16'b0000000000011010;
    assign weights1[30][323] = 16'b0000000000010110;
    assign weights1[30][324] = 16'b0000000000011000;
    assign weights1[30][325] = 16'b1111111111111111;
    assign weights1[30][326] = 16'b0000000000001110;
    assign weights1[30][327] = 16'b1111111111110010;
    assign weights1[30][328] = 16'b1111111111111010;
    assign weights1[30][329] = 16'b1111111111011010;
    assign weights1[30][330] = 16'b1111111111011011;
    assign weights1[30][331] = 16'b1111111111110011;
    assign weights1[30][332] = 16'b1111111111110101;
    assign weights1[30][333] = 16'b1111111111111011;
    assign weights1[30][334] = 16'b1111111111111011;
    assign weights1[30][335] = 16'b1111111111111000;
    assign weights1[30][336] = 16'b1111111111110011;
    assign weights1[30][337] = 16'b1111111111100011;
    assign weights1[30][338] = 16'b1111111111010100;
    assign weights1[30][339] = 16'b1111111111000000;
    assign weights1[30][340] = 16'b1111111110101101;
    assign weights1[30][341] = 16'b1111111110011000;
    assign weights1[30][342] = 16'b1111111101101101;
    assign weights1[30][343] = 16'b1111111100110110;
    assign weights1[30][344] = 16'b1111111100110010;
    assign weights1[30][345] = 16'b1111111110111010;
    assign weights1[30][346] = 16'b0000000000001000;
    assign weights1[30][347] = 16'b0000000000100001;
    assign weights1[30][348] = 16'b0000000000010011;
    assign weights1[30][349] = 16'b0000000000001001;
    assign weights1[30][350] = 16'b0000000000010010;
    assign weights1[30][351] = 16'b0000000000001010;
    assign weights1[30][352] = 16'b0000000000011010;
    assign weights1[30][353] = 16'b0000000000010100;
    assign weights1[30][354] = 16'b0000000000001011;
    assign weights1[30][355] = 16'b1111111111101111;
    assign weights1[30][356] = 16'b1111111111011011;
    assign weights1[30][357] = 16'b1111111111101010;
    assign weights1[30][358] = 16'b1111111111101100;
    assign weights1[30][359] = 16'b1111111111111110;
    assign weights1[30][360] = 16'b1111111111111010;
    assign weights1[30][361] = 16'b1111111111111010;
    assign weights1[30][362] = 16'b1111111111111001;
    assign weights1[30][363] = 16'b0000000000000011;
    assign weights1[30][364] = 16'b1111111111100010;
    assign weights1[30][365] = 16'b1111111111010111;
    assign weights1[30][366] = 16'b1111111111000011;
    assign weights1[30][367] = 16'b1111111110101001;
    assign weights1[30][368] = 16'b1111111110100101;
    assign weights1[30][369] = 16'b1111111110000110;
    assign weights1[30][370] = 16'b1111111101101101;
    assign weights1[30][371] = 16'b1111111110001110;
    assign weights1[30][372] = 16'b1111111111000101;
    assign weights1[30][373] = 16'b0000000000000110;
    assign weights1[30][374] = 16'b0000000000101010;
    assign weights1[30][375] = 16'b0000000000011011;
    assign weights1[30][376] = 16'b0000000000010100;
    assign weights1[30][377] = 16'b0000000000001000;
    assign weights1[30][378] = 16'b0000000000100101;
    assign weights1[30][379] = 16'b0000000000001011;
    assign weights1[30][380] = 16'b0000000000000001;
    assign weights1[30][381] = 16'b0000000000001110;
    assign weights1[30][382] = 16'b0000000000000100;
    assign weights1[30][383] = 16'b1111111111101111;
    assign weights1[30][384] = 16'b1111111111101111;
    assign weights1[30][385] = 16'b1111111111111111;
    assign weights1[30][386] = 16'b1111111111110110;
    assign weights1[30][387] = 16'b1111111111111100;
    assign weights1[30][388] = 16'b1111111111110111;
    assign weights1[30][389] = 16'b1111111111111011;
    assign weights1[30][390] = 16'b0000000000000011;
    assign weights1[30][391] = 16'b0000000000000010;
    assign weights1[30][392] = 16'b1111111111100101;
    assign weights1[30][393] = 16'b1111111111001110;
    assign weights1[30][394] = 16'b1111111110110111;
    assign weights1[30][395] = 16'b1111111110100100;
    assign weights1[30][396] = 16'b1111111110100011;
    assign weights1[30][397] = 16'b1111111110000111;
    assign weights1[30][398] = 16'b1111111110101000;
    assign weights1[30][399] = 16'b1111111111101000;
    assign weights1[30][400] = 16'b0000000000100000;
    assign weights1[30][401] = 16'b1111111111110111;
    assign weights1[30][402] = 16'b0000000000000100;
    assign weights1[30][403] = 16'b0000000000000011;
    assign weights1[30][404] = 16'b0000000000001000;
    assign weights1[30][405] = 16'b0000000000000101;
    assign weights1[30][406] = 16'b0000000000010001;
    assign weights1[30][407] = 16'b0000000000010101;
    assign weights1[30][408] = 16'b0000000000000100;
    assign weights1[30][409] = 16'b0000000000001000;
    assign weights1[30][410] = 16'b1111111111110000;
    assign weights1[30][411] = 16'b1111111111111000;
    assign weights1[30][412] = 16'b1111111111111111;
    assign weights1[30][413] = 16'b1111111111111010;
    assign weights1[30][414] = 16'b1111111111110011;
    assign weights1[30][415] = 16'b1111111111111001;
    assign weights1[30][416] = 16'b0000000000000010;
    assign weights1[30][417] = 16'b0000000000000011;
    assign weights1[30][418] = 16'b0000000000001011;
    assign weights1[30][419] = 16'b0000000000000110;
    assign weights1[30][420] = 16'b1111111111100010;
    assign weights1[30][421] = 16'b1111111111001100;
    assign weights1[30][422] = 16'b1111111110111101;
    assign weights1[30][423] = 16'b1111111110111010;
    assign weights1[30][424] = 16'b1111111110110010;
    assign weights1[30][425] = 16'b1111111111011100;
    assign weights1[30][426] = 16'b1111111111111011;
    assign weights1[30][427] = 16'b1111111111110011;
    assign weights1[30][428] = 16'b1111111111100001;
    assign weights1[30][429] = 16'b0000000000010011;
    assign weights1[30][430] = 16'b1111111111110100;
    assign weights1[30][431] = 16'b0000000000000011;
    assign weights1[30][432] = 16'b1111111111111101;
    assign weights1[30][433] = 16'b1111111111111100;
    assign weights1[30][434] = 16'b0000000000001000;
    assign weights1[30][435] = 16'b0000000000000010;
    assign weights1[30][436] = 16'b1111111111110101;
    assign weights1[30][437] = 16'b1111111111111000;
    assign weights1[30][438] = 16'b1111111111101111;
    assign weights1[30][439] = 16'b1111111111101101;
    assign weights1[30][440] = 16'b1111111111101101;
    assign weights1[30][441] = 16'b1111111111111011;
    assign weights1[30][442] = 16'b0000000000001000;
    assign weights1[30][443] = 16'b0000000000000101;
    assign weights1[30][444] = 16'b1111111111111000;
    assign weights1[30][445] = 16'b0000000000001000;
    assign weights1[30][446] = 16'b0000000000000000;
    assign weights1[30][447] = 16'b0000000000000001;
    assign weights1[30][448] = 16'b1111111111101011;
    assign weights1[30][449] = 16'b1111111111010101;
    assign weights1[30][450] = 16'b1111111111010011;
    assign weights1[30][451] = 16'b1111111111011101;
    assign weights1[30][452] = 16'b1111111111100110;
    assign weights1[30][453] = 16'b1111111111101111;
    assign weights1[30][454] = 16'b1111111111111110;
    assign weights1[30][455] = 16'b1111111111110110;
    assign weights1[30][456] = 16'b0000000000000001;
    assign weights1[30][457] = 16'b0000000000010000;
    assign weights1[30][458] = 16'b1111111111110100;
    assign weights1[30][459] = 16'b1111111111111100;
    assign weights1[30][460] = 16'b0000000000000000;
    assign weights1[30][461] = 16'b0000000000000101;
    assign weights1[30][462] = 16'b0000000000000010;
    assign weights1[30][463] = 16'b1111111111101000;
    assign weights1[30][464] = 16'b1111111111111101;
    assign weights1[30][465] = 16'b1111111111110110;
    assign weights1[30][466] = 16'b0000000000000111;
    assign weights1[30][467] = 16'b0000000000011110;
    assign weights1[30][468] = 16'b1111111111111100;
    assign weights1[30][469] = 16'b0000000000000010;
    assign weights1[30][470] = 16'b1111111111111111;
    assign weights1[30][471] = 16'b1111111111111000;
    assign weights1[30][472] = 16'b0000000000010011;
    assign weights1[30][473] = 16'b0000000000010001;
    assign weights1[30][474] = 16'b0000000000001110;
    assign weights1[30][475] = 16'b0000000000000101;
    assign weights1[30][476] = 16'b1111111111111000;
    assign weights1[30][477] = 16'b1111111111100011;
    assign weights1[30][478] = 16'b1111111111101110;
    assign weights1[30][479] = 16'b1111111111101000;
    assign weights1[30][480] = 16'b1111111111101110;
    assign weights1[30][481] = 16'b1111111111110101;
    assign weights1[30][482] = 16'b1111111111100000;
    assign weights1[30][483] = 16'b1111111111110101;
    assign weights1[30][484] = 16'b1111111111101011;
    assign weights1[30][485] = 16'b1111111111100011;
    assign weights1[30][486] = 16'b1111111111010010;
    assign weights1[30][487] = 16'b1111111111111001;
    assign weights1[30][488] = 16'b1111111111101011;
    assign weights1[30][489] = 16'b1111111111111001;
    assign weights1[30][490] = 16'b1111111111111100;
    assign weights1[30][491] = 16'b1111111111111011;
    assign weights1[30][492] = 16'b1111111111110000;
    assign weights1[30][493] = 16'b1111111111110010;
    assign weights1[30][494] = 16'b1111111111101101;
    assign weights1[30][495] = 16'b0000000000000001;
    assign weights1[30][496] = 16'b0000000000000110;
    assign weights1[30][497] = 16'b0000000000000011;
    assign weights1[30][498] = 16'b0000000000001011;
    assign weights1[30][499] = 16'b0000000000011011;
    assign weights1[30][500] = 16'b0000000000001111;
    assign weights1[30][501] = 16'b0000000000000011;
    assign weights1[30][502] = 16'b0000000000000001;
    assign weights1[30][503] = 16'b1111111111111100;
    assign weights1[30][504] = 16'b1111111111111111;
    assign weights1[30][505] = 16'b1111111111111101;
    assign weights1[30][506] = 16'b1111111111110110;
    assign weights1[30][507] = 16'b1111111111110110;
    assign weights1[30][508] = 16'b1111111111101001;
    assign weights1[30][509] = 16'b0000000000000101;
    assign weights1[30][510] = 16'b1111111111100110;
    assign weights1[30][511] = 16'b1111111111111000;
    assign weights1[30][512] = 16'b1111111111011000;
    assign weights1[30][513] = 16'b1111111111110011;
    assign weights1[30][514] = 16'b1111111111010110;
    assign weights1[30][515] = 16'b1111111111001110;
    assign weights1[30][516] = 16'b1111111111001111;
    assign weights1[30][517] = 16'b1111111111111011;
    assign weights1[30][518] = 16'b1111111111110111;
    assign weights1[30][519] = 16'b1111111111110010;
    assign weights1[30][520] = 16'b1111111111100011;
    assign weights1[30][521] = 16'b1111111111111111;
    assign weights1[30][522] = 16'b1111111111101111;
    assign weights1[30][523] = 16'b0000000000001000;
    assign weights1[30][524] = 16'b1111111111101000;
    assign weights1[30][525] = 16'b0000000000001111;
    assign weights1[30][526] = 16'b1111111111110000;
    assign weights1[30][527] = 16'b1111111111110101;
    assign weights1[30][528] = 16'b1111111111110111;
    assign weights1[30][529] = 16'b0000000000010101;
    assign weights1[30][530] = 16'b0000000000001100;
    assign weights1[30][531] = 16'b0000000000001000;
    assign weights1[30][532] = 16'b0000000000010000;
    assign weights1[30][533] = 16'b0000000000000001;
    assign weights1[30][534] = 16'b0000000000000100;
    assign weights1[30][535] = 16'b0000000000011110;
    assign weights1[30][536] = 16'b1111111111011001;
    assign weights1[30][537] = 16'b1111111111111001;
    assign weights1[30][538] = 16'b0000000000001000;
    assign weights1[30][539] = 16'b1111111111110111;
    assign weights1[30][540] = 16'b1111111111101100;
    assign weights1[30][541] = 16'b1111111111111101;
    assign weights1[30][542] = 16'b1111111111110100;
    assign weights1[30][543] = 16'b1111111111110000;
    assign weights1[30][544] = 16'b0000000000000100;
    assign weights1[30][545] = 16'b0000000000000000;
    assign weights1[30][546] = 16'b1111111111111100;
    assign weights1[30][547] = 16'b1111111111110100;
    assign weights1[30][548] = 16'b0000000000001011;
    assign weights1[30][549] = 16'b1111111111011111;
    assign weights1[30][550] = 16'b1111111111101111;
    assign weights1[30][551] = 16'b1111111111100111;
    assign weights1[30][552] = 16'b1111111111101111;
    assign weights1[30][553] = 16'b0000000000001100;
    assign weights1[30][554] = 16'b0000000000000001;
    assign weights1[30][555] = 16'b1111111111111111;
    assign weights1[30][556] = 16'b1111111111111111;
    assign weights1[30][557] = 16'b0000000000010000;
    assign weights1[30][558] = 16'b0000000000000100;
    assign weights1[30][559] = 16'b0000000000001111;
    assign weights1[30][560] = 16'b0000000000010100;
    assign weights1[30][561] = 16'b0000000000001100;
    assign weights1[30][562] = 16'b0000000000001001;
    assign weights1[30][563] = 16'b0000000000010110;
    assign weights1[30][564] = 16'b0000000000001101;
    assign weights1[30][565] = 16'b1111111111101001;
    assign weights1[30][566] = 16'b0000000000001011;
    assign weights1[30][567] = 16'b1111111111111111;
    assign weights1[30][568] = 16'b1111111111111100;
    assign weights1[30][569] = 16'b0000000000001011;
    assign weights1[30][570] = 16'b1111111111110101;
    assign weights1[30][571] = 16'b1111111111111101;
    assign weights1[30][572] = 16'b0000000000001111;
    assign weights1[30][573] = 16'b1111111111111101;
    assign weights1[30][574] = 16'b0000000000001000;
    assign weights1[30][575] = 16'b1111111111110110;
    assign weights1[30][576] = 16'b1111111111110111;
    assign weights1[30][577] = 16'b1111111111101101;
    assign weights1[30][578] = 16'b0000000000010011;
    assign weights1[30][579] = 16'b0000000000000100;
    assign weights1[30][580] = 16'b1111111111110001;
    assign weights1[30][581] = 16'b0000000000010100;
    assign weights1[30][582] = 16'b1111111111111010;
    assign weights1[30][583] = 16'b1111111111111000;
    assign weights1[30][584] = 16'b0000000000000110;
    assign weights1[30][585] = 16'b0000000000001000;
    assign weights1[30][586] = 16'b0000000000000111;
    assign weights1[30][587] = 16'b0000000000000110;
    assign weights1[30][588] = 16'b0000000000010100;
    assign weights1[30][589] = 16'b0000000000001010;
    assign weights1[30][590] = 16'b0000000000000000;
    assign weights1[30][591] = 16'b0000000000011000;
    assign weights1[30][592] = 16'b0000000000001011;
    assign weights1[30][593] = 16'b1111111111111100;
    assign weights1[30][594] = 16'b0000000000001011;
    assign weights1[30][595] = 16'b1111111111100001;
    assign weights1[30][596] = 16'b0000000000001100;
    assign weights1[30][597] = 16'b1111111111100111;
    assign weights1[30][598] = 16'b0000000000001000;
    assign weights1[30][599] = 16'b0000000000000000;
    assign weights1[30][600] = 16'b1111111111101101;
    assign weights1[30][601] = 16'b0000000000000101;
    assign weights1[30][602] = 16'b0000000000010010;
    assign weights1[30][603] = 16'b1111111111101110;
    assign weights1[30][604] = 16'b0000000000010100;
    assign weights1[30][605] = 16'b1111111111111111;
    assign weights1[30][606] = 16'b1111111111100111;
    assign weights1[30][607] = 16'b1111111111101010;
    assign weights1[30][608] = 16'b0000000000000101;
    assign weights1[30][609] = 16'b1111111111101111;
    assign weights1[30][610] = 16'b1111111111100111;
    assign weights1[30][611] = 16'b0000000000001100;
    assign weights1[30][612] = 16'b0000000000010010;
    assign weights1[30][613] = 16'b1111111111110100;
    assign weights1[30][614] = 16'b1111111111111100;
    assign weights1[30][615] = 16'b0000000000000100;
    assign weights1[30][616] = 16'b0000000000000101;
    assign weights1[30][617] = 16'b0000000000001111;
    assign weights1[30][618] = 16'b0000000000000111;
    assign weights1[30][619] = 16'b0000000000000000;
    assign weights1[30][620] = 16'b0000000000010100;
    assign weights1[30][621] = 16'b0000000000010000;
    assign weights1[30][622] = 16'b0000000000010010;
    assign weights1[30][623] = 16'b0000000000010111;
    assign weights1[30][624] = 16'b1111111111111000;
    assign weights1[30][625] = 16'b0000000000100110;
    assign weights1[30][626] = 16'b0000000000000001;
    assign weights1[30][627] = 16'b1111111111111011;
    assign weights1[30][628] = 16'b1111111111110000;
    assign weights1[30][629] = 16'b1111111111111001;
    assign weights1[30][630] = 16'b0000000000010100;
    assign weights1[30][631] = 16'b0000000000001011;
    assign weights1[30][632] = 16'b0000000000000001;
    assign weights1[30][633] = 16'b1111111111111110;
    assign weights1[30][634] = 16'b1111111111111000;
    assign weights1[30][635] = 16'b1111111111111010;
    assign weights1[30][636] = 16'b1111111111011011;
    assign weights1[30][637] = 16'b1111111111100110;
    assign weights1[30][638] = 16'b1111111111100111;
    assign weights1[30][639] = 16'b1111111111101110;
    assign weights1[30][640] = 16'b1111111111111010;
    assign weights1[30][641] = 16'b1111111111101100;
    assign weights1[30][642] = 16'b1111111111111101;
    assign weights1[30][643] = 16'b1111111111111100;
    assign weights1[30][644] = 16'b0000000000001000;
    assign weights1[30][645] = 16'b0000000000001101;
    assign weights1[30][646] = 16'b0000000000001101;
    assign weights1[30][647] = 16'b0000000000001001;
    assign weights1[30][648] = 16'b1111111111111111;
    assign weights1[30][649] = 16'b0000000000000111;
    assign weights1[30][650] = 16'b1111111111111010;
    assign weights1[30][651] = 16'b0000000000010001;
    assign weights1[30][652] = 16'b0000000000011010;
    assign weights1[30][653] = 16'b0000000000000111;
    assign weights1[30][654] = 16'b1111111111111000;
    assign weights1[30][655] = 16'b0000000000001100;
    assign weights1[30][656] = 16'b0000000000001010;
    assign weights1[30][657] = 16'b1111111111111100;
    assign weights1[30][658] = 16'b1111111111111110;
    assign weights1[30][659] = 16'b1111111111111100;
    assign weights1[30][660] = 16'b0000000000000000;
    assign weights1[30][661] = 16'b0000000000000010;
    assign weights1[30][662] = 16'b1111111111111010;
    assign weights1[30][663] = 16'b1111111111110101;
    assign weights1[30][664] = 16'b0000000000000000;
    assign weights1[30][665] = 16'b1111111111011011;
    assign weights1[30][666] = 16'b1111111111101101;
    assign weights1[30][667] = 16'b1111111111110111;
    assign weights1[30][668] = 16'b1111111111110110;
    assign weights1[30][669] = 16'b1111111111110110;
    assign weights1[30][670] = 16'b1111111111111111;
    assign weights1[30][671] = 16'b1111111111111100;
    assign weights1[30][672] = 16'b0000000000001000;
    assign weights1[30][673] = 16'b0000000000010010;
    assign weights1[30][674] = 16'b0000000000001011;
    assign weights1[30][675] = 16'b0000000000010010;
    assign weights1[30][676] = 16'b0000000000001001;
    assign weights1[30][677] = 16'b0000000000000001;
    assign weights1[30][678] = 16'b0000000000000001;
    assign weights1[30][679] = 16'b0000000000010011;
    assign weights1[30][680] = 16'b0000000000000011;
    assign weights1[30][681] = 16'b0000000000001110;
    assign weights1[30][682] = 16'b1111111111111001;
    assign weights1[30][683] = 16'b0000000000000010;
    assign weights1[30][684] = 16'b1111111111110000;
    assign weights1[30][685] = 16'b1111111111101111;
    assign weights1[30][686] = 16'b0000000000001000;
    assign weights1[30][687] = 16'b1111111111110001;
    assign weights1[30][688] = 16'b1111111111100010;
    assign weights1[30][689] = 16'b1111111111111010;
    assign weights1[30][690] = 16'b1111111111111000;
    assign weights1[30][691] = 16'b1111111111110110;
    assign weights1[30][692] = 16'b1111111111110001;
    assign weights1[30][693] = 16'b1111111111110100;
    assign weights1[30][694] = 16'b1111111111110010;
    assign weights1[30][695] = 16'b1111111111110011;
    assign weights1[30][696] = 16'b1111111111110001;
    assign weights1[30][697] = 16'b0000000000000001;
    assign weights1[30][698] = 16'b1111111111111100;
    assign weights1[30][699] = 16'b1111111111111011;
    assign weights1[30][700] = 16'b0000000000001010;
    assign weights1[30][701] = 16'b0000000000001111;
    assign weights1[30][702] = 16'b0000000000010000;
    assign weights1[30][703] = 16'b1111111111111101;
    assign weights1[30][704] = 16'b0000000000000100;
    assign weights1[30][705] = 16'b0000000000001011;
    assign weights1[30][706] = 16'b0000000000010101;
    assign weights1[30][707] = 16'b0000000000001011;
    assign weights1[30][708] = 16'b1111111111111110;
    assign weights1[30][709] = 16'b1111111111101100;
    assign weights1[30][710] = 16'b1111111111111100;
    assign weights1[30][711] = 16'b1111111111111100;
    assign weights1[30][712] = 16'b0000000000001010;
    assign weights1[30][713] = 16'b1111111111110111;
    assign weights1[30][714] = 16'b1111111111111011;
    assign weights1[30][715] = 16'b1111111111100001;
    assign weights1[30][716] = 16'b0000000000010010;
    assign weights1[30][717] = 16'b0000000000001110;
    assign weights1[30][718] = 16'b0000000000001000;
    assign weights1[30][719] = 16'b0000000000000001;
    assign weights1[30][720] = 16'b0000000000001110;
    assign weights1[30][721] = 16'b1111111111111100;
    assign weights1[30][722] = 16'b0000000000000100;
    assign weights1[30][723] = 16'b1111111111111001;
    assign weights1[30][724] = 16'b1111111111111100;
    assign weights1[30][725] = 16'b0000000000000010;
    assign weights1[30][726] = 16'b1111111111111101;
    assign weights1[30][727] = 16'b1111111111111100;
    assign weights1[30][728] = 16'b0000000000000011;
    assign weights1[30][729] = 16'b0000000000001001;
    assign weights1[30][730] = 16'b0000000000010010;
    assign weights1[30][731] = 16'b0000000000001010;
    assign weights1[30][732] = 16'b1111111111110111;
    assign weights1[30][733] = 16'b1111111111110111;
    assign weights1[30][734] = 16'b0000000000001111;
    assign weights1[30][735] = 16'b0000000000010011;
    assign weights1[30][736] = 16'b1111111111110010;
    assign weights1[30][737] = 16'b1111111111100110;
    assign weights1[30][738] = 16'b1111111111111100;
    assign weights1[30][739] = 16'b1111111111111000;
    assign weights1[30][740] = 16'b1111111111110101;
    assign weights1[30][741] = 16'b0000000000000111;
    assign weights1[30][742] = 16'b0000000000000101;
    assign weights1[30][743] = 16'b0000000000001110;
    assign weights1[30][744] = 16'b0000000000000001;
    assign weights1[30][745] = 16'b1111111111111110;
    assign weights1[30][746] = 16'b0000000000000111;
    assign weights1[30][747] = 16'b0000000000000110;
    assign weights1[30][748] = 16'b0000000000001010;
    assign weights1[30][749] = 16'b0000000000000100;
    assign weights1[30][750] = 16'b0000000000000000;
    assign weights1[30][751] = 16'b1111111111111011;
    assign weights1[30][752] = 16'b1111111111111101;
    assign weights1[30][753] = 16'b0000000000000001;
    assign weights1[30][754] = 16'b1111111111111111;
    assign weights1[30][755] = 16'b1111111111111111;
    assign weights1[30][756] = 16'b0000000000000010;
    assign weights1[30][757] = 16'b0000000000000111;
    assign weights1[30][758] = 16'b0000000000001011;
    assign weights1[30][759] = 16'b0000000000011000;
    assign weights1[30][760] = 16'b0000000000010100;
    assign weights1[30][761] = 16'b0000000000011010;
    assign weights1[30][762] = 16'b0000000000100000;
    assign weights1[30][763] = 16'b0000000000010110;
    assign weights1[30][764] = 16'b0000000000010010;
    assign weights1[30][765] = 16'b0000000000001100;
    assign weights1[30][766] = 16'b0000000000000111;
    assign weights1[30][767] = 16'b0000000000000110;
    assign weights1[30][768] = 16'b0000000000001100;
    assign weights1[30][769] = 16'b0000000000000011;
    assign weights1[30][770] = 16'b1111111111110011;
    assign weights1[30][771] = 16'b0000000000001101;
    assign weights1[30][772] = 16'b0000000000010011;
    assign weights1[30][773] = 16'b1111111111111001;
    assign weights1[30][774] = 16'b1111111111111010;
    assign weights1[30][775] = 16'b0000000000010101;
    assign weights1[30][776] = 16'b0000000000001110;
    assign weights1[30][777] = 16'b0000000000000001;
    assign weights1[30][778] = 16'b1111111111111110;
    assign weights1[30][779] = 16'b0000000000000011;
    assign weights1[30][780] = 16'b0000000000000001;
    assign weights1[30][781] = 16'b0000000000000001;
    assign weights1[30][782] = 16'b0000000000000001;
    assign weights1[30][783] = 16'b0000000000000000;
    assign weights1[31][0] = 16'b0000000000000001;
    assign weights1[31][1] = 16'b0000000000000001;
    assign weights1[31][2] = 16'b0000000000000000;
    assign weights1[31][3] = 16'b1111111111111100;
    assign weights1[31][4] = 16'b0000000000000000;
    assign weights1[31][5] = 16'b1111111111111000;
    assign weights1[31][6] = 16'b1111111111110111;
    assign weights1[31][7] = 16'b1111111111111000;
    assign weights1[31][8] = 16'b1111111111111000;
    assign weights1[31][9] = 16'b1111111111110111;
    assign weights1[31][10] = 16'b1111111111111010;
    assign weights1[31][11] = 16'b0000000000000011;
    assign weights1[31][12] = 16'b1111111111111110;
    assign weights1[31][13] = 16'b1111111111110101;
    assign weights1[31][14] = 16'b1111111111111000;
    assign weights1[31][15] = 16'b1111111111101001;
    assign weights1[31][16] = 16'b1111111111110011;
    assign weights1[31][17] = 16'b1111111111110101;
    assign weights1[31][18] = 16'b1111111111111101;
    assign weights1[31][19] = 16'b1111111111101011;
    assign weights1[31][20] = 16'b1111111111110011;
    assign weights1[31][21] = 16'b1111111111111001;
    assign weights1[31][22] = 16'b1111111111111110;
    assign weights1[31][23] = 16'b0000000000000101;
    assign weights1[31][24] = 16'b0000000000000110;
    assign weights1[31][25] = 16'b0000000000000100;
    assign weights1[31][26] = 16'b0000000000000101;
    assign weights1[31][27] = 16'b0000000000000001;
    assign weights1[31][28] = 16'b0000000000000000;
    assign weights1[31][29] = 16'b1111111111111111;
    assign weights1[31][30] = 16'b1111111111111011;
    assign weights1[31][31] = 16'b1111111111111100;
    assign weights1[31][32] = 16'b1111111111111011;
    assign weights1[31][33] = 16'b1111111111110111;
    assign weights1[31][34] = 16'b1111111111110000;
    assign weights1[31][35] = 16'b1111111111101011;
    assign weights1[31][36] = 16'b1111111111111100;
    assign weights1[31][37] = 16'b1111111111111010;
    assign weights1[31][38] = 16'b0000000000000001;
    assign weights1[31][39] = 16'b0000000000001001;
    assign weights1[31][40] = 16'b1111111111111000;
    assign weights1[31][41] = 16'b1111111111111111;
    assign weights1[31][42] = 16'b1111111111111011;
    assign weights1[31][43] = 16'b1111111111110110;
    assign weights1[31][44] = 16'b1111111111110110;
    assign weights1[31][45] = 16'b1111111111111000;
    assign weights1[31][46] = 16'b1111111111111010;
    assign weights1[31][47] = 16'b1111111111110100;
    assign weights1[31][48] = 16'b0000000000000000;
    assign weights1[31][49] = 16'b0000000000000011;
    assign weights1[31][50] = 16'b0000000000000111;
    assign weights1[31][51] = 16'b0000000000000000;
    assign weights1[31][52] = 16'b1111111111111111;
    assign weights1[31][53] = 16'b0000000000000101;
    assign weights1[31][54] = 16'b0000000000000011;
    assign weights1[31][55] = 16'b0000000000000011;
    assign weights1[31][56] = 16'b0000000000000000;
    assign weights1[31][57] = 16'b1111111111111111;
    assign weights1[31][58] = 16'b1111111111110111;
    assign weights1[31][59] = 16'b1111111111111100;
    assign weights1[31][60] = 16'b1111111111111011;
    assign weights1[31][61] = 16'b1111111111110011;
    assign weights1[31][62] = 16'b1111111111110110;
    assign weights1[31][63] = 16'b1111111111101101;
    assign weights1[31][64] = 16'b1111111111111000;
    assign weights1[31][65] = 16'b1111111111111000;
    assign weights1[31][66] = 16'b0000000000000011;
    assign weights1[31][67] = 16'b1111111111111100;
    assign weights1[31][68] = 16'b1111111111111001;
    assign weights1[31][69] = 16'b0000000000000010;
    assign weights1[31][70] = 16'b0000000000000100;
    assign weights1[31][71] = 16'b1111111111111001;
    assign weights1[31][72] = 16'b1111111111110010;
    assign weights1[31][73] = 16'b1111111111111010;
    assign weights1[31][74] = 16'b1111111111110111;
    assign weights1[31][75] = 16'b1111111111110011;
    assign weights1[31][76] = 16'b1111111111111101;
    assign weights1[31][77] = 16'b0000000000000100;
    assign weights1[31][78] = 16'b0000000000001100;
    assign weights1[31][79] = 16'b0000000000000001;
    assign weights1[31][80] = 16'b1111111111111101;
    assign weights1[31][81] = 16'b1111111111111000;
    assign weights1[31][82] = 16'b0000000000000001;
    assign weights1[31][83] = 16'b1111111111111111;
    assign weights1[31][84] = 16'b0000000000000000;
    assign weights1[31][85] = 16'b1111111111111100;
    assign weights1[31][86] = 16'b1111111111111011;
    assign weights1[31][87] = 16'b1111111111111001;
    assign weights1[31][88] = 16'b1111111111111101;
    assign weights1[31][89] = 16'b1111111111111101;
    assign weights1[31][90] = 16'b0000000000000111;
    assign weights1[31][91] = 16'b1111111111110000;
    assign weights1[31][92] = 16'b0000000000001010;
    assign weights1[31][93] = 16'b1111111111101011;
    assign weights1[31][94] = 16'b1111111111110011;
    assign weights1[31][95] = 16'b1111111111110001;
    assign weights1[31][96] = 16'b0000000000000010;
    assign weights1[31][97] = 16'b1111111111110110;
    assign weights1[31][98] = 16'b0000000000001111;
    assign weights1[31][99] = 16'b0000000000001000;
    assign weights1[31][100] = 16'b0000000000000001;
    assign weights1[31][101] = 16'b1111111111110010;
    assign weights1[31][102] = 16'b1111111111111001;
    assign weights1[31][103] = 16'b1111111111111100;
    assign weights1[31][104] = 16'b0000000000001001;
    assign weights1[31][105] = 16'b0000000000010000;
    assign weights1[31][106] = 16'b1111111111111101;
    assign weights1[31][107] = 16'b1111111111111000;
    assign weights1[31][108] = 16'b0000000000001000;
    assign weights1[31][109] = 16'b0000000000000000;
    assign weights1[31][110] = 16'b0000000000000100;
    assign weights1[31][111] = 16'b1111111111111011;
    assign weights1[31][112] = 16'b1111111111111111;
    assign weights1[31][113] = 16'b1111111111111111;
    assign weights1[31][114] = 16'b0000000000000010;
    assign weights1[31][115] = 16'b1111111111111101;
    assign weights1[31][116] = 16'b1111111111111010;
    assign weights1[31][117] = 16'b1111111111110110;
    assign weights1[31][118] = 16'b0000000000001111;
    assign weights1[31][119] = 16'b1111111111101111;
    assign weights1[31][120] = 16'b0000000000001010;
    assign weights1[31][121] = 16'b1111111111111001;
    assign weights1[31][122] = 16'b1111111111111000;
    assign weights1[31][123] = 16'b1111111111111000;
    assign weights1[31][124] = 16'b0000000000000011;
    assign weights1[31][125] = 16'b1111111111110101;
    assign weights1[31][126] = 16'b0000000000000010;
    assign weights1[31][127] = 16'b0000000000000011;
    assign weights1[31][128] = 16'b1111111111111111;
    assign weights1[31][129] = 16'b0000000000010011;
    assign weights1[31][130] = 16'b1111111111111001;
    assign weights1[31][131] = 16'b1111111111101110;
    assign weights1[31][132] = 16'b1111111111111111;
    assign weights1[31][133] = 16'b0000000000001110;
    assign weights1[31][134] = 16'b1111111111110111;
    assign weights1[31][135] = 16'b0000000000000001;
    assign weights1[31][136] = 16'b0000000000010011;
    assign weights1[31][137] = 16'b0000000000010101;
    assign weights1[31][138] = 16'b1111111111111101;
    assign weights1[31][139] = 16'b0000000000000111;
    assign weights1[31][140] = 16'b1111111111111101;
    assign weights1[31][141] = 16'b0000000000000010;
    assign weights1[31][142] = 16'b0000000000000101;
    assign weights1[31][143] = 16'b1111111111110111;
    assign weights1[31][144] = 16'b1111111111111110;
    assign weights1[31][145] = 16'b1111111111111011;
    assign weights1[31][146] = 16'b1111111111110101;
    assign weights1[31][147] = 16'b0000000000001001;
    assign weights1[31][148] = 16'b1111111111111111;
    assign weights1[31][149] = 16'b0000000000001010;
    assign weights1[31][150] = 16'b0000000000000111;
    assign weights1[31][151] = 16'b0000000000000100;
    assign weights1[31][152] = 16'b0000000000001100;
    assign weights1[31][153] = 16'b1111111111111101;
    assign weights1[31][154] = 16'b0000000000000010;
    assign weights1[31][155] = 16'b1111111111111111;
    assign weights1[31][156] = 16'b0000000000000000;
    assign weights1[31][157] = 16'b0000000000000010;
    assign weights1[31][158] = 16'b1111111111110000;
    assign weights1[31][159] = 16'b1111111111111011;
    assign weights1[31][160] = 16'b0000000000000001;
    assign weights1[31][161] = 16'b0000000000000011;
    assign weights1[31][162] = 16'b0000000000000111;
    assign weights1[31][163] = 16'b0000000000000011;
    assign weights1[31][164] = 16'b0000000000001011;
    assign weights1[31][165] = 16'b1111111111110101;
    assign weights1[31][166] = 16'b1111111111111011;
    assign weights1[31][167] = 16'b1111111111111010;
    assign weights1[31][168] = 16'b0000000000000010;
    assign weights1[31][169] = 16'b0000000000000001;
    assign weights1[31][170] = 16'b1111111111111010;
    assign weights1[31][171] = 16'b1111111111111101;
    assign weights1[31][172] = 16'b0000000000001011;
    assign weights1[31][173] = 16'b0000000000000101;
    assign weights1[31][174] = 16'b1111111111111101;
    assign weights1[31][175] = 16'b1111111111011110;
    assign weights1[31][176] = 16'b1111111111111101;
    assign weights1[31][177] = 16'b1111111111110101;
    assign weights1[31][178] = 16'b1111111111111100;
    assign weights1[31][179] = 16'b1111111111100000;
    assign weights1[31][180] = 16'b0000000000000101;
    assign weights1[31][181] = 16'b0000000000000111;
    assign weights1[31][182] = 16'b0000000000000011;
    assign weights1[31][183] = 16'b0000000000001010;
    assign weights1[31][184] = 16'b1111111111111111;
    assign weights1[31][185] = 16'b1111111111110000;
    assign weights1[31][186] = 16'b1111111111111000;
    assign weights1[31][187] = 16'b1111111111110010;
    assign weights1[31][188] = 16'b1111111111110000;
    assign weights1[31][189] = 16'b0000000000000111;
    assign weights1[31][190] = 16'b1111111111101101;
    assign weights1[31][191] = 16'b1111111111111100;
    assign weights1[31][192] = 16'b0000000000001011;
    assign weights1[31][193] = 16'b0000000000001011;
    assign weights1[31][194] = 16'b0000000000000100;
    assign weights1[31][195] = 16'b1111111111111110;
    assign weights1[31][196] = 16'b0000000000000000;
    assign weights1[31][197] = 16'b0000000000000111;
    assign weights1[31][198] = 16'b0000000000000100;
    assign weights1[31][199] = 16'b0000000000000111;
    assign weights1[31][200] = 16'b1111111111111110;
    assign weights1[31][201] = 16'b0000000000000101;
    assign weights1[31][202] = 16'b0000000000001011;
    assign weights1[31][203] = 16'b0000000000000110;
    assign weights1[31][204] = 16'b1111111111110001;
    assign weights1[31][205] = 16'b0000000000000100;
    assign weights1[31][206] = 16'b1111111111110111;
    assign weights1[31][207] = 16'b0000000000001000;
    assign weights1[31][208] = 16'b1111111111110001;
    assign weights1[31][209] = 16'b1111111111110111;
    assign weights1[31][210] = 16'b1111111111110110;
    assign weights1[31][211] = 16'b1111111111110000;
    assign weights1[31][212] = 16'b1111111111110111;
    assign weights1[31][213] = 16'b1111111111111111;
    assign weights1[31][214] = 16'b1111111111111001;
    assign weights1[31][215] = 16'b0000000000000001;
    assign weights1[31][216] = 16'b1111111111110110;
    assign weights1[31][217] = 16'b0000000000001001;
    assign weights1[31][218] = 16'b1111111111111001;
    assign weights1[31][219] = 16'b0000000000010101;
    assign weights1[31][220] = 16'b0000000000000010;
    assign weights1[31][221] = 16'b1111111111111101;
    assign weights1[31][222] = 16'b1111111111111001;
    assign weights1[31][223] = 16'b1111111111111110;
    assign weights1[31][224] = 16'b0000000000001010;
    assign weights1[31][225] = 16'b0000000000000000;
    assign weights1[31][226] = 16'b0000000000001001;
    assign weights1[31][227] = 16'b0000000000001000;
    assign weights1[31][228] = 16'b0000000000001001;
    assign weights1[31][229] = 16'b0000000000000100;
    assign weights1[31][230] = 16'b0000000000001100;
    assign weights1[31][231] = 16'b0000000000000000;
    assign weights1[31][232] = 16'b0000000000010010;
    assign weights1[31][233] = 16'b1111111111111001;
    assign weights1[31][234] = 16'b0000000000000101;
    assign weights1[31][235] = 16'b1111111111111010;
    assign weights1[31][236] = 16'b0000000000001000;
    assign weights1[31][237] = 16'b1111111111111001;
    assign weights1[31][238] = 16'b0000000000001110;
    assign weights1[31][239] = 16'b1111111111111101;
    assign weights1[31][240] = 16'b1111111111111110;
    assign weights1[31][241] = 16'b0000000000010010;
    assign weights1[31][242] = 16'b1111111111110101;
    assign weights1[31][243] = 16'b1111111111111100;
    assign weights1[31][244] = 16'b1111111111111011;
    assign weights1[31][245] = 16'b0000000000001100;
    assign weights1[31][246] = 16'b1111111111110011;
    assign weights1[31][247] = 16'b1111111111110110;
    assign weights1[31][248] = 16'b0000000000000011;
    assign weights1[31][249] = 16'b0000000000001001;
    assign weights1[31][250] = 16'b1111111111110110;
    assign weights1[31][251] = 16'b1111111111110110;
    assign weights1[31][252] = 16'b0000000000000011;
    assign weights1[31][253] = 16'b0000000000000110;
    assign weights1[31][254] = 16'b0000000000001101;
    assign weights1[31][255] = 16'b1111111111111100;
    assign weights1[31][256] = 16'b0000000000001111;
    assign weights1[31][257] = 16'b0000000000001001;
    assign weights1[31][258] = 16'b1111111111111101;
    assign weights1[31][259] = 16'b0000000000001011;
    assign weights1[31][260] = 16'b1111111111111010;
    assign weights1[31][261] = 16'b0000000000000110;
    assign weights1[31][262] = 16'b0000000000001111;
    assign weights1[31][263] = 16'b1111111111111000;
    assign weights1[31][264] = 16'b1111111111110100;
    assign weights1[31][265] = 16'b1111111111110111;
    assign weights1[31][266] = 16'b0000000000000000;
    assign weights1[31][267] = 16'b0000000000000000;
    assign weights1[31][268] = 16'b1111111111111101;
    assign weights1[31][269] = 16'b1111111111111011;
    assign weights1[31][270] = 16'b0000000000000110;
    assign weights1[31][271] = 16'b0000000000000011;
    assign weights1[31][272] = 16'b1111111111111110;
    assign weights1[31][273] = 16'b0000000000010101;
    assign weights1[31][274] = 16'b0000000000001011;
    assign weights1[31][275] = 16'b0000000000000101;
    assign weights1[31][276] = 16'b1111111111110110;
    assign weights1[31][277] = 16'b0000000000000001;
    assign weights1[31][278] = 16'b1111111111101000;
    assign weights1[31][279] = 16'b1111111111110000;
    assign weights1[31][280] = 16'b0000000000000010;
    assign weights1[31][281] = 16'b1111111111110011;
    assign weights1[31][282] = 16'b1111111111111001;
    assign weights1[31][283] = 16'b1111111111110110;
    assign weights1[31][284] = 16'b1111111111101011;
    assign weights1[31][285] = 16'b1111111111111110;
    assign weights1[31][286] = 16'b1111111111110110;
    assign weights1[31][287] = 16'b1111111111111001;
    assign weights1[31][288] = 16'b1111111111111111;
    assign weights1[31][289] = 16'b1111111111111100;
    assign weights1[31][290] = 16'b1111111111110011;
    assign weights1[31][291] = 16'b1111111111111010;
    assign weights1[31][292] = 16'b0000000000001001;
    assign weights1[31][293] = 16'b0000000000010011;
    assign weights1[31][294] = 16'b1111111111110010;
    assign weights1[31][295] = 16'b0000000000000100;
    assign weights1[31][296] = 16'b1111111111111101;
    assign weights1[31][297] = 16'b0000000000000101;
    assign weights1[31][298] = 16'b0000000000000110;
    assign weights1[31][299] = 16'b0000000000000010;
    assign weights1[31][300] = 16'b1111111111110010;
    assign weights1[31][301] = 16'b0000000000000000;
    assign weights1[31][302] = 16'b1111111111110111;
    assign weights1[31][303] = 16'b0000000000000111;
    assign weights1[31][304] = 16'b1111111111111101;
    assign weights1[31][305] = 16'b1111111111111110;
    assign weights1[31][306] = 16'b1111111111101011;
    assign weights1[31][307] = 16'b1111111111110100;
    assign weights1[31][308] = 16'b0000000000001001;
    assign weights1[31][309] = 16'b0000000000000110;
    assign weights1[31][310] = 16'b0000000000000100;
    assign weights1[31][311] = 16'b0000000000000011;
    assign weights1[31][312] = 16'b0000000000001100;
    assign weights1[31][313] = 16'b0000000000001100;
    assign weights1[31][314] = 16'b0000000000000010;
    assign weights1[31][315] = 16'b0000000000000010;
    assign weights1[31][316] = 16'b1111111111101011;
    assign weights1[31][317] = 16'b0000000000001111;
    assign weights1[31][318] = 16'b0000000000010111;
    assign weights1[31][319] = 16'b1111111111101101;
    assign weights1[31][320] = 16'b1111111111111010;
    assign weights1[31][321] = 16'b0000000000000001;
    assign weights1[31][322] = 16'b1111111111111001;
    assign weights1[31][323] = 16'b1111111111110111;
    assign weights1[31][324] = 16'b1111111111110110;
    assign weights1[31][325] = 16'b1111111111111111;
    assign weights1[31][326] = 16'b1111111111111100;
    assign weights1[31][327] = 16'b1111111111111011;
    assign weights1[31][328] = 16'b1111111111110110;
    assign weights1[31][329] = 16'b0000000000001101;
    assign weights1[31][330] = 16'b1111111111111111;
    assign weights1[31][331] = 16'b1111111111111001;
    assign weights1[31][332] = 16'b0000000000000010;
    assign weights1[31][333] = 16'b1111111111111110;
    assign weights1[31][334] = 16'b0000000000000011;
    assign weights1[31][335] = 16'b0000000000000010;
    assign weights1[31][336] = 16'b0000000000001001;
    assign weights1[31][337] = 16'b0000000000001010;
    assign weights1[31][338] = 16'b0000000000010111;
    assign weights1[31][339] = 16'b0000000000001010;
    assign weights1[31][340] = 16'b0000000000000111;
    assign weights1[31][341] = 16'b0000000000010001;
    assign weights1[31][342] = 16'b0000000000010011;
    assign weights1[31][343] = 16'b0000000000010000;
    assign weights1[31][344] = 16'b0000000000010100;
    assign weights1[31][345] = 16'b0000000000000110;
    assign weights1[31][346] = 16'b1111111111111000;
    assign weights1[31][347] = 16'b0000000000001011;
    assign weights1[31][348] = 16'b0000000000001010;
    assign weights1[31][349] = 16'b1111111111111100;
    assign weights1[31][350] = 16'b1111111111110100;
    assign weights1[31][351] = 16'b0000000000001101;
    assign weights1[31][352] = 16'b0000000000001110;
    assign weights1[31][353] = 16'b1111111111111110;
    assign weights1[31][354] = 16'b1111111111110101;
    assign weights1[31][355] = 16'b0000000000010001;
    assign weights1[31][356] = 16'b0000000000000011;
    assign weights1[31][357] = 16'b0000000000001001;
    assign weights1[31][358] = 16'b0000000000010100;
    assign weights1[31][359] = 16'b1111111111111101;
    assign weights1[31][360] = 16'b0000000000001100;
    assign weights1[31][361] = 16'b0000000000000011;
    assign weights1[31][362] = 16'b1111111111111000;
    assign weights1[31][363] = 16'b0000000000000101;
    assign weights1[31][364] = 16'b0000000000000011;
    assign weights1[31][365] = 16'b0000000000000101;
    assign weights1[31][366] = 16'b0000000000011010;
    assign weights1[31][367] = 16'b0000000000001001;
    assign weights1[31][368] = 16'b0000000000000101;
    assign weights1[31][369] = 16'b0000000000100110;
    assign weights1[31][370] = 16'b1111111111111000;
    assign weights1[31][371] = 16'b0000000000010001;
    assign weights1[31][372] = 16'b0000000000001100;
    assign weights1[31][373] = 16'b0000000000001110;
    assign weights1[31][374] = 16'b0000000000001011;
    assign weights1[31][375] = 16'b1111111111110010;
    assign weights1[31][376] = 16'b0000000000000001;
    assign weights1[31][377] = 16'b1111111111110010;
    assign weights1[31][378] = 16'b1111111111111011;
    assign weights1[31][379] = 16'b0000000000000101;
    assign weights1[31][380] = 16'b1111111111111100;
    assign weights1[31][381] = 16'b0000000000010011;
    assign weights1[31][382] = 16'b0000000000010001;
    assign weights1[31][383] = 16'b1111111111110011;
    assign weights1[31][384] = 16'b0000000000000000;
    assign weights1[31][385] = 16'b0000000000000101;
    assign weights1[31][386] = 16'b1111111111111100;
    assign weights1[31][387] = 16'b1111111111110111;
    assign weights1[31][388] = 16'b0000000000000000;
    assign weights1[31][389] = 16'b0000000000000011;
    assign weights1[31][390] = 16'b1111111111111011;
    assign weights1[31][391] = 16'b0000000000000011;
    assign weights1[31][392] = 16'b1111111111111101;
    assign weights1[31][393] = 16'b0000000000010010;
    assign weights1[31][394] = 16'b0000000000001101;
    assign weights1[31][395] = 16'b0000000000001001;
    assign weights1[31][396] = 16'b0000000000001001;
    assign weights1[31][397] = 16'b0000000000000010;
    assign weights1[31][398] = 16'b0000000000001110;
    assign weights1[31][399] = 16'b0000000000000101;
    assign weights1[31][400] = 16'b0000000000000100;
    assign weights1[31][401] = 16'b1111111111111101;
    assign weights1[31][402] = 16'b0000000000000010;
    assign weights1[31][403] = 16'b0000000000001011;
    assign weights1[31][404] = 16'b0000000000000100;
    assign weights1[31][405] = 16'b1111111111111111;
    assign weights1[31][406] = 16'b1111111111111110;
    assign weights1[31][407] = 16'b1111111111110110;
    assign weights1[31][408] = 16'b0000000000000101;
    assign weights1[31][409] = 16'b0000000000001101;
    assign weights1[31][410] = 16'b0000000000000001;
    assign weights1[31][411] = 16'b0000000000000101;
    assign weights1[31][412] = 16'b1111111111111000;
    assign weights1[31][413] = 16'b1111111111111010;
    assign weights1[31][414] = 16'b1111111111110101;
    assign weights1[31][415] = 16'b0000000000000110;
    assign weights1[31][416] = 16'b0000000000001100;
    assign weights1[31][417] = 16'b0000000000000000;
    assign weights1[31][418] = 16'b1111111111110000;
    assign weights1[31][419] = 16'b0000000000000101;
    assign weights1[31][420] = 16'b0000000000001101;
    assign weights1[31][421] = 16'b0000000000001011;
    assign weights1[31][422] = 16'b0000000000001001;
    assign weights1[31][423] = 16'b0000000000001011;
    assign weights1[31][424] = 16'b1111111111111010;
    assign weights1[31][425] = 16'b1111111111101100;
    assign weights1[31][426] = 16'b0000000000000000;
    assign weights1[31][427] = 16'b1111111111101101;
    assign weights1[31][428] = 16'b0000000000000111;
    assign weights1[31][429] = 16'b1111111111101101;
    assign weights1[31][430] = 16'b1111111111111101;
    assign weights1[31][431] = 16'b0000000000000001;
    assign weights1[31][432] = 16'b1111111111101101;
    assign weights1[31][433] = 16'b1111111111110010;
    assign weights1[31][434] = 16'b1111111111100101;
    assign weights1[31][435] = 16'b1111111111101101;
    assign weights1[31][436] = 16'b0000000000001011;
    assign weights1[31][437] = 16'b1111111111111100;
    assign weights1[31][438] = 16'b0000000000001100;
    assign weights1[31][439] = 16'b0000000000001000;
    assign weights1[31][440] = 16'b1111111111111101;
    assign weights1[31][441] = 16'b0000000000001100;
    assign weights1[31][442] = 16'b0000000000000110;
    assign weights1[31][443] = 16'b0000000000001000;
    assign weights1[31][444] = 16'b0000000000001011;
    assign weights1[31][445] = 16'b1111111111111001;
    assign weights1[31][446] = 16'b0000000000000111;
    assign weights1[31][447] = 16'b1111111111111110;
    assign weights1[31][448] = 16'b0000000000001111;
    assign weights1[31][449] = 16'b0000000000001011;
    assign weights1[31][450] = 16'b0000000000001110;
    assign weights1[31][451] = 16'b0000000000000111;
    assign weights1[31][452] = 16'b0000000000001101;
    assign weights1[31][453] = 16'b1111111111110101;
    assign weights1[31][454] = 16'b1111111111110111;
    assign weights1[31][455] = 16'b1111111111101110;
    assign weights1[31][456] = 16'b0000000000000110;
    assign weights1[31][457] = 16'b0000000000000010;
    assign weights1[31][458] = 16'b0000000000000001;
    assign weights1[31][459] = 16'b0000000000010010;
    assign weights1[31][460] = 16'b0000000000000010;
    assign weights1[31][461] = 16'b1111111111101101;
    assign weights1[31][462] = 16'b1111111111011110;
    assign weights1[31][463] = 16'b1111111111100111;
    assign weights1[31][464] = 16'b0000000000000001;
    assign weights1[31][465] = 16'b0000000000001110;
    assign weights1[31][466] = 16'b0000000000001101;
    assign weights1[31][467] = 16'b0000000000001011;
    assign weights1[31][468] = 16'b1111111111111100;
    assign weights1[31][469] = 16'b0000000000000011;
    assign weights1[31][470] = 16'b1111111111110111;
    assign weights1[31][471] = 16'b0000000000001001;
    assign weights1[31][472] = 16'b0000000000010000;
    assign weights1[31][473] = 16'b0000000000010101;
    assign weights1[31][474] = 16'b0000000000000110;
    assign weights1[31][475] = 16'b0000000000000011;
    assign weights1[31][476] = 16'b0000000000000010;
    assign weights1[31][477] = 16'b1111111111111001;
    assign weights1[31][478] = 16'b0000000000000110;
    assign weights1[31][479] = 16'b1111111111100111;
    assign weights1[31][480] = 16'b0000000000000100;
    assign weights1[31][481] = 16'b1111111111101101;
    assign weights1[31][482] = 16'b1111111111100011;
    assign weights1[31][483] = 16'b1111111111110000;
    assign weights1[31][484] = 16'b1111111111101100;
    assign weights1[31][485] = 16'b0000000000000010;
    assign weights1[31][486] = 16'b0000000000100001;
    assign weights1[31][487] = 16'b0000000000001100;
    assign weights1[31][488] = 16'b1111111111110000;
    assign weights1[31][489] = 16'b1111111111101010;
    assign weights1[31][490] = 16'b1111111111101000;
    assign weights1[31][491] = 16'b1111111111101100;
    assign weights1[31][492] = 16'b0000000000010000;
    assign weights1[31][493] = 16'b0000000000011101;
    assign weights1[31][494] = 16'b0000000000000101;
    assign weights1[31][495] = 16'b0000000000001000;
    assign weights1[31][496] = 16'b1111111111110101;
    assign weights1[31][497] = 16'b0000000000000001;
    assign weights1[31][498] = 16'b1111111111111110;
    assign weights1[31][499] = 16'b0000000000000000;
    assign weights1[31][500] = 16'b0000000000011011;
    assign weights1[31][501] = 16'b0000000000000111;
    assign weights1[31][502] = 16'b0000000000001010;
    assign weights1[31][503] = 16'b0000000000000011;
    assign weights1[31][504] = 16'b1111111111111010;
    assign weights1[31][505] = 16'b1111111111101110;
    assign weights1[31][506] = 16'b1111111111110100;
    assign weights1[31][507] = 16'b1111111111101011;
    assign weights1[31][508] = 16'b1111111111110001;
    assign weights1[31][509] = 16'b1111111111100100;
    assign weights1[31][510] = 16'b1111111111010011;
    assign weights1[31][511] = 16'b1111111111101100;
    assign weights1[31][512] = 16'b0000000000100000;
    assign weights1[31][513] = 16'b0000000000100100;
    assign weights1[31][514] = 16'b0000000000101000;
    assign weights1[31][515] = 16'b0000000000010110;
    assign weights1[31][516] = 16'b1111111111110110;
    assign weights1[31][517] = 16'b1111111111100011;
    assign weights1[31][518] = 16'b1111111111000000;
    assign weights1[31][519] = 16'b1111111111011011;
    assign weights1[31][520] = 16'b0000000000101000;
    assign weights1[31][521] = 16'b0000000000101010;
    assign weights1[31][522] = 16'b0000000000010101;
    assign weights1[31][523] = 16'b1111111111111101;
    assign weights1[31][524] = 16'b1111111111111011;
    assign weights1[31][525] = 16'b1111111111100111;
    assign weights1[31][526] = 16'b0000000000000100;
    assign weights1[31][527] = 16'b0000000000010100;
    assign weights1[31][528] = 16'b0000000000010110;
    assign weights1[31][529] = 16'b0000000000001100;
    assign weights1[31][530] = 16'b0000000000001010;
    assign weights1[31][531] = 16'b0000000000001000;
    assign weights1[31][532] = 16'b1111111111110010;
    assign weights1[31][533] = 16'b1111111111101001;
    assign weights1[31][534] = 16'b1111111111100100;
    assign weights1[31][535] = 16'b1111111111010000;
    assign weights1[31][536] = 16'b1111111111000101;
    assign weights1[31][537] = 16'b1111111111100100;
    assign weights1[31][538] = 16'b1111111111110011;
    assign weights1[31][539] = 16'b1111111111111100;
    assign weights1[31][540] = 16'b0000000000110100;
    assign weights1[31][541] = 16'b0000000000011011;
    assign weights1[31][542] = 16'b0000000000010001;
    assign weights1[31][543] = 16'b0000000000000000;
    assign weights1[31][544] = 16'b1111111111101101;
    assign weights1[31][545] = 16'b1111111111010001;
    assign weights1[31][546] = 16'b1111111110100010;
    assign weights1[31][547] = 16'b1111111111101100;
    assign weights1[31][548] = 16'b0000000000101101;
    assign weights1[31][549] = 16'b0000000000010111;
    assign weights1[31][550] = 16'b0000000000010011;
    assign weights1[31][551] = 16'b0000000000001000;
    assign weights1[31][552] = 16'b1111111111100000;
    assign weights1[31][553] = 16'b1111111111010110;
    assign weights1[31][554] = 16'b1111111111111000;
    assign weights1[31][555] = 16'b1111111111111010;
    assign weights1[31][556] = 16'b0000000000001101;
    assign weights1[31][557] = 16'b0000000000010111;
    assign weights1[31][558] = 16'b0000000000001101;
    assign weights1[31][559] = 16'b0000000000001111;
    assign weights1[31][560] = 16'b1111111111101101;
    assign weights1[31][561] = 16'b1111111111100101;
    assign weights1[31][562] = 16'b1111111111011111;
    assign weights1[31][563] = 16'b1111111111001000;
    assign weights1[31][564] = 16'b1111111111001000;
    assign weights1[31][565] = 16'b1111111111011101;
    assign weights1[31][566] = 16'b1111111111110111;
    assign weights1[31][567] = 16'b0000000000101000;
    assign weights1[31][568] = 16'b0000000000110101;
    assign weights1[31][569] = 16'b0000000000010001;
    assign weights1[31][570] = 16'b0000000000010011;
    assign weights1[31][571] = 16'b1111111111100001;
    assign weights1[31][572] = 16'b1111111111011010;
    assign weights1[31][573] = 16'b1111111110011011;
    assign weights1[31][574] = 16'b1111111110110111;
    assign weights1[31][575] = 16'b0000000000001010;
    assign weights1[31][576] = 16'b0000000000111010;
    assign weights1[31][577] = 16'b0000000000100000;
    assign weights1[31][578] = 16'b0000000000000101;
    assign weights1[31][579] = 16'b0000000000010011;
    assign weights1[31][580] = 16'b1111111111101101;
    assign weights1[31][581] = 16'b1111111111001100;
    assign weights1[31][582] = 16'b1111111111001000;
    assign weights1[31][583] = 16'b1111111111101001;
    assign weights1[31][584] = 16'b0000000000000010;
    assign weights1[31][585] = 16'b0000000000010000;
    assign weights1[31][586] = 16'b0000000000010001;
    assign weights1[31][587] = 16'b0000000000000110;
    assign weights1[31][588] = 16'b1111111111101001;
    assign weights1[31][589] = 16'b1111111111011100;
    assign weights1[31][590] = 16'b1111111111001100;
    assign weights1[31][591] = 16'b1111111111011011;
    assign weights1[31][592] = 16'b1111111111101000;
    assign weights1[31][593] = 16'b0000000000000111;
    assign weights1[31][594] = 16'b0000000000001110;
    assign weights1[31][595] = 16'b0000000000101101;
    assign weights1[31][596] = 16'b0000000001010101;
    assign weights1[31][597] = 16'b0000000000010111;
    assign weights1[31][598] = 16'b0000000000011000;
    assign weights1[31][599] = 16'b1111111111001101;
    assign weights1[31][600] = 16'b1111111110110100;
    assign weights1[31][601] = 16'b1111111101111100;
    assign weights1[31][602] = 16'b1111111111000101;
    assign weights1[31][603] = 16'b0000000000100111;
    assign weights1[31][604] = 16'b0000000000111110;
    assign weights1[31][605] = 16'b0000000000100001;
    assign weights1[31][606] = 16'b0000000000001001;
    assign weights1[31][607] = 16'b1111111111111110;
    assign weights1[31][608] = 16'b1111111111111001;
    assign weights1[31][609] = 16'b1111111111010001;
    assign weights1[31][610] = 16'b1111111110111001;
    assign weights1[31][611] = 16'b1111111111100111;
    assign weights1[31][612] = 16'b1111111111110100;
    assign weights1[31][613] = 16'b0000000000000110;
    assign weights1[31][614] = 16'b0000000000010000;
    assign weights1[31][615] = 16'b0000000000001000;
    assign weights1[31][616] = 16'b1111111111101100;
    assign weights1[31][617] = 16'b1111111111100011;
    assign weights1[31][618] = 16'b1111111111110010;
    assign weights1[31][619] = 16'b1111111111110111;
    assign weights1[31][620] = 16'b1111111111111111;
    assign weights1[31][621] = 16'b0000000000101000;
    assign weights1[31][622] = 16'b0000000001000000;
    assign weights1[31][623] = 16'b0000000001001001;
    assign weights1[31][624] = 16'b0000000000100111;
    assign weights1[31][625] = 16'b0000000000000000;
    assign weights1[31][626] = 16'b1111111111000000;
    assign weights1[31][627] = 16'b1111111110011110;
    assign weights1[31][628] = 16'b1111111110001101;
    assign weights1[31][629] = 16'b1111111101110101;
    assign weights1[31][630] = 16'b1111111111100011;
    assign weights1[31][631] = 16'b0000000000110000;
    assign weights1[31][632] = 16'b0000000000101101;
    assign weights1[31][633] = 16'b0000000000101001;
    assign weights1[31][634] = 16'b0000000000101111;
    assign weights1[31][635] = 16'b0000000000010000;
    assign weights1[31][636] = 16'b0000000000000010;
    assign weights1[31][637] = 16'b1111111111000000;
    assign weights1[31][638] = 16'b1111111110011011;
    assign weights1[31][639] = 16'b1111111110111101;
    assign weights1[31][640] = 16'b1111111111011111;
    assign weights1[31][641] = 16'b1111111111111110;
    assign weights1[31][642] = 16'b0000000000000100;
    assign weights1[31][643] = 16'b0000000000000011;
    assign weights1[31][644] = 16'b1111111111101101;
    assign weights1[31][645] = 16'b1111111111110110;
    assign weights1[31][646] = 16'b0000000000010110;
    assign weights1[31][647] = 16'b0000000000011001;
    assign weights1[31][648] = 16'b0000000000101001;
    assign weights1[31][649] = 16'b0000000000111001;
    assign weights1[31][650] = 16'b0000000000101011;
    assign weights1[31][651] = 16'b0000000000100110;
    assign weights1[31][652] = 16'b1111111111110110;
    assign weights1[31][653] = 16'b1111111111001001;
    assign weights1[31][654] = 16'b1111111110011111;
    assign weights1[31][655] = 16'b1111111110001100;
    assign weights1[31][656] = 16'b1111111110001010;
    assign weights1[31][657] = 16'b1111111110001000;
    assign weights1[31][658] = 16'b1111111111010101;
    assign weights1[31][659] = 16'b0000000000111110;
    assign weights1[31][660] = 16'b0000000000111101;
    assign weights1[31][661] = 16'b0000000000110111;
    assign weights1[31][662] = 16'b0000000000101101;
    assign weights1[31][663] = 16'b0000000000011101;
    assign weights1[31][664] = 16'b1111111111110010;
    assign weights1[31][665] = 16'b1111111110110011;
    assign weights1[31][666] = 16'b1111111110101101;
    assign weights1[31][667] = 16'b1111111110111011;
    assign weights1[31][668] = 16'b1111111111001110;
    assign weights1[31][669] = 16'b1111111111100111;
    assign weights1[31][670] = 16'b1111111111110110;
    assign weights1[31][671] = 16'b1111111111111011;
    assign weights1[31][672] = 16'b0000000000001000;
    assign weights1[31][673] = 16'b0000000000001110;
    assign weights1[31][674] = 16'b0000000000011110;
    assign weights1[31][675] = 16'b0000000000100100;
    assign weights1[31][676] = 16'b0000000000101011;
    assign weights1[31][677] = 16'b0000000000110110;
    assign weights1[31][678] = 16'b0000000000110001;
    assign weights1[31][679] = 16'b0000000000000111;
    assign weights1[31][680] = 16'b1111111111000100;
    assign weights1[31][681] = 16'b1111111110001011;
    assign weights1[31][682] = 16'b1111111101111001;
    assign weights1[31][683] = 16'b1111111101100000;
    assign weights1[31][684] = 16'b1111111110011000;
    assign weights1[31][685] = 16'b1111111111010101;
    assign weights1[31][686] = 16'b0000000000001110;
    assign weights1[31][687] = 16'b0000000000111010;
    assign weights1[31][688] = 16'b0000000001000011;
    assign weights1[31][689] = 16'b0000000000101100;
    assign weights1[31][690] = 16'b0000000000100110;
    assign weights1[31][691] = 16'b0000000000100000;
    assign weights1[31][692] = 16'b1111111111111100;
    assign weights1[31][693] = 16'b1111111110111100;
    assign weights1[31][694] = 16'b1111111110111001;
    assign weights1[31][695] = 16'b1111111110111100;
    assign weights1[31][696] = 16'b1111111111001110;
    assign weights1[31][697] = 16'b1111111111100000;
    assign weights1[31][698] = 16'b1111111111110100;
    assign weights1[31][699] = 16'b1111111111110111;
    assign weights1[31][700] = 16'b0000000000001000;
    assign weights1[31][701] = 16'b0000000000001101;
    assign weights1[31][702] = 16'b0000000000100000;
    assign weights1[31][703] = 16'b0000000000100011;
    assign weights1[31][704] = 16'b0000000000101110;
    assign weights1[31][705] = 16'b0000000000100000;
    assign weights1[31][706] = 16'b1111111111111110;
    assign weights1[31][707] = 16'b1111111111011000;
    assign weights1[31][708] = 16'b1111111110100001;
    assign weights1[31][709] = 16'b1111111110001000;
    assign weights1[31][710] = 16'b1111111101111000;
    assign weights1[31][711] = 16'b1111111101111010;
    assign weights1[31][712] = 16'b1111111110100000;
    assign weights1[31][713] = 16'b1111111110110110;
    assign weights1[31][714] = 16'b1111111111111111;
    assign weights1[31][715] = 16'b0000000000101010;
    assign weights1[31][716] = 16'b0000000000001111;
    assign weights1[31][717] = 16'b0000000000101011;
    assign weights1[31][718] = 16'b0000000000101010;
    assign weights1[31][719] = 16'b0000000000100000;
    assign weights1[31][720] = 16'b1111111111111000;
    assign weights1[31][721] = 16'b1111111111011010;
    assign weights1[31][722] = 16'b1111111110111011;
    assign weights1[31][723] = 16'b1111111110111101;
    assign weights1[31][724] = 16'b1111111111010011;
    assign weights1[31][725] = 16'b1111111111101001;
    assign weights1[31][726] = 16'b1111111111110001;
    assign weights1[31][727] = 16'b1111111111111000;
    assign weights1[31][728] = 16'b0000000000000111;
    assign weights1[31][729] = 16'b0000000000000001;
    assign weights1[31][730] = 16'b0000000000000110;
    assign weights1[31][731] = 16'b0000000000001001;
    assign weights1[31][732] = 16'b1111111111111111;
    assign weights1[31][733] = 16'b1111111111111011;
    assign weights1[31][734] = 16'b1111111111010101;
    assign weights1[31][735] = 16'b1111111110100111;
    assign weights1[31][736] = 16'b1111111110001110;
    assign weights1[31][737] = 16'b1111111101111110;
    assign weights1[31][738] = 16'b1111111101111011;
    assign weights1[31][739] = 16'b1111111110111011;
    assign weights1[31][740] = 16'b1111111111111100;
    assign weights1[31][741] = 16'b1111111111111110;
    assign weights1[31][742] = 16'b0000000000100111;
    assign weights1[31][743] = 16'b0000000000000001;
    assign weights1[31][744] = 16'b0000000000010001;
    assign weights1[31][745] = 16'b0000000000100001;
    assign weights1[31][746] = 16'b0000000000100101;
    assign weights1[31][747] = 16'b0000000000100100;
    assign weights1[31][748] = 16'b0000000000001001;
    assign weights1[31][749] = 16'b1111111111001111;
    assign weights1[31][750] = 16'b1111111111000110;
    assign weights1[31][751] = 16'b1111111111010101;
    assign weights1[31][752] = 16'b1111111111100011;
    assign weights1[31][753] = 16'b1111111111101111;
    assign weights1[31][754] = 16'b1111111111110101;
    assign weights1[31][755] = 16'b1111111111111110;
    assign weights1[31][756] = 16'b0000000000000100;
    assign weights1[31][757] = 16'b0000000000000010;
    assign weights1[31][758] = 16'b0000000000000001;
    assign weights1[31][759] = 16'b0000000000000000;
    assign weights1[31][760] = 16'b1111111111110111;
    assign weights1[31][761] = 16'b1111111111010111;
    assign weights1[31][762] = 16'b1111111110111111;
    assign weights1[31][763] = 16'b1111111110010101;
    assign weights1[31][764] = 16'b1111111110000111;
    assign weights1[31][765] = 16'b1111111101111000;
    assign weights1[31][766] = 16'b1111111110010010;
    assign weights1[31][767] = 16'b1111111110110010;
    assign weights1[31][768] = 16'b1111111111101100;
    assign weights1[31][769] = 16'b1111111111110100;
    assign weights1[31][770] = 16'b0000000000000000;
    assign weights1[31][771] = 16'b0000000000011110;
    assign weights1[31][772] = 16'b0000000001000111;
    assign weights1[31][773] = 16'b0000000001010100;
    assign weights1[31][774] = 16'b0000000001000100;
    assign weights1[31][775] = 16'b0000000000110011;
    assign weights1[31][776] = 16'b0000000000010100;
    assign weights1[31][777] = 16'b1111111111101000;
    assign weights1[31][778] = 16'b1111111111011111;
    assign weights1[31][779] = 16'b1111111111100100;
    assign weights1[31][780] = 16'b1111111111110001;
    assign weights1[31][781] = 16'b1111111111111000;
    assign weights1[31][782] = 16'b1111111111111010;
    assign weights1[31][783] = 16'b0000000000000001;
    assign weights1[32][0] = 16'b0000000000000000;
    assign weights1[32][1] = 16'b1111111111111111;
    assign weights1[32][2] = 16'b1111111111111110;
    assign weights1[32][3] = 16'b1111111111111100;
    assign weights1[32][4] = 16'b1111111111111101;
    assign weights1[32][5] = 16'b1111111111111010;
    assign weights1[32][6] = 16'b1111111111111000;
    assign weights1[32][7] = 16'b1111111111111001;
    assign weights1[32][8] = 16'b1111111111110100;
    assign weights1[32][9] = 16'b1111111111110110;
    assign weights1[32][10] = 16'b1111111111111011;
    assign weights1[32][11] = 16'b1111111111111110;
    assign weights1[32][12] = 16'b0000000000001001;
    assign weights1[32][13] = 16'b0000000000001001;
    assign weights1[32][14] = 16'b1111111111111110;
    assign weights1[32][15] = 16'b1111111111111111;
    assign weights1[32][16] = 16'b1111111111111001;
    assign weights1[32][17] = 16'b1111111111110100;
    assign weights1[32][18] = 16'b1111111111100011;
    assign weights1[32][19] = 16'b1111111111010001;
    assign weights1[32][20] = 16'b1111111111011100;
    assign weights1[32][21] = 16'b1111111111011001;
    assign weights1[32][22] = 16'b1111111111011011;
    assign weights1[32][23] = 16'b1111111111011111;
    assign weights1[32][24] = 16'b1111111111101000;
    assign weights1[32][25] = 16'b1111111111110000;
    assign weights1[32][26] = 16'b1111111111110111;
    assign weights1[32][27] = 16'b1111111111111010;
    assign weights1[32][28] = 16'b1111111111111111;
    assign weights1[32][29] = 16'b1111111111111100;
    assign weights1[32][30] = 16'b1111111111110110;
    assign weights1[32][31] = 16'b1111111111111010;
    assign weights1[32][32] = 16'b1111111111111011;
    assign weights1[32][33] = 16'b1111111111111000;
    assign weights1[32][34] = 16'b1111111111110001;
    assign weights1[32][35] = 16'b1111111111110111;
    assign weights1[32][36] = 16'b1111111111111011;
    assign weights1[32][37] = 16'b1111111111110000;
    assign weights1[32][38] = 16'b1111111111111011;
    assign weights1[32][39] = 16'b0000000000000100;
    assign weights1[32][40] = 16'b0000000000001001;
    assign weights1[32][41] = 16'b0000000000000100;
    assign weights1[32][42] = 16'b0000000000000010;
    assign weights1[32][43] = 16'b1111111111111000;
    assign weights1[32][44] = 16'b0000000000000000;
    assign weights1[32][45] = 16'b0000000000001010;
    assign weights1[32][46] = 16'b1111111111111011;
    assign weights1[32][47] = 16'b1111111111101100;
    assign weights1[32][48] = 16'b1111111111010011;
    assign weights1[32][49] = 16'b1111111111010101;
    assign weights1[32][50] = 16'b1111111111001010;
    assign weights1[32][51] = 16'b1111111111010100;
    assign weights1[32][52] = 16'b1111111111011101;
    assign weights1[32][53] = 16'b1111111111100101;
    assign weights1[32][54] = 16'b1111111111110100;
    assign weights1[32][55] = 16'b1111111111110111;
    assign weights1[32][56] = 16'b1111111111111111;
    assign weights1[32][57] = 16'b1111111111111001;
    assign weights1[32][58] = 16'b1111111111111001;
    assign weights1[32][59] = 16'b1111111111110111;
    assign weights1[32][60] = 16'b1111111111110101;
    assign weights1[32][61] = 16'b1111111111110011;
    assign weights1[32][62] = 16'b1111111111101011;
    assign weights1[32][63] = 16'b1111111111111010;
    assign weights1[32][64] = 16'b0000000000000100;
    assign weights1[32][65] = 16'b0000000000000110;
    assign weights1[32][66] = 16'b1111111111111100;
    assign weights1[32][67] = 16'b1111111111101101;
    assign weights1[32][68] = 16'b1111111111111101;
    assign weights1[32][69] = 16'b0000000000000011;
    assign weights1[32][70] = 16'b0000000000010110;
    assign weights1[32][71] = 16'b0000000000001001;
    assign weights1[32][72] = 16'b0000000000000110;
    assign weights1[32][73] = 16'b0000000000001100;
    assign weights1[32][74] = 16'b0000000000001111;
    assign weights1[32][75] = 16'b0000000000001001;
    assign weights1[32][76] = 16'b1111111111110000;
    assign weights1[32][77] = 16'b1111111111100111;
    assign weights1[32][78] = 16'b1111111111001001;
    assign weights1[32][79] = 16'b1111111111001110;
    assign weights1[32][80] = 16'b1111111111010110;
    assign weights1[32][81] = 16'b1111111111011001;
    assign weights1[32][82] = 16'b1111111111101100;
    assign weights1[32][83] = 16'b1111111111101111;
    assign weights1[32][84] = 16'b1111111111111101;
    assign weights1[32][85] = 16'b1111111111111100;
    assign weights1[32][86] = 16'b1111111111111011;
    assign weights1[32][87] = 16'b1111111111110001;
    assign weights1[32][88] = 16'b1111111111110010;
    assign weights1[32][89] = 16'b1111111111110100;
    assign weights1[32][90] = 16'b1111111111110100;
    assign weights1[32][91] = 16'b1111111111111001;
    assign weights1[32][92] = 16'b1111111111111110;
    assign weights1[32][93] = 16'b1111111111111001;
    assign weights1[32][94] = 16'b1111111111101111;
    assign weights1[32][95] = 16'b1111111111110010;
    assign weights1[32][96] = 16'b0000000000001000;
    assign weights1[32][97] = 16'b0000000000001011;
    assign weights1[32][98] = 16'b0000000000011000;
    assign weights1[32][99] = 16'b1111111111111101;
    assign weights1[32][100] = 16'b0000000000011011;
    assign weights1[32][101] = 16'b0000000000100101;
    assign weights1[32][102] = 16'b0000000000001111;
    assign weights1[32][103] = 16'b0000000000010010;
    assign weights1[32][104] = 16'b0000000000010011;
    assign weights1[32][105] = 16'b1111111111110101;
    assign weights1[32][106] = 16'b1111111111011010;
    assign weights1[32][107] = 16'b1111111111001010;
    assign weights1[32][108] = 16'b1111111111001000;
    assign weights1[32][109] = 16'b1111111111001111;
    assign weights1[32][110] = 16'b1111111111011101;
    assign weights1[32][111] = 16'b1111111111100110;
    assign weights1[32][112] = 16'b1111111111111111;
    assign weights1[32][113] = 16'b1111111111111001;
    assign weights1[32][114] = 16'b1111111111110011;
    assign weights1[32][115] = 16'b1111111111101110;
    assign weights1[32][116] = 16'b1111111111101101;
    assign weights1[32][117] = 16'b1111111111110000;
    assign weights1[32][118] = 16'b1111111111111001;
    assign weights1[32][119] = 16'b1111111111101111;
    assign weights1[32][120] = 16'b1111111111111011;
    assign weights1[32][121] = 16'b1111111111111001;
    assign weights1[32][122] = 16'b1111111111110111;
    assign weights1[32][123] = 16'b0000000000000001;
    assign weights1[32][124] = 16'b0000000000001010;
    assign weights1[32][125] = 16'b1111111111110101;
    assign weights1[32][126] = 16'b0000000000010001;
    assign weights1[32][127] = 16'b0000000000011100;
    assign weights1[32][128] = 16'b0000000000100000;
    assign weights1[32][129] = 16'b0000000000110110;
    assign weights1[32][130] = 16'b0000000000101100;
    assign weights1[32][131] = 16'b0000000000010101;
    assign weights1[32][132] = 16'b0000000000101001;
    assign weights1[32][133] = 16'b0000000000001011;
    assign weights1[32][134] = 16'b1111111111110101;
    assign weights1[32][135] = 16'b1111111111011100;
    assign weights1[32][136] = 16'b1111111111001110;
    assign weights1[32][137] = 16'b1111111111000110;
    assign weights1[32][138] = 16'b1111111111010100;
    assign weights1[32][139] = 16'b1111111111101010;
    assign weights1[32][140] = 16'b0000000000000000;
    assign weights1[32][141] = 16'b1111111111110110;
    assign weights1[32][142] = 16'b1111111111101100;
    assign weights1[32][143] = 16'b1111111111101101;
    assign weights1[32][144] = 16'b1111111111100100;
    assign weights1[32][145] = 16'b1111111111100010;
    assign weights1[32][146] = 16'b1111111111101011;
    assign weights1[32][147] = 16'b1111111111110101;
    assign weights1[32][148] = 16'b1111111111011110;
    assign weights1[32][149] = 16'b1111111111101011;
    assign weights1[32][150] = 16'b1111111111110011;
    assign weights1[32][151] = 16'b1111111111101100;
    assign weights1[32][152] = 16'b0000000000000101;
    assign weights1[32][153] = 16'b0000000000000010;
    assign weights1[32][154] = 16'b0000000000000000;
    assign weights1[32][155] = 16'b0000000000011011;
    assign weights1[32][156] = 16'b0000000000010111;
    assign weights1[32][157] = 16'b0000000000101000;
    assign weights1[32][158] = 16'b0000000000011011;
    assign weights1[32][159] = 16'b0000000000101011;
    assign weights1[32][160] = 16'b0000000000110111;
    assign weights1[32][161] = 16'b0000000000010110;
    assign weights1[32][162] = 16'b0000000000000110;
    assign weights1[32][163] = 16'b1111111111101000;
    assign weights1[32][164] = 16'b1111111111011011;
    assign weights1[32][165] = 16'b1111111111010110;
    assign weights1[32][166] = 16'b1111111111011001;
    assign weights1[32][167] = 16'b1111111111011111;
    assign weights1[32][168] = 16'b1111111111111100;
    assign weights1[32][169] = 16'b1111111111110100;
    assign weights1[32][170] = 16'b1111111111101110;
    assign weights1[32][171] = 16'b1111111111110111;
    assign weights1[32][172] = 16'b1111111111101101;
    assign weights1[32][173] = 16'b1111111111101100;
    assign weights1[32][174] = 16'b1111111111111010;
    assign weights1[32][175] = 16'b1111111111101111;
    assign weights1[32][176] = 16'b1111111111101011;
    assign weights1[32][177] = 16'b1111111111101101;
    assign weights1[32][178] = 16'b1111111111100010;
    assign weights1[32][179] = 16'b1111111111110001;
    assign weights1[32][180] = 16'b1111111111110010;
    assign weights1[32][181] = 16'b1111111111111111;
    assign weights1[32][182] = 16'b1111111111101110;
    assign weights1[32][183] = 16'b0000000000000000;
    assign weights1[32][184] = 16'b0000000000001000;
    assign weights1[32][185] = 16'b0000000000100100;
    assign weights1[32][186] = 16'b0000000000101001;
    assign weights1[32][187] = 16'b0000000000101011;
    assign weights1[32][188] = 16'b0000000000110101;
    assign weights1[32][189] = 16'b0000000000101010;
    assign weights1[32][190] = 16'b0000000000011000;
    assign weights1[32][191] = 16'b0000000000000101;
    assign weights1[32][192] = 16'b1111111111011111;
    assign weights1[32][193] = 16'b1111111111010110;
    assign weights1[32][194] = 16'b1111111111010101;
    assign weights1[32][195] = 16'b1111111111011001;
    assign weights1[32][196] = 16'b1111111111111100;
    assign weights1[32][197] = 16'b1111111111110111;
    assign weights1[32][198] = 16'b1111111111110011;
    assign weights1[32][199] = 16'b1111111111110111;
    assign weights1[32][200] = 16'b1111111111110110;
    assign weights1[32][201] = 16'b1111111111101000;
    assign weights1[32][202] = 16'b1111111111110010;
    assign weights1[32][203] = 16'b1111111111111001;
    assign weights1[32][204] = 16'b1111111111110000;
    assign weights1[32][205] = 16'b1111111111110110;
    assign weights1[32][206] = 16'b1111111111110110;
    assign weights1[32][207] = 16'b1111111111111010;
    assign weights1[32][208] = 16'b1111111111110011;
    assign weights1[32][209] = 16'b1111111111101111;
    assign weights1[32][210] = 16'b1111111111101111;
    assign weights1[32][211] = 16'b1111111111110110;
    assign weights1[32][212] = 16'b0000000000001010;
    assign weights1[32][213] = 16'b0000000000101011;
    assign weights1[32][214] = 16'b0000000001000000;
    assign weights1[32][215] = 16'b0000000000110010;
    assign weights1[32][216] = 16'b0000000000110001;
    assign weights1[32][217] = 16'b0000000000101000;
    assign weights1[32][218] = 16'b0000000000011111;
    assign weights1[32][219] = 16'b0000000000010100;
    assign weights1[32][220] = 16'b1111111111110100;
    assign weights1[32][221] = 16'b1111111111100111;
    assign weights1[32][222] = 16'b1111111111011001;
    assign weights1[32][223] = 16'b1111111111100000;
    assign weights1[32][224] = 16'b1111111111111010;
    assign weights1[32][225] = 16'b1111111111111001;
    assign weights1[32][226] = 16'b1111111111110001;
    assign weights1[32][227] = 16'b1111111111110000;
    assign weights1[32][228] = 16'b1111111111111011;
    assign weights1[32][229] = 16'b1111111111101111;
    assign weights1[32][230] = 16'b1111111111011101;
    assign weights1[32][231] = 16'b0000000000000111;
    assign weights1[32][232] = 16'b1111111111111110;
    assign weights1[32][233] = 16'b1111111111100010;
    assign weights1[32][234] = 16'b1111111111110101;
    assign weights1[32][235] = 16'b1111111111101110;
    assign weights1[32][236] = 16'b1111111111110000;
    assign weights1[32][237] = 16'b1111111111100101;
    assign weights1[32][238] = 16'b1111111111011111;
    assign weights1[32][239] = 16'b1111111111110001;
    assign weights1[32][240] = 16'b1111111111110011;
    assign weights1[32][241] = 16'b0000000000011001;
    assign weights1[32][242] = 16'b0000000001000001;
    assign weights1[32][243] = 16'b0000000000110110;
    assign weights1[32][244] = 16'b0000000000100110;
    assign weights1[32][245] = 16'b0000000000111011;
    assign weights1[32][246] = 16'b0000000000100010;
    assign weights1[32][247] = 16'b0000000000011001;
    assign weights1[32][248] = 16'b1111111111110101;
    assign weights1[32][249] = 16'b1111111111011111;
    assign weights1[32][250] = 16'b1111111111100000;
    assign weights1[32][251] = 16'b1111111111011101;
    assign weights1[32][252] = 16'b0000000000000010;
    assign weights1[32][253] = 16'b1111111111111001;
    assign weights1[32][254] = 16'b1111111111110011;
    assign weights1[32][255] = 16'b1111111111110110;
    assign weights1[32][256] = 16'b0000000000000101;
    assign weights1[32][257] = 16'b1111111111111011;
    assign weights1[32][258] = 16'b0000000000001100;
    assign weights1[32][259] = 16'b1111111111111101;
    assign weights1[32][260] = 16'b1111111111111011;
    assign weights1[32][261] = 16'b1111111111111010;
    assign weights1[32][262] = 16'b0000000000000001;
    assign weights1[32][263] = 16'b0000000000000101;
    assign weights1[32][264] = 16'b1111111111110100;
    assign weights1[32][265] = 16'b1111111111101001;
    assign weights1[32][266] = 16'b1111111111100010;
    assign weights1[32][267] = 16'b1111111111010010;
    assign weights1[32][268] = 16'b1111111111010011;
    assign weights1[32][269] = 16'b1111111111111100;
    assign weights1[32][270] = 16'b0000000000111001;
    assign weights1[32][271] = 16'b0000000001000010;
    assign weights1[32][272] = 16'b0000000000101011;
    assign weights1[32][273] = 16'b0000000000101000;
    assign weights1[32][274] = 16'b0000000000011100;
    assign weights1[32][275] = 16'b0000000000010001;
    assign weights1[32][276] = 16'b0000000000000101;
    assign weights1[32][277] = 16'b1111111111101010;
    assign weights1[32][278] = 16'b1111111111100110;
    assign weights1[32][279] = 16'b1111111111100011;
    assign weights1[32][280] = 16'b0000000000000010;
    assign weights1[32][281] = 16'b0000000000000011;
    assign weights1[32][282] = 16'b1111111111111101;
    assign weights1[32][283] = 16'b0000000000001011;
    assign weights1[32][284] = 16'b0000000000000010;
    assign weights1[32][285] = 16'b0000000000001001;
    assign weights1[32][286] = 16'b1111111111111010;
    assign weights1[32][287] = 16'b1111111111111010;
    assign weights1[32][288] = 16'b1111111111110101;
    assign weights1[32][289] = 16'b0000000000000000;
    assign weights1[32][290] = 16'b1111111111100100;
    assign weights1[32][291] = 16'b1111111111101010;
    assign weights1[32][292] = 16'b1111111111101010;
    assign weights1[32][293] = 16'b1111111111100000;
    assign weights1[32][294] = 16'b1111111111010101;
    assign weights1[32][295] = 16'b1111111111011110;
    assign weights1[32][296] = 16'b1111111111000001;
    assign weights1[32][297] = 16'b1111111111111100;
    assign weights1[32][298] = 16'b0000000000101111;
    assign weights1[32][299] = 16'b0000000000111111;
    assign weights1[32][300] = 16'b0000000000111111;
    assign weights1[32][301] = 16'b0000000000101000;
    assign weights1[32][302] = 16'b0000000000101110;
    assign weights1[32][303] = 16'b0000000000100110;
    assign weights1[32][304] = 16'b1111111111111100;
    assign weights1[32][305] = 16'b1111111111110000;
    assign weights1[32][306] = 16'b1111111111100000;
    assign weights1[32][307] = 16'b1111111111100011;
    assign weights1[32][308] = 16'b0000000000000011;
    assign weights1[32][309] = 16'b0000000000001010;
    assign weights1[32][310] = 16'b0000000000001111;
    assign weights1[32][311] = 16'b0000000000001011;
    assign weights1[32][312] = 16'b1111111111111011;
    assign weights1[32][313] = 16'b1111111111111011;
    assign weights1[32][314] = 16'b1111111111110100;
    assign weights1[32][315] = 16'b1111111111110111;
    assign weights1[32][316] = 16'b1111111111101110;
    assign weights1[32][317] = 16'b1111111111111011;
    assign weights1[32][318] = 16'b1111111111101101;
    assign weights1[32][319] = 16'b1111111111111000;
    assign weights1[32][320] = 16'b1111111111101001;
    assign weights1[32][321] = 16'b1111111111110010;
    assign weights1[32][322] = 16'b1111111111101100;
    assign weights1[32][323] = 16'b1111111111011001;
    assign weights1[32][324] = 16'b1111111111001110;
    assign weights1[32][325] = 16'b1111111111101101;
    assign weights1[32][326] = 16'b0000000000010011;
    assign weights1[32][327] = 16'b0000000000101000;
    assign weights1[32][328] = 16'b0000000000110011;
    assign weights1[32][329] = 16'b0000000000100110;
    assign weights1[32][330] = 16'b0000000000101110;
    assign weights1[32][331] = 16'b0000000000100110;
    assign weights1[32][332] = 16'b0000000000000100;
    assign weights1[32][333] = 16'b1111111111101110;
    assign weights1[32][334] = 16'b1111111111100010;
    assign weights1[32][335] = 16'b1111111111111000;
    assign weights1[32][336] = 16'b0000000000000111;
    assign weights1[32][337] = 16'b0000000000001100;
    assign weights1[32][338] = 16'b0000000000001000;
    assign weights1[32][339] = 16'b1111111111111010;
    assign weights1[32][340] = 16'b1111111111110100;
    assign weights1[32][341] = 16'b0000000000000100;
    assign weights1[32][342] = 16'b1111111111110010;
    assign weights1[32][343] = 16'b1111111111100001;
    assign weights1[32][344] = 16'b0000000000000100;
    assign weights1[32][345] = 16'b1111111111101101;
    assign weights1[32][346] = 16'b1111111111101000;
    assign weights1[32][347] = 16'b1111111111111000;
    assign weights1[32][348] = 16'b1111111111110010;
    assign weights1[32][349] = 16'b1111111111110001;
    assign weights1[32][350] = 16'b1111111111101011;
    assign weights1[32][351] = 16'b1111111111010011;
    assign weights1[32][352] = 16'b1111111110111001;
    assign weights1[32][353] = 16'b1111111111001100;
    assign weights1[32][354] = 16'b0000000000000100;
    assign weights1[32][355] = 16'b0000000000011100;
    assign weights1[32][356] = 16'b0000000000100000;
    assign weights1[32][357] = 16'b0000000000010110;
    assign weights1[32][358] = 16'b0000000000011110;
    assign weights1[32][359] = 16'b0000000000001101;
    assign weights1[32][360] = 16'b0000000000000101;
    assign weights1[32][361] = 16'b1111111111111000;
    assign weights1[32][362] = 16'b1111111111100100;
    assign weights1[32][363] = 16'b1111111111101111;
    assign weights1[32][364] = 16'b0000000000000111;
    assign weights1[32][365] = 16'b0000000000010000;
    assign weights1[32][366] = 16'b0000000000000000;
    assign weights1[32][367] = 16'b1111111111101101;
    assign weights1[32][368] = 16'b1111111111111010;
    assign weights1[32][369] = 16'b1111111111111011;
    assign weights1[32][370] = 16'b1111111111110100;
    assign weights1[32][371] = 16'b1111111111101111;
    assign weights1[32][372] = 16'b0000000000000000;
    assign weights1[32][373] = 16'b1111111111101101;
    assign weights1[32][374] = 16'b1111111111110011;
    assign weights1[32][375] = 16'b1111111111111000;
    assign weights1[32][376] = 16'b1111111111111010;
    assign weights1[32][377] = 16'b1111111111110110;
    assign weights1[32][378] = 16'b1111111111011110;
    assign weights1[32][379] = 16'b1111111110111001;
    assign weights1[32][380] = 16'b1111111110111101;
    assign weights1[32][381] = 16'b1111111111011000;
    assign weights1[32][382] = 16'b0000000000000101;
    assign weights1[32][383] = 16'b0000000000011010;
    assign weights1[32][384] = 16'b0000000000000101;
    assign weights1[32][385] = 16'b0000000000010110;
    assign weights1[32][386] = 16'b0000000000001001;
    assign weights1[32][387] = 16'b0000000000011011;
    assign weights1[32][388] = 16'b1111111111111110;
    assign weights1[32][389] = 16'b1111111111110111;
    assign weights1[32][390] = 16'b1111111111100110;
    assign weights1[32][391] = 16'b1111111111101110;
    assign weights1[32][392] = 16'b0000000000001011;
    assign weights1[32][393] = 16'b0000000000001001;
    assign weights1[32][394] = 16'b1111111111111010;
    assign weights1[32][395] = 16'b1111111111111011;
    assign weights1[32][396] = 16'b1111111111100101;
    assign weights1[32][397] = 16'b0000000000000101;
    assign weights1[32][398] = 16'b1111111111101010;
    assign weights1[32][399] = 16'b1111111111111011;
    assign weights1[32][400] = 16'b1111111111110010;
    assign weights1[32][401] = 16'b1111111111111110;
    assign weights1[32][402] = 16'b0000000000000010;
    assign weights1[32][403] = 16'b0000000000000010;
    assign weights1[32][404] = 16'b1111111111110110;
    assign weights1[32][405] = 16'b1111111111111000;
    assign weights1[32][406] = 16'b1111111111011010;
    assign weights1[32][407] = 16'b1111111111010010;
    assign weights1[32][408] = 16'b1111111110111100;
    assign weights1[32][409] = 16'b1111111111101000;
    assign weights1[32][410] = 16'b0000000000001101;
    assign weights1[32][411] = 16'b0000000000000001;
    assign weights1[32][412] = 16'b0000000000010100;
    assign weights1[32][413] = 16'b0000000000001101;
    assign weights1[32][414] = 16'b0000000000010011;
    assign weights1[32][415] = 16'b0000000000011011;
    assign weights1[32][416] = 16'b1111111111111001;
    assign weights1[32][417] = 16'b1111111111110001;
    assign weights1[32][418] = 16'b1111111111101111;
    assign weights1[32][419] = 16'b1111111111111001;
    assign weights1[32][420] = 16'b0000000000001101;
    assign weights1[32][421] = 16'b0000000000000100;
    assign weights1[32][422] = 16'b0000000000000110;
    assign weights1[32][423] = 16'b0000000000000011;
    assign weights1[32][424] = 16'b1111111111111010;
    assign weights1[32][425] = 16'b0000000000010001;
    assign weights1[32][426] = 16'b1111111111110010;
    assign weights1[32][427] = 16'b0000000000001100;
    assign weights1[32][428] = 16'b0000000000000110;
    assign weights1[32][429] = 16'b0000000000001111;
    assign weights1[32][430] = 16'b1111111111110101;
    assign weights1[32][431] = 16'b1111111111101111;
    assign weights1[32][432] = 16'b1111111111101100;
    assign weights1[32][433] = 16'b1111111111110001;
    assign weights1[32][434] = 16'b1111111111011011;
    assign weights1[32][435] = 16'b1111111111010010;
    assign weights1[32][436] = 16'b1111111111010110;
    assign weights1[32][437] = 16'b1111111111110100;
    assign weights1[32][438] = 16'b0000000000010011;
    assign weights1[32][439] = 16'b0000000000010111;
    assign weights1[32][440] = 16'b0000000000001000;
    assign weights1[32][441] = 16'b0000000000001000;
    assign weights1[32][442] = 16'b0000000000010010;
    assign weights1[32][443] = 16'b0000000000000001;
    assign weights1[32][444] = 16'b1111111111110001;
    assign weights1[32][445] = 16'b1111111111110010;
    assign weights1[32][446] = 16'b1111111111101110;
    assign weights1[32][447] = 16'b0000000000000110;
    assign weights1[32][448] = 16'b0000000000001001;
    assign weights1[32][449] = 16'b0000000000001010;
    assign weights1[32][450] = 16'b0000000000010000;
    assign weights1[32][451] = 16'b1111111111111110;
    assign weights1[32][452] = 16'b0000000000001010;
    assign weights1[32][453] = 16'b0000000000000101;
    assign weights1[32][454] = 16'b1111111111111101;
    assign weights1[32][455] = 16'b0000000000000000;
    assign weights1[32][456] = 16'b0000000000001011;
    assign weights1[32][457] = 16'b1111111111111001;
    assign weights1[32][458] = 16'b1111111111101101;
    assign weights1[32][459] = 16'b1111111111110100;
    assign weights1[32][460] = 16'b1111111111100011;
    assign weights1[32][461] = 16'b1111111111011110;
    assign weights1[32][462] = 16'b1111111111010100;
    assign weights1[32][463] = 16'b1111111111011111;
    assign weights1[32][464] = 16'b1111111111110001;
    assign weights1[32][465] = 16'b0000000000000111;
    assign weights1[32][466] = 16'b0000000000001100;
    assign weights1[32][467] = 16'b0000000000001010;
    assign weights1[32][468] = 16'b0000000000010111;
    assign weights1[32][469] = 16'b0000000000010110;
    assign weights1[32][470] = 16'b0000000000000101;
    assign weights1[32][471] = 16'b1111111111111000;
    assign weights1[32][472] = 16'b0000000000000000;
    assign weights1[32][473] = 16'b1111111111111100;
    assign weights1[32][474] = 16'b1111111111110110;
    assign weights1[32][475] = 16'b0000000000000010;
    assign weights1[32][476] = 16'b0000000000001001;
    assign weights1[32][477] = 16'b0000000000001001;
    assign weights1[32][478] = 16'b0000000000011000;
    assign weights1[32][479] = 16'b0000000000000010;
    assign weights1[32][480] = 16'b0000000000011010;
    assign weights1[32][481] = 16'b0000000000000001;
    assign weights1[32][482] = 16'b1111111111111111;
    assign weights1[32][483] = 16'b1111111111111100;
    assign weights1[32][484] = 16'b1111111111111111;
    assign weights1[32][485] = 16'b1111111111111111;
    assign weights1[32][486] = 16'b1111111111111011;
    assign weights1[32][487] = 16'b1111111111110011;
    assign weights1[32][488] = 16'b1111111111100000;
    assign weights1[32][489] = 16'b1111111111110100;
    assign weights1[32][490] = 16'b1111111111101001;
    assign weights1[32][491] = 16'b1111111111110010;
    assign weights1[32][492] = 16'b1111111111110110;
    assign weights1[32][493] = 16'b0000000000000000;
    assign weights1[32][494] = 16'b0000000000001111;
    assign weights1[32][495] = 16'b0000000000010110;
    assign weights1[32][496] = 16'b0000000000001100;
    assign weights1[32][497] = 16'b1111111111110010;
    assign weights1[32][498] = 16'b1111111111110111;
    assign weights1[32][499] = 16'b1111111111100100;
    assign weights1[32][500] = 16'b1111111111101111;
    assign weights1[32][501] = 16'b1111111111110111;
    assign weights1[32][502] = 16'b1111111111111100;
    assign weights1[32][503] = 16'b0000000000000010;
    assign weights1[32][504] = 16'b0000000000000100;
    assign weights1[32][505] = 16'b0000000000000000;
    assign weights1[32][506] = 16'b0000000000001010;
    assign weights1[32][507] = 16'b0000000000000110;
    assign weights1[32][508] = 16'b0000000000001011;
    assign weights1[32][509] = 16'b0000000000010000;
    assign weights1[32][510] = 16'b0000000000010000;
    assign weights1[32][511] = 16'b1111111111111110;
    assign weights1[32][512] = 16'b0000000000000101;
    assign weights1[32][513] = 16'b0000000000000001;
    assign weights1[32][514] = 16'b0000000000010011;
    assign weights1[32][515] = 16'b1111111111101001;
    assign weights1[32][516] = 16'b1111111111100011;
    assign weights1[32][517] = 16'b1111111111101100;
    assign weights1[32][518] = 16'b1111111111110110;
    assign weights1[32][519] = 16'b1111111111110010;
    assign weights1[32][520] = 16'b1111111111110101;
    assign weights1[32][521] = 16'b1111111111111111;
    assign weights1[32][522] = 16'b1111111111111000;
    assign weights1[32][523] = 16'b0000000000001011;
    assign weights1[32][524] = 16'b1111111111101110;
    assign weights1[32][525] = 16'b1111111111101101;
    assign weights1[32][526] = 16'b1111111111101010;
    assign weights1[32][527] = 16'b1111111111100000;
    assign weights1[32][528] = 16'b1111111111101110;
    assign weights1[32][529] = 16'b1111111111110001;
    assign weights1[32][530] = 16'b1111111111111000;
    assign weights1[32][531] = 16'b1111111111111011;
    assign weights1[32][532] = 16'b0000000000000000;
    assign weights1[32][533] = 16'b1111111111111111;
    assign weights1[32][534] = 16'b1111111111111010;
    assign weights1[32][535] = 16'b0000000000000001;
    assign weights1[32][536] = 16'b1111111111110101;
    assign weights1[32][537] = 16'b0000000000000001;
    assign weights1[32][538] = 16'b0000000000000010;
    assign weights1[32][539] = 16'b1111111111111001;
    assign weights1[32][540] = 16'b0000000000001100;
    assign weights1[32][541] = 16'b0000000000010010;
    assign weights1[32][542] = 16'b0000000000000110;
    assign weights1[32][543] = 16'b0000000000000000;
    assign weights1[32][544] = 16'b1111111111111000;
    assign weights1[32][545] = 16'b1111111111111101;
    assign weights1[32][546] = 16'b0000000000001001;
    assign weights1[32][547] = 16'b0000000000000000;
    assign weights1[32][548] = 16'b1111111111111111;
    assign weights1[32][549] = 16'b0000000000000011;
    assign weights1[32][550] = 16'b1111111111111100;
    assign weights1[32][551] = 16'b0000000000000100;
    assign weights1[32][552] = 16'b1111111111110100;
    assign weights1[32][553] = 16'b1111111111110100;
    assign weights1[32][554] = 16'b1111111111111011;
    assign weights1[32][555] = 16'b1111111111111010;
    assign weights1[32][556] = 16'b1111111111110100;
    assign weights1[32][557] = 16'b1111111111111000;
    assign weights1[32][558] = 16'b1111111111111010;
    assign weights1[32][559] = 16'b0000000000000100;
    assign weights1[32][560] = 16'b1111111111111100;
    assign weights1[32][561] = 16'b1111111111111001;
    assign weights1[32][562] = 16'b1111111111110110;
    assign weights1[32][563] = 16'b0000000000000101;
    assign weights1[32][564] = 16'b0000000000000111;
    assign weights1[32][565] = 16'b0000000000001101;
    assign weights1[32][566] = 16'b0000000000000011;
    assign weights1[32][567] = 16'b1111111111110101;
    assign weights1[32][568] = 16'b1111111111111001;
    assign weights1[32][569] = 16'b1111111111111111;
    assign weights1[32][570] = 16'b0000000000011010;
    assign weights1[32][571] = 16'b0000000000000011;
    assign weights1[32][572] = 16'b0000000000001011;
    assign weights1[32][573] = 16'b0000000000001000;
    assign weights1[32][574] = 16'b0000000000001000;
    assign weights1[32][575] = 16'b0000000000000001;
    assign weights1[32][576] = 16'b1111111111110011;
    assign weights1[32][577] = 16'b0000000000001001;
    assign weights1[32][578] = 16'b0000000000000110;
    assign weights1[32][579] = 16'b1111111111111111;
    assign weights1[32][580] = 16'b1111111111110110;
    assign weights1[32][581] = 16'b0000000000000101;
    assign weights1[32][582] = 16'b1111111111111010;
    assign weights1[32][583] = 16'b0000000000001010;
    assign weights1[32][584] = 16'b1111111111110101;
    assign weights1[32][585] = 16'b0000000000000000;
    assign weights1[32][586] = 16'b0000000000000000;
    assign weights1[32][587] = 16'b0000000000001101;
    assign weights1[32][588] = 16'b1111111111111011;
    assign weights1[32][589] = 16'b0000000000000001;
    assign weights1[32][590] = 16'b1111111111110010;
    assign weights1[32][591] = 16'b1111111111111001;
    assign weights1[32][592] = 16'b0000000000001000;
    assign weights1[32][593] = 16'b0000000000010110;
    assign weights1[32][594] = 16'b0000000000000001;
    assign weights1[32][595] = 16'b1111111111111111;
    assign weights1[32][596] = 16'b1111111111110100;
    assign weights1[32][597] = 16'b1111111111111010;
    assign weights1[32][598] = 16'b1111111111111110;
    assign weights1[32][599] = 16'b0000000000010110;
    assign weights1[32][600] = 16'b0000000000001011;
    assign weights1[32][601] = 16'b0000000000000111;
    assign weights1[32][602] = 16'b0000000000000001;
    assign weights1[32][603] = 16'b1111111111111000;
    assign weights1[32][604] = 16'b0000000000000001;
    assign weights1[32][605] = 16'b1111111111111101;
    assign weights1[32][606] = 16'b1111111111110001;
    assign weights1[32][607] = 16'b1111111111111111;
    assign weights1[32][608] = 16'b1111111111110010;
    assign weights1[32][609] = 16'b1111111111111111;
    assign weights1[32][610] = 16'b1111111111111100;
    assign weights1[32][611] = 16'b0000000000010000;
    assign weights1[32][612] = 16'b0000000000001110;
    assign weights1[32][613] = 16'b0000000000000001;
    assign weights1[32][614] = 16'b0000000000000000;
    assign weights1[32][615] = 16'b0000000000001111;
    assign weights1[32][616] = 16'b1111111111111110;
    assign weights1[32][617] = 16'b1111111111111101;
    assign weights1[32][618] = 16'b1111111111111111;
    assign weights1[32][619] = 16'b1111111111111110;
    assign weights1[32][620] = 16'b1111111111111011;
    assign weights1[32][621] = 16'b1111111111111000;
    assign weights1[32][622] = 16'b1111111111110011;
    assign weights1[32][623] = 16'b0000000000001001;
    assign weights1[32][624] = 16'b1111111111111010;
    assign weights1[32][625] = 16'b0000000000001011;
    assign weights1[32][626] = 16'b0000000000010111;
    assign weights1[32][627] = 16'b0000000000010011;
    assign weights1[32][628] = 16'b0000000000010011;
    assign weights1[32][629] = 16'b0000000000000001;
    assign weights1[32][630] = 16'b1111111111111111;
    assign weights1[32][631] = 16'b1111111111110010;
    assign weights1[32][632] = 16'b0000000000001101;
    assign weights1[32][633] = 16'b1111111111111101;
    assign weights1[32][634] = 16'b1111111111111101;
    assign weights1[32][635] = 16'b1111111111111110;
    assign weights1[32][636] = 16'b1111111111111110;
    assign weights1[32][637] = 16'b0000000000000010;
    assign weights1[32][638] = 16'b1111111111111001;
    assign weights1[32][639] = 16'b0000000000011011;
    assign weights1[32][640] = 16'b0000000000000000;
    assign weights1[32][641] = 16'b1111111111111001;
    assign weights1[32][642] = 16'b0000000000001001;
    assign weights1[32][643] = 16'b0000000000001001;
    assign weights1[32][644] = 16'b1111111111111110;
    assign weights1[32][645] = 16'b0000000000000000;
    assign weights1[32][646] = 16'b1111111111111111;
    assign weights1[32][647] = 16'b1111111111111010;
    assign weights1[32][648] = 16'b1111111111111101;
    assign weights1[32][649] = 16'b1111111111110101;
    assign weights1[32][650] = 16'b0000000000001111;
    assign weights1[32][651] = 16'b0000000000001101;
    assign weights1[32][652] = 16'b0000000000000010;
    assign weights1[32][653] = 16'b1111111111111011;
    assign weights1[32][654] = 16'b0000000000011100;
    assign weights1[32][655] = 16'b0000000000010111;
    assign weights1[32][656] = 16'b0000000000001100;
    assign weights1[32][657] = 16'b0000000000000101;
    assign weights1[32][658] = 16'b0000000000001010;
    assign weights1[32][659] = 16'b1111111111111100;
    assign weights1[32][660] = 16'b0000000000010001;
    assign weights1[32][661] = 16'b0000000000000101;
    assign weights1[32][662] = 16'b1111111111110101;
    assign weights1[32][663] = 16'b1111111111111111;
    assign weights1[32][664] = 16'b1111111111111101;
    assign weights1[32][665] = 16'b0000000000001110;
    assign weights1[32][666] = 16'b0000000000000101;
    assign weights1[32][667] = 16'b0000000000001011;
    assign weights1[32][668] = 16'b0000000000000001;
    assign weights1[32][669] = 16'b1111111111111110;
    assign weights1[32][670] = 16'b1111111111111111;
    assign weights1[32][671] = 16'b0000000000000101;
    assign weights1[32][672] = 16'b0000000000000000;
    assign weights1[32][673] = 16'b1111111111111101;
    assign weights1[32][674] = 16'b1111111111111011;
    assign weights1[32][675] = 16'b1111111111111001;
    assign weights1[32][676] = 16'b0000000000000110;
    assign weights1[32][677] = 16'b0000000000011000;
    assign weights1[32][678] = 16'b0000000000010011;
    assign weights1[32][679] = 16'b0000000000000000;
    assign weights1[32][680] = 16'b1111111111111001;
    assign weights1[32][681] = 16'b0000000000010000;
    assign weights1[32][682] = 16'b0000000000011110;
    assign weights1[32][683] = 16'b0000000000001010;
    assign weights1[32][684] = 16'b0000000000000111;
    assign weights1[32][685] = 16'b1111111111110111;
    assign weights1[32][686] = 16'b1111111111101101;
    assign weights1[32][687] = 16'b1111111111101011;
    assign weights1[32][688] = 16'b0000000000001000;
    assign weights1[32][689] = 16'b1111111111111011;
    assign weights1[32][690] = 16'b1111111111111000;
    assign weights1[32][691] = 16'b0000000000000000;
    assign weights1[32][692] = 16'b0000000000000010;
    assign weights1[32][693] = 16'b0000000000001000;
    assign weights1[32][694] = 16'b1111111111111010;
    assign weights1[32][695] = 16'b1111111111111111;
    assign weights1[32][696] = 16'b0000000000000000;
    assign weights1[32][697] = 16'b0000000000000101;
    assign weights1[32][698] = 16'b1111111111111011;
    assign weights1[32][699] = 16'b1111111111111110;
    assign weights1[32][700] = 16'b1111111111111111;
    assign weights1[32][701] = 16'b1111111111111110;
    assign weights1[32][702] = 16'b1111111111111001;
    assign weights1[32][703] = 16'b1111111111111000;
    assign weights1[32][704] = 16'b1111111111111111;
    assign weights1[32][705] = 16'b0000000000000011;
    assign weights1[32][706] = 16'b0000000000000100;
    assign weights1[32][707] = 16'b0000000000001010;
    assign weights1[32][708] = 16'b0000000000010101;
    assign weights1[32][709] = 16'b0000000000011101;
    assign weights1[32][710] = 16'b0000000000011101;
    assign weights1[32][711] = 16'b0000000000000000;
    assign weights1[32][712] = 16'b1111111111111011;
    assign weights1[32][713] = 16'b1111111111111101;
    assign weights1[32][714] = 16'b1111111111110101;
    assign weights1[32][715] = 16'b1111111111110010;
    assign weights1[32][716] = 16'b1111111111110011;
    assign weights1[32][717] = 16'b1111111111111010;
    assign weights1[32][718] = 16'b1111111111111010;
    assign weights1[32][719] = 16'b1111111111110101;
    assign weights1[32][720] = 16'b1111111111110110;
    assign weights1[32][721] = 16'b0000000000001001;
    assign weights1[32][722] = 16'b1111111111111000;
    assign weights1[32][723] = 16'b1111111111111100;
    assign weights1[32][724] = 16'b1111111111111100;
    assign weights1[32][725] = 16'b1111111111111011;
    assign weights1[32][726] = 16'b1111111111111000;
    assign weights1[32][727] = 16'b1111111111111110;
    assign weights1[32][728] = 16'b1111111111111110;
    assign weights1[32][729] = 16'b0000000000000001;
    assign weights1[32][730] = 16'b1111111111111000;
    assign weights1[32][731] = 16'b1111111111111011;
    assign weights1[32][732] = 16'b1111111111111111;
    assign weights1[32][733] = 16'b1111111111110010;
    assign weights1[32][734] = 16'b1111111111110010;
    assign weights1[32][735] = 16'b1111111111111110;
    assign weights1[32][736] = 16'b0000000000001101;
    assign weights1[32][737] = 16'b0000000000001110;
    assign weights1[32][738] = 16'b0000000000000101;
    assign weights1[32][739] = 16'b1111111111110001;
    assign weights1[32][740] = 16'b1111111111101000;
    assign weights1[32][741] = 16'b1111111111111000;
    assign weights1[32][742] = 16'b1111111111111001;
    assign weights1[32][743] = 16'b0000000000000000;
    assign weights1[32][744] = 16'b1111111111111000;
    assign weights1[32][745] = 16'b0000000000000000;
    assign weights1[32][746] = 16'b1111111111110001;
    assign weights1[32][747] = 16'b1111111111110101;
    assign weights1[32][748] = 16'b0000000000001010;
    assign weights1[32][749] = 16'b0000000000000010;
    assign weights1[32][750] = 16'b1111111111111111;
    assign weights1[32][751] = 16'b1111111111111000;
    assign weights1[32][752] = 16'b1111111111110110;
    assign weights1[32][753] = 16'b1111111111110100;
    assign weights1[32][754] = 16'b1111111111111110;
    assign weights1[32][755] = 16'b1111111111111111;
    assign weights1[32][756] = 16'b1111111111111111;
    assign weights1[32][757] = 16'b1111111111111111;
    assign weights1[32][758] = 16'b1111111111111111;
    assign weights1[32][759] = 16'b0000000000000001;
    assign weights1[32][760] = 16'b1111111111111101;
    assign weights1[32][761] = 16'b0000000000000100;
    assign weights1[32][762] = 16'b0000000000000110;
    assign weights1[32][763] = 16'b0000000000000000;
    assign weights1[32][764] = 16'b1111111111110111;
    assign weights1[32][765] = 16'b1111111111100100;
    assign weights1[32][766] = 16'b1111111111101001;
    assign weights1[32][767] = 16'b1111111111110011;
    assign weights1[32][768] = 16'b1111111111110000;
    assign weights1[32][769] = 16'b1111111111101110;
    assign weights1[32][770] = 16'b1111111111101110;
    assign weights1[32][771] = 16'b1111111111110000;
    assign weights1[32][772] = 16'b1111111111101101;
    assign weights1[32][773] = 16'b1111111111110111;
    assign weights1[32][774] = 16'b1111111111110101;
    assign weights1[32][775] = 16'b1111111111110110;
    assign weights1[32][776] = 16'b1111111111111011;
    assign weights1[32][777] = 16'b1111111111110110;
    assign weights1[32][778] = 16'b1111111111111000;
    assign weights1[32][779] = 16'b1111111111111000;
    assign weights1[32][780] = 16'b1111111111111010;
    assign weights1[32][781] = 16'b1111111111111101;
    assign weights1[32][782] = 16'b1111111111111111;
    assign weights1[32][783] = 16'b0000000000000001;
    assign weights1[33][0] = 16'b0000000000000000;
    assign weights1[33][1] = 16'b0000000000000001;
    assign weights1[33][2] = 16'b0000000000000011;
    assign weights1[33][3] = 16'b0000000000001011;
    assign weights1[33][4] = 16'b0000000000001001;
    assign weights1[33][5] = 16'b0000000000001010;
    assign weights1[33][6] = 16'b0000000000001101;
    assign weights1[33][7] = 16'b0000000000010100;
    assign weights1[33][8] = 16'b0000000000000110;
    assign weights1[33][9] = 16'b0000000000001101;
    assign weights1[33][10] = 16'b0000000000001110;
    assign weights1[33][11] = 16'b0000000000011100;
    assign weights1[33][12] = 16'b0000000000001100;
    assign weights1[33][13] = 16'b0000000000011111;
    assign weights1[33][14] = 16'b0000000000010110;
    assign weights1[33][15] = 16'b0000000000001110;
    assign weights1[33][16] = 16'b0000000000001111;
    assign weights1[33][17] = 16'b0000000000001111;
    assign weights1[33][18] = 16'b0000000000010010;
    assign weights1[33][19] = 16'b0000000000000100;
    assign weights1[33][20] = 16'b0000000000000000;
    assign weights1[33][21] = 16'b0000000000011001;
    assign weights1[33][22] = 16'b1111111111111001;
    assign weights1[33][23] = 16'b1111111111111010;
    assign weights1[33][24] = 16'b1111111111111101;
    assign weights1[33][25] = 16'b1111111111101110;
    assign weights1[33][26] = 16'b1111111111111010;
    assign weights1[33][27] = 16'b1111111111111100;
    assign weights1[33][28] = 16'b0000000000000001;
    assign weights1[33][29] = 16'b0000000000000001;
    assign weights1[33][30] = 16'b0000000000000001;
    assign weights1[33][31] = 16'b0000000000000010;
    assign weights1[33][32] = 16'b0000000000001100;
    assign weights1[33][33] = 16'b0000000000001101;
    assign weights1[33][34] = 16'b0000000000000000;
    assign weights1[33][35] = 16'b0000000000010100;
    assign weights1[33][36] = 16'b1111111111111101;
    assign weights1[33][37] = 16'b0000000000001000;
    assign weights1[33][38] = 16'b0000000000001000;
    assign weights1[33][39] = 16'b0000000000000000;
    assign weights1[33][40] = 16'b0000000000000110;
    assign weights1[33][41] = 16'b0000000000001001;
    assign weights1[33][42] = 16'b1111111111111011;
    assign weights1[33][43] = 16'b1111111111110011;
    assign weights1[33][44] = 16'b1111111111111111;
    assign weights1[33][45] = 16'b0000000000000001;
    assign weights1[33][46] = 16'b0000000000000000;
    assign weights1[33][47] = 16'b1111111111111100;
    assign weights1[33][48] = 16'b0000000000000101;
    assign weights1[33][49] = 16'b0000000000000000;
    assign weights1[33][50] = 16'b0000000000000111;
    assign weights1[33][51] = 16'b0000000000000000;
    assign weights1[33][52] = 16'b0000000000000000;
    assign weights1[33][53] = 16'b1111111111111011;
    assign weights1[33][54] = 16'b1111111111110000;
    assign weights1[33][55] = 16'b1111111111111010;
    assign weights1[33][56] = 16'b0000000000000001;
    assign weights1[33][57] = 16'b0000000000000010;
    assign weights1[33][58] = 16'b1111111111111101;
    assign weights1[33][59] = 16'b1111111111111110;
    assign weights1[33][60] = 16'b0000000000001011;
    assign weights1[33][61] = 16'b0000000000001001;
    assign weights1[33][62] = 16'b0000000000001000;
    assign weights1[33][63] = 16'b0000000000000011;
    assign weights1[33][64] = 16'b1111111111110010;
    assign weights1[33][65] = 16'b1111111111111000;
    assign weights1[33][66] = 16'b0000000000000001;
    assign weights1[33][67] = 16'b1111111111110011;
    assign weights1[33][68] = 16'b1111111111111110;
    assign weights1[33][69] = 16'b1111111111110001;
    assign weights1[33][70] = 16'b0000000000001110;
    assign weights1[33][71] = 16'b1111111111110011;
    assign weights1[33][72] = 16'b0000000000000010;
    assign weights1[33][73] = 16'b0000000000001000;
    assign weights1[33][74] = 16'b1111111111110010;
    assign weights1[33][75] = 16'b1111111111111000;
    assign weights1[33][76] = 16'b1111111111101111;
    assign weights1[33][77] = 16'b1111111111111010;
    assign weights1[33][78] = 16'b0000000000001100;
    assign weights1[33][79] = 16'b1111111111110100;
    assign weights1[33][80] = 16'b1111111111111101;
    assign weights1[33][81] = 16'b1111111111111001;
    assign weights1[33][82] = 16'b1111111111111001;
    assign weights1[33][83] = 16'b1111111111110010;
    assign weights1[33][84] = 16'b1111111111111111;
    assign weights1[33][85] = 16'b0000000000000001;
    assign weights1[33][86] = 16'b0000000000000000;
    assign weights1[33][87] = 16'b0000000000000100;
    assign weights1[33][88] = 16'b0000000000010011;
    assign weights1[33][89] = 16'b0000000000000001;
    assign weights1[33][90] = 16'b0000000000000111;
    assign weights1[33][91] = 16'b1111111111111000;
    assign weights1[33][92] = 16'b1111111111110000;
    assign weights1[33][93] = 16'b0000000000000000;
    assign weights1[33][94] = 16'b0000000000000010;
    assign weights1[33][95] = 16'b0000000000000101;
    assign weights1[33][96] = 16'b0000000000000100;
    assign weights1[33][97] = 16'b0000000000001110;
    assign weights1[33][98] = 16'b1111111111111110;
    assign weights1[33][99] = 16'b0000000000001000;
    assign weights1[33][100] = 16'b0000000000000001;
    assign weights1[33][101] = 16'b1111111111111100;
    assign weights1[33][102] = 16'b1111111111111100;
    assign weights1[33][103] = 16'b0000000000001110;
    assign weights1[33][104] = 16'b1111111111111101;
    assign weights1[33][105] = 16'b1111111111111100;
    assign weights1[33][106] = 16'b1111111111111001;
    assign weights1[33][107] = 16'b0000000000001100;
    assign weights1[33][108] = 16'b1111111111111100;
    assign weights1[33][109] = 16'b1111111111111001;
    assign weights1[33][110] = 16'b1111111111101100;
    assign weights1[33][111] = 16'b1111111111110010;
    assign weights1[33][112] = 16'b1111111111111101;
    assign weights1[33][113] = 16'b1111111111111100;
    assign weights1[33][114] = 16'b1111111111111100;
    assign weights1[33][115] = 16'b1111111111110100;
    assign weights1[33][116] = 16'b0000000000001100;
    assign weights1[33][117] = 16'b0000000000000111;
    assign weights1[33][118] = 16'b1111111111111000;
    assign weights1[33][119] = 16'b1111111111110001;
    assign weights1[33][120] = 16'b1111111111110011;
    assign weights1[33][121] = 16'b1111111111101101;
    assign weights1[33][122] = 16'b1111111111111110;
    assign weights1[33][123] = 16'b1111111111101100;
    assign weights1[33][124] = 16'b1111111111101011;
    assign weights1[33][125] = 16'b1111111111111110;
    assign weights1[33][126] = 16'b1111111111110001;
    assign weights1[33][127] = 16'b1111111111111101;
    assign weights1[33][128] = 16'b1111111111110000;
    assign weights1[33][129] = 16'b1111111111110110;
    assign weights1[33][130] = 16'b1111111111111110;
    assign weights1[33][131] = 16'b1111111111101111;
    assign weights1[33][132] = 16'b1111111111101010;
    assign weights1[33][133] = 16'b1111111111110101;
    assign weights1[33][134] = 16'b1111111111111110;
    assign weights1[33][135] = 16'b1111111111110001;
    assign weights1[33][136] = 16'b1111111111101000;
    assign weights1[33][137] = 16'b1111111111110100;
    assign weights1[33][138] = 16'b1111111111101100;
    assign weights1[33][139] = 16'b1111111111101001;
    assign weights1[33][140] = 16'b1111111111111000;
    assign weights1[33][141] = 16'b1111111111110010;
    assign weights1[33][142] = 16'b1111111111110101;
    assign weights1[33][143] = 16'b1111111111110111;
    assign weights1[33][144] = 16'b1111111111110010;
    assign weights1[33][145] = 16'b1111111111110110;
    assign weights1[33][146] = 16'b1111111111111111;
    assign weights1[33][147] = 16'b1111111111011011;
    assign weights1[33][148] = 16'b1111111111100101;
    assign weights1[33][149] = 16'b1111111111101110;
    assign weights1[33][150] = 16'b1111111111101111;
    assign weights1[33][151] = 16'b1111111111011010;
    assign weights1[33][152] = 16'b1111111111111011;
    assign weights1[33][153] = 16'b1111111111101111;
    assign weights1[33][154] = 16'b0000000000000001;
    assign weights1[33][155] = 16'b1111111111110111;
    assign weights1[33][156] = 16'b0000000000000111;
    assign weights1[33][157] = 16'b0000000000000001;
    assign weights1[33][158] = 16'b0000000000000111;
    assign weights1[33][159] = 16'b1111111111110011;
    assign weights1[33][160] = 16'b1111111111111101;
    assign weights1[33][161] = 16'b0000000000000010;
    assign weights1[33][162] = 16'b1111111111111000;
    assign weights1[33][163] = 16'b1111111111101100;
    assign weights1[33][164] = 16'b1111111111110011;
    assign weights1[33][165] = 16'b1111111111110100;
    assign weights1[33][166] = 16'b1111111111101110;
    assign weights1[33][167] = 16'b1111111111100101;
    assign weights1[33][168] = 16'b1111111111111000;
    assign weights1[33][169] = 16'b1111111111110011;
    assign weights1[33][170] = 16'b1111111111101001;
    assign weights1[33][171] = 16'b1111111111011111;
    assign weights1[33][172] = 16'b1111111111110011;
    assign weights1[33][173] = 16'b0000000000001110;
    assign weights1[33][174] = 16'b1111111111111010;
    assign weights1[33][175] = 16'b1111111111101100;
    assign weights1[33][176] = 16'b1111111111101011;
    assign weights1[33][177] = 16'b1111111111110101;
    assign weights1[33][178] = 16'b1111111111100111;
    assign weights1[33][179] = 16'b1111111111111000;
    assign weights1[33][180] = 16'b1111111111100001;
    assign weights1[33][181] = 16'b1111111111110011;
    assign weights1[33][182] = 16'b1111111111010001;
    assign weights1[33][183] = 16'b1111111111101001;
    assign weights1[33][184] = 16'b1111111111101110;
    assign weights1[33][185] = 16'b1111111111101000;
    assign weights1[33][186] = 16'b1111111111110010;
    assign weights1[33][187] = 16'b1111111111011100;
    assign weights1[33][188] = 16'b1111111111110111;
    assign weights1[33][189] = 16'b1111111111100001;
    assign weights1[33][190] = 16'b1111111111101101;
    assign weights1[33][191] = 16'b1111111111110001;
    assign weights1[33][192] = 16'b1111111111111000;
    assign weights1[33][193] = 16'b1111111111110100;
    assign weights1[33][194] = 16'b1111111111100100;
    assign weights1[33][195] = 16'b1111111111010001;
    assign weights1[33][196] = 16'b1111111111110011;
    assign weights1[33][197] = 16'b1111111111100101;
    assign weights1[33][198] = 16'b1111111111101001;
    assign weights1[33][199] = 16'b1111111111100101;
    assign weights1[33][200] = 16'b1111111111100111;
    assign weights1[33][201] = 16'b0000000000010001;
    assign weights1[33][202] = 16'b1111111111100110;
    assign weights1[33][203] = 16'b1111111111101110;
    assign weights1[33][204] = 16'b1111111111101000;
    assign weights1[33][205] = 16'b0000000000001010;
    assign weights1[33][206] = 16'b1111111111100011;
    assign weights1[33][207] = 16'b1111111111101101;
    assign weights1[33][208] = 16'b1111111111110001;
    assign weights1[33][209] = 16'b1111111111010011;
    assign weights1[33][210] = 16'b1111111111101110;
    assign weights1[33][211] = 16'b1111111111111100;
    assign weights1[33][212] = 16'b1111111111101011;
    assign weights1[33][213] = 16'b1111111111110110;
    assign weights1[33][214] = 16'b1111111111011001;
    assign weights1[33][215] = 16'b1111111111100101;
    assign weights1[33][216] = 16'b1111111111010010;
    assign weights1[33][217] = 16'b1111111111010010;
    assign weights1[33][218] = 16'b1111111111101111;
    assign weights1[33][219] = 16'b1111111111100000;
    assign weights1[33][220] = 16'b1111111111101011;
    assign weights1[33][221] = 16'b1111111111010111;
    assign weights1[33][222] = 16'b1111111111100001;
    assign weights1[33][223] = 16'b1111111111010100;
    assign weights1[33][224] = 16'b1111111111111000;
    assign weights1[33][225] = 16'b1111111111100110;
    assign weights1[33][226] = 16'b1111111111011010;
    assign weights1[33][227] = 16'b1111111111011110;
    assign weights1[33][228] = 16'b1111111111010110;
    assign weights1[33][229] = 16'b1111111111011000;
    assign weights1[33][230] = 16'b1111111111011110;
    assign weights1[33][231] = 16'b1111111111100100;
    assign weights1[33][232] = 16'b1111111111010110;
    assign weights1[33][233] = 16'b1111111111110001;
    assign weights1[33][234] = 16'b1111111111110010;
    assign weights1[33][235] = 16'b1111111111101011;
    assign weights1[33][236] = 16'b1111111111100100;
    assign weights1[33][237] = 16'b1111111111110000;
    assign weights1[33][238] = 16'b1111111111100010;
    assign weights1[33][239] = 16'b1111111111101100;
    assign weights1[33][240] = 16'b1111111111101011;
    assign weights1[33][241] = 16'b1111111111110000;
    assign weights1[33][242] = 16'b1111111111101111;
    assign weights1[33][243] = 16'b1111111111100010;
    assign weights1[33][244] = 16'b1111111111011110;
    assign weights1[33][245] = 16'b1111111111010101;
    assign weights1[33][246] = 16'b1111111111010011;
    assign weights1[33][247] = 16'b1111111111100110;
    assign weights1[33][248] = 16'b1111111111100111;
    assign weights1[33][249] = 16'b1111111111010110;
    assign weights1[33][250] = 16'b1111111111101000;
    assign weights1[33][251] = 16'b1111111111011011;
    assign weights1[33][252] = 16'b1111111111111010;
    assign weights1[33][253] = 16'b1111111111101111;
    assign weights1[33][254] = 16'b1111111111011000;
    assign weights1[33][255] = 16'b1111111111011010;
    assign weights1[33][256] = 16'b1111111111100101;
    assign weights1[33][257] = 16'b1111111111001101;
    assign weights1[33][258] = 16'b1111111111000001;
    assign weights1[33][259] = 16'b1111111111100001;
    assign weights1[33][260] = 16'b1111111111011010;
    assign weights1[33][261] = 16'b1111111111011010;
    assign weights1[33][262] = 16'b1111111111011111;
    assign weights1[33][263] = 16'b1111111111100101;
    assign weights1[33][264] = 16'b1111111111010101;
    assign weights1[33][265] = 16'b1111111111101000;
    assign weights1[33][266] = 16'b1111111111100010;
    assign weights1[33][267] = 16'b1111111111110100;
    assign weights1[33][268] = 16'b1111111111100011;
    assign weights1[33][269] = 16'b1111111111100110;
    assign weights1[33][270] = 16'b1111111111011111;
    assign weights1[33][271] = 16'b1111111111010111;
    assign weights1[33][272] = 16'b1111111111110000;
    assign weights1[33][273] = 16'b1111111111110110;
    assign weights1[33][274] = 16'b1111111111101011;
    assign weights1[33][275] = 16'b1111111111011010;
    assign weights1[33][276] = 16'b1111111111100100;
    assign weights1[33][277] = 16'b1111111111001010;
    assign weights1[33][278] = 16'b1111111111011101;
    assign weights1[33][279] = 16'b1111111111011011;
    assign weights1[33][280] = 16'b1111111111110100;
    assign weights1[33][281] = 16'b1111111111110001;
    assign weights1[33][282] = 16'b1111111111011101;
    assign weights1[33][283] = 16'b1111111111010101;
    assign weights1[33][284] = 16'b1111111111001011;
    assign weights1[33][285] = 16'b1111111111101111;
    assign weights1[33][286] = 16'b1111111111110011;
    assign weights1[33][287] = 16'b1111111111111011;
    assign weights1[33][288] = 16'b1111111111110001;
    assign weights1[33][289] = 16'b0000000000000000;
    assign weights1[33][290] = 16'b1111111111110000;
    assign weights1[33][291] = 16'b1111111111101111;
    assign weights1[33][292] = 16'b1111111111110011;
    assign weights1[33][293] = 16'b1111111111110010;
    assign weights1[33][294] = 16'b1111111111100111;
    assign weights1[33][295] = 16'b1111111111100110;
    assign weights1[33][296] = 16'b1111111111110011;
    assign weights1[33][297] = 16'b1111111111111011;
    assign weights1[33][298] = 16'b1111111111110111;
    assign weights1[33][299] = 16'b1111111111111010;
    assign weights1[33][300] = 16'b1111111111111000;
    assign weights1[33][301] = 16'b1111111111110111;
    assign weights1[33][302] = 16'b1111111111111110;
    assign weights1[33][303] = 16'b1111111111010111;
    assign weights1[33][304] = 16'b1111111111010111;
    assign weights1[33][305] = 16'b1111111111010000;
    assign weights1[33][306] = 16'b1111111111010110;
    assign weights1[33][307] = 16'b1111111111011000;
    assign weights1[33][308] = 16'b1111111111111100;
    assign weights1[33][309] = 16'b0000000000000100;
    assign weights1[33][310] = 16'b1111111111110001;
    assign weights1[33][311] = 16'b1111111111110000;
    assign weights1[33][312] = 16'b0000000000011110;
    assign weights1[33][313] = 16'b0000000000101100;
    assign weights1[33][314] = 16'b0000000000001101;
    assign weights1[33][315] = 16'b1111111111111101;
    assign weights1[33][316] = 16'b0000000000010000;
    assign weights1[33][317] = 16'b0000000000001100;
    assign weights1[33][318] = 16'b0000000000000101;
    assign weights1[33][319] = 16'b0000000000001010;
    assign weights1[33][320] = 16'b0000000000001000;
    assign weights1[33][321] = 16'b0000000000000001;
    assign weights1[33][322] = 16'b0000000000000010;
    assign weights1[33][323] = 16'b1111111111110111;
    assign weights1[33][324] = 16'b0000000000010000;
    assign weights1[33][325] = 16'b1111111111110000;
    assign weights1[33][326] = 16'b1111111111101101;
    assign weights1[33][327] = 16'b1111111111110110;
    assign weights1[33][328] = 16'b1111111111111001;
    assign weights1[33][329] = 16'b0000000000000011;
    assign weights1[33][330] = 16'b1111111111011100;
    assign weights1[33][331] = 16'b1111111111100100;
    assign weights1[33][332] = 16'b1111111111101110;
    assign weights1[33][333] = 16'b1111111111110110;
    assign weights1[33][334] = 16'b1111111111010011;
    assign weights1[33][335] = 16'b1111111111111010;
    assign weights1[33][336] = 16'b0000000000000110;
    assign weights1[33][337] = 16'b0000000000010001;
    assign weights1[33][338] = 16'b0000000000011001;
    assign weights1[33][339] = 16'b0000000000010000;
    assign weights1[33][340] = 16'b0000000000010111;
    assign weights1[33][341] = 16'b0000000000000111;
    assign weights1[33][342] = 16'b0000000000011101;
    assign weights1[33][343] = 16'b0000000000010111;
    assign weights1[33][344] = 16'b0000000001000000;
    assign weights1[33][345] = 16'b0000000000010101;
    assign weights1[33][346] = 16'b0000000000100101;
    assign weights1[33][347] = 16'b0000000000100010;
    assign weights1[33][348] = 16'b0000000000011001;
    assign weights1[33][349] = 16'b0000000000001000;
    assign weights1[33][350] = 16'b0000000000001000;
    assign weights1[33][351] = 16'b0000000000001011;
    assign weights1[33][352] = 16'b0000000000011100;
    assign weights1[33][353] = 16'b0000000000010000;
    assign weights1[33][354] = 16'b1111111111111111;
    assign weights1[33][355] = 16'b0000000000001000;
    assign weights1[33][356] = 16'b1111111111110000;
    assign weights1[33][357] = 16'b1111111111111011;
    assign weights1[33][358] = 16'b0000000000010100;
    assign weights1[33][359] = 16'b0000000000000110;
    assign weights1[33][360] = 16'b1111111111101000;
    assign weights1[33][361] = 16'b1111111111110101;
    assign weights1[33][362] = 16'b1111111111111011;
    assign weights1[33][363] = 16'b0000000000010111;
    assign weights1[33][364] = 16'b0000000000010101;
    assign weights1[33][365] = 16'b0000000000100100;
    assign weights1[33][366] = 16'b0000000000011111;
    assign weights1[33][367] = 16'b0000000000011111;
    assign weights1[33][368] = 16'b0000000000001011;
    assign weights1[33][369] = 16'b0000000000010011;
    assign weights1[33][370] = 16'b0000000000100001;
    assign weights1[33][371] = 16'b0000000000001011;
    assign weights1[33][372] = 16'b0000000000000000;
    assign weights1[33][373] = 16'b0000000000010101;
    assign weights1[33][374] = 16'b0000000000101010;
    assign weights1[33][375] = 16'b0000000000011001;
    assign weights1[33][376] = 16'b0000000000001100;
    assign weights1[33][377] = 16'b0000000000101010;
    assign weights1[33][378] = 16'b0000000000010110;
    assign weights1[33][379] = 16'b0000000000010100;
    assign weights1[33][380] = 16'b0000000000101100;
    assign weights1[33][381] = 16'b0000000000010111;
    assign weights1[33][382] = 16'b0000000000010011;
    assign weights1[33][383] = 16'b0000000000101000;
    assign weights1[33][384] = 16'b0000000000001011;
    assign weights1[33][385] = 16'b0000000000001110;
    assign weights1[33][386] = 16'b0000000000000100;
    assign weights1[33][387] = 16'b0000000000101001;
    assign weights1[33][388] = 16'b0000000000110111;
    assign weights1[33][389] = 16'b0000000000010001;
    assign weights1[33][390] = 16'b0000000000010000;
    assign weights1[33][391] = 16'b0000000000010011;
    assign weights1[33][392] = 16'b0000000000010000;
    assign weights1[33][393] = 16'b0000000000010100;
    assign weights1[33][394] = 16'b0000000000100001;
    assign weights1[33][395] = 16'b0000000000010001;
    assign weights1[33][396] = 16'b0000000000011001;
    assign weights1[33][397] = 16'b0000000000111001;
    assign weights1[33][398] = 16'b0000000000010000;
    assign weights1[33][399] = 16'b0000000000100011;
    assign weights1[33][400] = 16'b0000000000011001;
    assign weights1[33][401] = 16'b0000000000011111;
    assign weights1[33][402] = 16'b0000000000010011;
    assign weights1[33][403] = 16'b0000000000100100;
    assign weights1[33][404] = 16'b0000000000101000;
    assign weights1[33][405] = 16'b0000000000011001;
    assign weights1[33][406] = 16'b0000000000100000;
    assign weights1[33][407] = 16'b0000000000100001;
    assign weights1[33][408] = 16'b0000000000101101;
    assign weights1[33][409] = 16'b0000000000100001;
    assign weights1[33][410] = 16'b0000000000010011;
    assign weights1[33][411] = 16'b0000000000100111;
    assign weights1[33][412] = 16'b0000000000100001;
    assign weights1[33][413] = 16'b0000000000010111;
    assign weights1[33][414] = 16'b0000000000110000;
    assign weights1[33][415] = 16'b0000000000100111;
    assign weights1[33][416] = 16'b0000000000011010;
    assign weights1[33][417] = 16'b0000000000101111;
    assign weights1[33][418] = 16'b0000000000011111;
    assign weights1[33][419] = 16'b0000000000010000;
    assign weights1[33][420] = 16'b0000000000001111;
    assign weights1[33][421] = 16'b0000000000011101;
    assign weights1[33][422] = 16'b0000000000010011;
    assign weights1[33][423] = 16'b0000000000100011;
    assign weights1[33][424] = 16'b0000000000001010;
    assign weights1[33][425] = 16'b1111111111111100;
    assign weights1[33][426] = 16'b0000000000010111;
    assign weights1[33][427] = 16'b0000000000011001;
    assign weights1[33][428] = 16'b0000000000011010;
    assign weights1[33][429] = 16'b0000000000010110;
    assign weights1[33][430] = 16'b0000000000011001;
    assign weights1[33][431] = 16'b0000000000100001;
    assign weights1[33][432] = 16'b0000000000011010;
    assign weights1[33][433] = 16'b0000000000001001;
    assign weights1[33][434] = 16'b0000000000001011;
    assign weights1[33][435] = 16'b0000000000101001;
    assign weights1[33][436] = 16'b0000000000011010;
    assign weights1[33][437] = 16'b0000000000101001;
    assign weights1[33][438] = 16'b0000000000000110;
    assign weights1[33][439] = 16'b0000000000101101;
    assign weights1[33][440] = 16'b0000000000010000;
    assign weights1[33][441] = 16'b0000000000010011;
    assign weights1[33][442] = 16'b0000000000011110;
    assign weights1[33][443] = 16'b0000000000100100;
    assign weights1[33][444] = 16'b0000000000011001;
    assign weights1[33][445] = 16'b0000000000101101;
    assign weights1[33][446] = 16'b0000000001001011;
    assign weights1[33][447] = 16'b0000000000101000;
    assign weights1[33][448] = 16'b0000000000001101;
    assign weights1[33][449] = 16'b0000000000001101;
    assign weights1[33][450] = 16'b0000000000010001;
    assign weights1[33][451] = 16'b0000000000010011;
    assign weights1[33][452] = 16'b0000000000000110;
    assign weights1[33][453] = 16'b0000000000001111;
    assign weights1[33][454] = 16'b0000000000100000;
    assign weights1[33][455] = 16'b0000000000010001;
    assign weights1[33][456] = 16'b0000000000001100;
    assign weights1[33][457] = 16'b0000000000001000;
    assign weights1[33][458] = 16'b0000000000010000;
    assign weights1[33][459] = 16'b0000000000001110;
    assign weights1[33][460] = 16'b0000000000011101;
    assign weights1[33][461] = 16'b0000000000101001;
    assign weights1[33][462] = 16'b0000000000010111;
    assign weights1[33][463] = 16'b0000000000101101;
    assign weights1[33][464] = 16'b0000000000011110;
    assign weights1[33][465] = 16'b0000000000110111;
    assign weights1[33][466] = 16'b0000000000110011;
    assign weights1[33][467] = 16'b0000000000100000;
    assign weights1[33][468] = 16'b0000000000110000;
    assign weights1[33][469] = 16'b0000000000101001;
    assign weights1[33][470] = 16'b0000000000100111;
    assign weights1[33][471] = 16'b0000000000100110;
    assign weights1[33][472] = 16'b0000000000111011;
    assign weights1[33][473] = 16'b0000000000101101;
    assign weights1[33][474] = 16'b0000000000100100;
    assign weights1[33][475] = 16'b0000000000101101;
    assign weights1[33][476] = 16'b1111111111111100;
    assign weights1[33][477] = 16'b0000000000000000;
    assign weights1[33][478] = 16'b1111111111110111;
    assign weights1[33][479] = 16'b0000000000010100;
    assign weights1[33][480] = 16'b0000000000001011;
    assign weights1[33][481] = 16'b1111111111110100;
    assign weights1[33][482] = 16'b0000000000010101;
    assign weights1[33][483] = 16'b1111111111111100;
    assign weights1[33][484] = 16'b0000000000001101;
    assign weights1[33][485] = 16'b0000000000001010;
    assign weights1[33][486] = 16'b0000000000000011;
    assign weights1[33][487] = 16'b0000000000011101;
    assign weights1[33][488] = 16'b1111111111111001;
    assign weights1[33][489] = 16'b0000000000001110;
    assign weights1[33][490] = 16'b0000000000011010;
    assign weights1[33][491] = 16'b0000000000010011;
    assign weights1[33][492] = 16'b0000000000001011;
    assign weights1[33][493] = 16'b1111111111111101;
    assign weights1[33][494] = 16'b0000000000100011;
    assign weights1[33][495] = 16'b0000000000010000;
    assign weights1[33][496] = 16'b0000000000101001;
    assign weights1[33][497] = 16'b0000000000101100;
    assign weights1[33][498] = 16'b0000000000001110;
    assign weights1[33][499] = 16'b0000000000101100;
    assign weights1[33][500] = 16'b0000000000110110;
    assign weights1[33][501] = 16'b0000000000111010;
    assign weights1[33][502] = 16'b0000000000100011;
    assign weights1[33][503] = 16'b0000000000011010;
    assign weights1[33][504] = 16'b0000000000000001;
    assign weights1[33][505] = 16'b1111111111111100;
    assign weights1[33][506] = 16'b1111111111011011;
    assign weights1[33][507] = 16'b0000000000000100;
    assign weights1[33][508] = 16'b0000000000000000;
    assign weights1[33][509] = 16'b1111111111100111;
    assign weights1[33][510] = 16'b1111111111110111;
    assign weights1[33][511] = 16'b1111111111101111;
    assign weights1[33][512] = 16'b0000000000000100;
    assign weights1[33][513] = 16'b0000000000010000;
    assign weights1[33][514] = 16'b0000000000001100;
    assign weights1[33][515] = 16'b1111111111110011;
    assign weights1[33][516] = 16'b0000000000000011;
    assign weights1[33][517] = 16'b1111111111110111;
    assign weights1[33][518] = 16'b1111111111111110;
    assign weights1[33][519] = 16'b1111111111101111;
    assign weights1[33][520] = 16'b1111111111111101;
    assign weights1[33][521] = 16'b0000000000001000;
    assign weights1[33][522] = 16'b0000000000001100;
    assign weights1[33][523] = 16'b1111111111110011;
    assign weights1[33][524] = 16'b0000000000100110;
    assign weights1[33][525] = 16'b0000000000010010;
    assign weights1[33][526] = 16'b0000000000100010;
    assign weights1[33][527] = 16'b0000000000011110;
    assign weights1[33][528] = 16'b0000000000011000;
    assign weights1[33][529] = 16'b0000000000011010;
    assign weights1[33][530] = 16'b0000000000000110;
    assign weights1[33][531] = 16'b0000000000000111;
    assign weights1[33][532] = 16'b1111111111111001;
    assign weights1[33][533] = 16'b1111111111101110;
    assign weights1[33][534] = 16'b1111111111100110;
    assign weights1[33][535] = 16'b1111111111100100;
    assign weights1[33][536] = 16'b0000000000000110;
    assign weights1[33][537] = 16'b1111111111011111;
    assign weights1[33][538] = 16'b0000000000000100;
    assign weights1[33][539] = 16'b0000000000001111;
    assign weights1[33][540] = 16'b1111111111101111;
    assign weights1[33][541] = 16'b1111111111100000;
    assign weights1[33][542] = 16'b1111111111111100;
    assign weights1[33][543] = 16'b0000000000000001;
    assign weights1[33][544] = 16'b1111111111111110;
    assign weights1[33][545] = 16'b1111111111101111;
    assign weights1[33][546] = 16'b1111111111101001;
    assign weights1[33][547] = 16'b1111111111111000;
    assign weights1[33][548] = 16'b1111111111110110;
    assign weights1[33][549] = 16'b1111111111110100;
    assign weights1[33][550] = 16'b1111111111100110;
    assign weights1[33][551] = 16'b1111111111100101;
    assign weights1[33][552] = 16'b1111111111111110;
    assign weights1[33][553] = 16'b0000000000000101;
    assign weights1[33][554] = 16'b0000000000000000;
    assign weights1[33][555] = 16'b0000000000010100;
    assign weights1[33][556] = 16'b0000000000010010;
    assign weights1[33][557] = 16'b1111111111100001;
    assign weights1[33][558] = 16'b1111111111111101;
    assign weights1[33][559] = 16'b1111111111111111;
    assign weights1[33][560] = 16'b1111111111110111;
    assign weights1[33][561] = 16'b1111111111011101;
    assign weights1[33][562] = 16'b1111111111011010;
    assign weights1[33][563] = 16'b1111111111001011;
    assign weights1[33][564] = 16'b1111111111101010;
    assign weights1[33][565] = 16'b1111111111100011;
    assign weights1[33][566] = 16'b1111111111111010;
    assign weights1[33][567] = 16'b0000000000000100;
    assign weights1[33][568] = 16'b0000000000000011;
    assign weights1[33][569] = 16'b1111111111111000;
    assign weights1[33][570] = 16'b1111111111110011;
    assign weights1[33][571] = 16'b1111111111111111;
    assign weights1[33][572] = 16'b0000000000000011;
    assign weights1[33][573] = 16'b0000000000000110;
    assign weights1[33][574] = 16'b1111111111111010;
    assign weights1[33][575] = 16'b0000000000001100;
    assign weights1[33][576] = 16'b1111111111110100;
    assign weights1[33][577] = 16'b1111111111111001;
    assign weights1[33][578] = 16'b1111111111111001;
    assign weights1[33][579] = 16'b1111111111100011;
    assign weights1[33][580] = 16'b1111111111011001;
    assign weights1[33][581] = 16'b1111111111100010;
    assign weights1[33][582] = 16'b1111111111100110;
    assign weights1[33][583] = 16'b1111111111100001;
    assign weights1[33][584] = 16'b1111111111010010;
    assign weights1[33][585] = 16'b1111111111000000;
    assign weights1[33][586] = 16'b1111111111010010;
    assign weights1[33][587] = 16'b1111111111011110;
    assign weights1[33][588] = 16'b1111111111111100;
    assign weights1[33][589] = 16'b1111111111110101;
    assign weights1[33][590] = 16'b1111111111100110;
    assign weights1[33][591] = 16'b1111111111001001;
    assign weights1[33][592] = 16'b1111111111000101;
    assign weights1[33][593] = 16'b1111111111000101;
    assign weights1[33][594] = 16'b1111111111011100;
    assign weights1[33][595] = 16'b1111111111110011;
    assign weights1[33][596] = 16'b1111111111111010;
    assign weights1[33][597] = 16'b1111111111100110;
    assign weights1[33][598] = 16'b1111111111111000;
    assign weights1[33][599] = 16'b1111111111110111;
    assign weights1[33][600] = 16'b0000000000100111;
    assign weights1[33][601] = 16'b0000000000010101;
    assign weights1[33][602] = 16'b0000000000000100;
    assign weights1[33][603] = 16'b1111111111111011;
    assign weights1[33][604] = 16'b1111111111011110;
    assign weights1[33][605] = 16'b1111111111111011;
    assign weights1[33][606] = 16'b1111111111110000;
    assign weights1[33][607] = 16'b1111111111100101;
    assign weights1[33][608] = 16'b1111111111010111;
    assign weights1[33][609] = 16'b1111111111010011;
    assign weights1[33][610] = 16'b1111111110111101;
    assign weights1[33][611] = 16'b1111111110111110;
    assign weights1[33][612] = 16'b1111111110100111;
    assign weights1[33][613] = 16'b1111111110110111;
    assign weights1[33][614] = 16'b1111111111000100;
    assign weights1[33][615] = 16'b1111111111011001;
    assign weights1[33][616] = 16'b1111111111111001;
    assign weights1[33][617] = 16'b1111111111111000;
    assign weights1[33][618] = 16'b1111111111101100;
    assign weights1[33][619] = 16'b1111111111011001;
    assign weights1[33][620] = 16'b1111111111010000;
    assign weights1[33][621] = 16'b1111111111000010;
    assign weights1[33][622] = 16'b1111111111001110;
    assign weights1[33][623] = 16'b1111111110111101;
    assign weights1[33][624] = 16'b1111111111011001;
    assign weights1[33][625] = 16'b1111111111001010;
    assign weights1[33][626] = 16'b0000000000000000;
    assign weights1[33][627] = 16'b1111111111100001;
    assign weights1[33][628] = 16'b1111111111100011;
    assign weights1[33][629] = 16'b1111111111101001;
    assign weights1[33][630] = 16'b1111111111100001;
    assign weights1[33][631] = 16'b1111111111101000;
    assign weights1[33][632] = 16'b1111111111110011;
    assign weights1[33][633] = 16'b1111111111100001;
    assign weights1[33][634] = 16'b1111111111110100;
    assign weights1[33][635] = 16'b1111111111011000;
    assign weights1[33][636] = 16'b1111111111010111;
    assign weights1[33][637] = 16'b1111111111000111;
    assign weights1[33][638] = 16'b1111111110110000;
    assign weights1[33][639] = 16'b1111111110100101;
    assign weights1[33][640] = 16'b1111111110101000;
    assign weights1[33][641] = 16'b1111111110111111;
    assign weights1[33][642] = 16'b1111111111010100;
    assign weights1[33][643] = 16'b1111111111011010;
    assign weights1[33][644] = 16'b1111111111111011;
    assign weights1[33][645] = 16'b1111111111110011;
    assign weights1[33][646] = 16'b1111111111101100;
    assign weights1[33][647] = 16'b1111111111010111;
    assign weights1[33][648] = 16'b1111111111000100;
    assign weights1[33][649] = 16'b1111111110111011;
    assign weights1[33][650] = 16'b1111111110111001;
    assign weights1[33][651] = 16'b1111111110100011;
    assign weights1[33][652] = 16'b1111111110110100;
    assign weights1[33][653] = 16'b1111111110001110;
    assign weights1[33][654] = 16'b1111111110101101;
    assign weights1[33][655] = 16'b1111111110100101;
    assign weights1[33][656] = 16'b1111111110111001;
    assign weights1[33][657] = 16'b1111111111010011;
    assign weights1[33][658] = 16'b1111111111001001;
    assign weights1[33][659] = 16'b1111111111101000;
    assign weights1[33][660] = 16'b1111111111011000;
    assign weights1[33][661] = 16'b1111111111001110;
    assign weights1[33][662] = 16'b1111111111011001;
    assign weights1[33][663] = 16'b1111111111011101;
    assign weights1[33][664] = 16'b1111111111011001;
    assign weights1[33][665] = 16'b1111111110110110;
    assign weights1[33][666] = 16'b1111111111000010;
    assign weights1[33][667] = 16'b1111111110110111;
    assign weights1[33][668] = 16'b1111111110110111;
    assign weights1[33][669] = 16'b1111111111010000;
    assign weights1[33][670] = 16'b1111111111100010;
    assign weights1[33][671] = 16'b1111111111100110;
    assign weights1[33][672] = 16'b1111111111111101;
    assign weights1[33][673] = 16'b1111111111110110;
    assign weights1[33][674] = 16'b1111111111100101;
    assign weights1[33][675] = 16'b1111111111011000;
    assign weights1[33][676] = 16'b1111111111010101;
    assign weights1[33][677] = 16'b1111111111001101;
    assign weights1[33][678] = 16'b1111111111000001;
    assign weights1[33][679] = 16'b1111111110110111;
    assign weights1[33][680] = 16'b1111111110110100;
    assign weights1[33][681] = 16'b1111111111000101;
    assign weights1[33][682] = 16'b1111111110101000;
    assign weights1[33][683] = 16'b1111111111010101;
    assign weights1[33][684] = 16'b1111111111000111;
    assign weights1[33][685] = 16'b1111111110110110;
    assign weights1[33][686] = 16'b1111111111011110;
    assign weights1[33][687] = 16'b1111111111011001;
    assign weights1[33][688] = 16'b1111111111010101;
    assign weights1[33][689] = 16'b1111111111010000;
    assign weights1[33][690] = 16'b1111111111011100;
    assign weights1[33][691] = 16'b1111111111000111;
    assign weights1[33][692] = 16'b1111111110100111;
    assign weights1[33][693] = 16'b1111111110111110;
    assign weights1[33][694] = 16'b1111111110111111;
    assign weights1[33][695] = 16'b1111111111010011;
    assign weights1[33][696] = 16'b1111111111010101;
    assign weights1[33][697] = 16'b1111111111011101;
    assign weights1[33][698] = 16'b1111111111100001;
    assign weights1[33][699] = 16'b1111111111100111;
    assign weights1[33][700] = 16'b0000000000000000;
    assign weights1[33][701] = 16'b1111111111110101;
    assign weights1[33][702] = 16'b1111111111100111;
    assign weights1[33][703] = 16'b1111111111100011;
    assign weights1[33][704] = 16'b1111111111100000;
    assign weights1[33][705] = 16'b1111111111010000;
    assign weights1[33][706] = 16'b1111111111000100;
    assign weights1[33][707] = 16'b1111111111000011;
    assign weights1[33][708] = 16'b1111111110111111;
    assign weights1[33][709] = 16'b1111111110011100;
    assign weights1[33][710] = 16'b1111111110011101;
    assign weights1[33][711] = 16'b1111111110100110;
    assign weights1[33][712] = 16'b1111111110001001;
    assign weights1[33][713] = 16'b1111111110010000;
    assign weights1[33][714] = 16'b1111111110101101;
    assign weights1[33][715] = 16'b1111111110010101;
    assign weights1[33][716] = 16'b1111111110010100;
    assign weights1[33][717] = 16'b1111111110011001;
    assign weights1[33][718] = 16'b1111111110000100;
    assign weights1[33][719] = 16'b1111111110010100;
    assign weights1[33][720] = 16'b1111111110010111;
    assign weights1[33][721] = 16'b1111111110110011;
    assign weights1[33][722] = 16'b1111111110111101;
    assign weights1[33][723] = 16'b1111111111010100;
    assign weights1[33][724] = 16'b1111111111011000;
    assign weights1[33][725] = 16'b1111111111100101;
    assign weights1[33][726] = 16'b1111111111101000;
    assign weights1[33][727] = 16'b1111111111110001;
    assign weights1[33][728] = 16'b1111111111111110;
    assign weights1[33][729] = 16'b1111111111111001;
    assign weights1[33][730] = 16'b1111111111110011;
    assign weights1[33][731] = 16'b1111111111110000;
    assign weights1[33][732] = 16'b1111111111101000;
    assign weights1[33][733] = 16'b1111111111011000;
    assign weights1[33][734] = 16'b1111111111001010;
    assign weights1[33][735] = 16'b1111111111000001;
    assign weights1[33][736] = 16'b1111111110111111;
    assign weights1[33][737] = 16'b1111111110111010;
    assign weights1[33][738] = 16'b1111111110110000;
    assign weights1[33][739] = 16'b1111111110011110;
    assign weights1[33][740] = 16'b1111111110011001;
    assign weights1[33][741] = 16'b1111111110001010;
    assign weights1[33][742] = 16'b1111111110001001;
    assign weights1[33][743] = 16'b1111111110010000;
    assign weights1[33][744] = 16'b1111111110011100;
    assign weights1[33][745] = 16'b1111111110010010;
    assign weights1[33][746] = 16'b1111111110101000;
    assign weights1[33][747] = 16'b1111111110101110;
    assign weights1[33][748] = 16'b1111111110110001;
    assign weights1[33][749] = 16'b1111111111000110;
    assign weights1[33][750] = 16'b1111111111010001;
    assign weights1[33][751] = 16'b1111111111100010;
    assign weights1[33][752] = 16'b1111111111100101;
    assign weights1[33][753] = 16'b1111111111101001;
    assign weights1[33][754] = 16'b1111111111110000;
    assign weights1[33][755] = 16'b1111111111110111;
    assign weights1[33][756] = 16'b1111111111111011;
    assign weights1[33][757] = 16'b1111111111111010;
    assign weights1[33][758] = 16'b1111111111111010;
    assign weights1[33][759] = 16'b1111111111111001;
    assign weights1[33][760] = 16'b1111111111110000;
    assign weights1[33][761] = 16'b1111111111101000;
    assign weights1[33][762] = 16'b1111111111100001;
    assign weights1[33][763] = 16'b1111111111001101;
    assign weights1[33][764] = 16'b1111111111001000;
    assign weights1[33][765] = 16'b1111111111001101;
    assign weights1[33][766] = 16'b1111111111000101;
    assign weights1[33][767] = 16'b1111111110110010;
    assign weights1[33][768] = 16'b1111111110110011;
    assign weights1[33][769] = 16'b1111111110110000;
    assign weights1[33][770] = 16'b1111111110100110;
    assign weights1[33][771] = 16'b1111111110111000;
    assign weights1[33][772] = 16'b1111111110111101;
    assign weights1[33][773] = 16'b1111111110111101;
    assign weights1[33][774] = 16'b1111111111000101;
    assign weights1[33][775] = 16'b1111111111001101;
    assign weights1[33][776] = 16'b1111111111010001;
    assign weights1[33][777] = 16'b1111111111010110;
    assign weights1[33][778] = 16'b1111111111100100;
    assign weights1[33][779] = 16'b1111111111101101;
    assign weights1[33][780] = 16'b1111111111101101;
    assign weights1[33][781] = 16'b1111111111110100;
    assign weights1[33][782] = 16'b1111111111111001;
    assign weights1[33][783] = 16'b1111111111111100;
    assign weights1[34][0] = 16'b0000000000000001;
    assign weights1[34][1] = 16'b1111111111111111;
    assign weights1[34][2] = 16'b1111111111111110;
    assign weights1[34][3] = 16'b0000000000000001;
    assign weights1[34][4] = 16'b0000000000000011;
    assign weights1[34][5] = 16'b0000000000001000;
    assign weights1[34][6] = 16'b0000000000000001;
    assign weights1[34][7] = 16'b0000000000001101;
    assign weights1[34][8] = 16'b0000000000010110;
    assign weights1[34][9] = 16'b0000000000001110;
    assign weights1[34][10] = 16'b0000000000000111;
    assign weights1[34][11] = 16'b0000000000000101;
    assign weights1[34][12] = 16'b1111111111110011;
    assign weights1[34][13] = 16'b1111111111011000;
    assign weights1[34][14] = 16'b1111111111000001;
    assign weights1[34][15] = 16'b1111111111000011;
    assign weights1[34][16] = 16'b1111111111010110;
    assign weights1[34][17] = 16'b1111111111011101;
    assign weights1[34][18] = 16'b1111111111110100;
    assign weights1[34][19] = 16'b1111111111111110;
    assign weights1[34][20] = 16'b0000000000010000;
    assign weights1[34][21] = 16'b0000000000011000;
    assign weights1[34][22] = 16'b0000000000010000;
    assign weights1[34][23] = 16'b0000000000010010;
    assign weights1[34][24] = 16'b0000000000001010;
    assign weights1[34][25] = 16'b0000000000000010;
    assign weights1[34][26] = 16'b0000000000000110;
    assign weights1[34][27] = 16'b0000000000000001;
    assign weights1[34][28] = 16'b1111111111111110;
    assign weights1[34][29] = 16'b1111111111111110;
    assign weights1[34][30] = 16'b0000000000000001;
    assign weights1[34][31] = 16'b0000000000000010;
    assign weights1[34][32] = 16'b0000000000000101;
    assign weights1[34][33] = 16'b0000000000000010;
    assign weights1[34][34] = 16'b1111111111111110;
    assign weights1[34][35] = 16'b0000000000010101;
    assign weights1[34][36] = 16'b0000000000100001;
    assign weights1[34][37] = 16'b0000000000001001;
    assign weights1[34][38] = 16'b0000000000010011;
    assign weights1[34][39] = 16'b0000000000001101;
    assign weights1[34][40] = 16'b0000000000010001;
    assign weights1[34][41] = 16'b1111111111100110;
    assign weights1[34][42] = 16'b1111111111001101;
    assign weights1[34][43] = 16'b1111111111000010;
    assign weights1[34][44] = 16'b1111111111001001;
    assign weights1[34][45] = 16'b1111111111011011;
    assign weights1[34][46] = 16'b1111111111011111;
    assign weights1[34][47] = 16'b0000000000010001;
    assign weights1[34][48] = 16'b0000000000011111;
    assign weights1[34][49] = 16'b0000000000011011;
    assign weights1[34][50] = 16'b0000000000010101;
    assign weights1[34][51] = 16'b0000000000010100;
    assign weights1[34][52] = 16'b0000000000001100;
    assign weights1[34][53] = 16'b0000000000010001;
    assign weights1[34][54] = 16'b0000000000001111;
    assign weights1[34][55] = 16'b0000000000001001;
    assign weights1[34][56] = 16'b0000000000000010;
    assign weights1[34][57] = 16'b0000000000000010;
    assign weights1[34][58] = 16'b0000000000000010;
    assign weights1[34][59] = 16'b0000000000000010;
    assign weights1[34][60] = 16'b0000000000000100;
    assign weights1[34][61] = 16'b1111111111111101;
    assign weights1[34][62] = 16'b1111111111110010;
    assign weights1[34][63] = 16'b0000000000000000;
    assign weights1[34][64] = 16'b0000000000011001;
    assign weights1[34][65] = 16'b0000000000001100;
    assign weights1[34][66] = 16'b1111111111110011;
    assign weights1[34][67] = 16'b0000000000000011;
    assign weights1[34][68] = 16'b0000000000000110;
    assign weights1[34][69] = 16'b1111111111010101;
    assign weights1[34][70] = 16'b1111111111000001;
    assign weights1[34][71] = 16'b1111111110101111;
    assign weights1[34][72] = 16'b1111111110101101;
    assign weights1[34][73] = 16'b1111111110111001;
    assign weights1[34][74] = 16'b1111111111010000;
    assign weights1[34][75] = 16'b0000000000000101;
    assign weights1[34][76] = 16'b0000000000101100;
    assign weights1[34][77] = 16'b0000000000100100;
    assign weights1[34][78] = 16'b0000000000011100;
    assign weights1[34][79] = 16'b0000000000100000;
    assign weights1[34][80] = 16'b0000000000010010;
    assign weights1[34][81] = 16'b0000000000010000;
    assign weights1[34][82] = 16'b0000000000010000;
    assign weights1[34][83] = 16'b0000000000001010;
    assign weights1[34][84] = 16'b0000000000000110;
    assign weights1[34][85] = 16'b0000000000001001;
    assign weights1[34][86] = 16'b0000000000000010;
    assign weights1[34][87] = 16'b0000000000000101;
    assign weights1[34][88] = 16'b0000000000000100;
    assign weights1[34][89] = 16'b1111111111101111;
    assign weights1[34][90] = 16'b1111111111111001;
    assign weights1[34][91] = 16'b0000000000001011;
    assign weights1[34][92] = 16'b0000000000010010;
    assign weights1[34][93] = 16'b0000000000000111;
    assign weights1[34][94] = 16'b1111111111111001;
    assign weights1[34][95] = 16'b1111111111110101;
    assign weights1[34][96] = 16'b1111111111110101;
    assign weights1[34][97] = 16'b1111111111001110;
    assign weights1[34][98] = 16'b1111111111010000;
    assign weights1[34][99] = 16'b1111111110101011;
    assign weights1[34][100] = 16'b1111111110000001;
    assign weights1[34][101] = 16'b1111111110100110;
    assign weights1[34][102] = 16'b1111111111001101;
    assign weights1[34][103] = 16'b1111111111111100;
    assign weights1[34][104] = 16'b0000000000010110;
    assign weights1[34][105] = 16'b0000000000000101;
    assign weights1[34][106] = 16'b0000000000010010;
    assign weights1[34][107] = 16'b0000000000011000;
    assign weights1[34][108] = 16'b0000000000011101;
    assign weights1[34][109] = 16'b0000000000010000;
    assign weights1[34][110] = 16'b0000000000001111;
    assign weights1[34][111] = 16'b0000000000001001;
    assign weights1[34][112] = 16'b0000000000000100;
    assign weights1[34][113] = 16'b0000000000000011;
    assign weights1[34][114] = 16'b1111111111111011;
    assign weights1[34][115] = 16'b1111111111111100;
    assign weights1[34][116] = 16'b1111111111111010;
    assign weights1[34][117] = 16'b1111111111110111;
    assign weights1[34][118] = 16'b1111111111111001;
    assign weights1[34][119] = 16'b1111111111111100;
    assign weights1[34][120] = 16'b0000000000001000;
    assign weights1[34][121] = 16'b0000000000011001;
    assign weights1[34][122] = 16'b1111111111110001;
    assign weights1[34][123] = 16'b0000000000000100;
    assign weights1[34][124] = 16'b1111111111111111;
    assign weights1[34][125] = 16'b1111111111010010;
    assign weights1[34][126] = 16'b1111111111011111;
    assign weights1[34][127] = 16'b1111111110100011;
    assign weights1[34][128] = 16'b1111111101101101;
    assign weights1[34][129] = 16'b1111111110000001;
    assign weights1[34][130] = 16'b1111111110111100;
    assign weights1[34][131] = 16'b1111111111100101;
    assign weights1[34][132] = 16'b0000000000010110;
    assign weights1[34][133] = 16'b0000000000010101;
    assign weights1[34][134] = 16'b0000000000011011;
    assign weights1[34][135] = 16'b0000000000100001;
    assign weights1[34][136] = 16'b0000000000101001;
    assign weights1[34][137] = 16'b0000000000001001;
    assign weights1[34][138] = 16'b0000000000000110;
    assign weights1[34][139] = 16'b0000000000001100;
    assign weights1[34][140] = 16'b0000000000000101;
    assign weights1[34][141] = 16'b1111111111111101;
    assign weights1[34][142] = 16'b1111111111111100;
    assign weights1[34][143] = 16'b1111111111111000;
    assign weights1[34][144] = 16'b1111111111101000;
    assign weights1[34][145] = 16'b1111111111111010;
    assign weights1[34][146] = 16'b1111111111101111;
    assign weights1[34][147] = 16'b0000000000000000;
    assign weights1[34][148] = 16'b0000000000001110;
    assign weights1[34][149] = 16'b1111111111111000;
    assign weights1[34][150] = 16'b0000000000000001;
    assign weights1[34][151] = 16'b1111111111111011;
    assign weights1[34][152] = 16'b0000000000001101;
    assign weights1[34][153] = 16'b1111111111110101;
    assign weights1[34][154] = 16'b1111111111010101;
    assign weights1[34][155] = 16'b1111111110111001;
    assign weights1[34][156] = 16'b1111111101011101;
    assign weights1[34][157] = 16'b1111111101010011;
    assign weights1[34][158] = 16'b1111111111100110;
    assign weights1[34][159] = 16'b0000000000010000;
    assign weights1[34][160] = 16'b0000000000011001;
    assign weights1[34][161] = 16'b0000000000101001;
    assign weights1[34][162] = 16'b0000000000011111;
    assign weights1[34][163] = 16'b0000000000101101;
    assign weights1[34][164] = 16'b0000000000001111;
    assign weights1[34][165] = 16'b0000000000001001;
    assign weights1[34][166] = 16'b0000000000000001;
    assign weights1[34][167] = 16'b1111111111111111;
    assign weights1[34][168] = 16'b0000000000000011;
    assign weights1[34][169] = 16'b0000000000000010;
    assign weights1[34][170] = 16'b1111111111110111;
    assign weights1[34][171] = 16'b1111111111111001;
    assign weights1[34][172] = 16'b1111111111111101;
    assign weights1[34][173] = 16'b0000000000000000;
    assign weights1[34][174] = 16'b0000000000000010;
    assign weights1[34][175] = 16'b0000000000000010;
    assign weights1[34][176] = 16'b0000000000001001;
    assign weights1[34][177] = 16'b0000000000010010;
    assign weights1[34][178] = 16'b0000000000000111;
    assign weights1[34][179] = 16'b1111111111111001;
    assign weights1[34][180] = 16'b1111111111111001;
    assign weights1[34][181] = 16'b1111111111101010;
    assign weights1[34][182] = 16'b1111111111111110;
    assign weights1[34][183] = 16'b1111111111000111;
    assign weights1[34][184] = 16'b1111111100110001;
    assign weights1[34][185] = 16'b1111111101000100;
    assign weights1[34][186] = 16'b1111111111011111;
    assign weights1[34][187] = 16'b0000000000111001;
    assign weights1[34][188] = 16'b0000000000010011;
    assign weights1[34][189] = 16'b0000000000010000;
    assign weights1[34][190] = 16'b0000000000011001;
    assign weights1[34][191] = 16'b0000000000100010;
    assign weights1[34][192] = 16'b0000000000010001;
    assign weights1[34][193] = 16'b1111111111111101;
    assign weights1[34][194] = 16'b1111111111111001;
    assign weights1[34][195] = 16'b1111111111111101;
    assign weights1[34][196] = 16'b0000000000001000;
    assign weights1[34][197] = 16'b0000000000000110;
    assign weights1[34][198] = 16'b1111111111111100;
    assign weights1[34][199] = 16'b1111111111110110;
    assign weights1[34][200] = 16'b1111111111111101;
    assign weights1[34][201] = 16'b1111111111100101;
    assign weights1[34][202] = 16'b1111111111101110;
    assign weights1[34][203] = 16'b1111111111111110;
    assign weights1[34][204] = 16'b0000000000010111;
    assign weights1[34][205] = 16'b0000000000001100;
    assign weights1[34][206] = 16'b0000000000010011;
    assign weights1[34][207] = 16'b0000000000000000;
    assign weights1[34][208] = 16'b0000000000001101;
    assign weights1[34][209] = 16'b1111111111111111;
    assign weights1[34][210] = 16'b1111111111110100;
    assign weights1[34][211] = 16'b1111111111100001;
    assign weights1[34][212] = 16'b1111111100001100;
    assign weights1[34][213] = 16'b1111111100110111;
    assign weights1[34][214] = 16'b0000000000100111;
    assign weights1[34][215] = 16'b0000000001000110;
    assign weights1[34][216] = 16'b0000000000100110;
    assign weights1[34][217] = 16'b0000000000010001;
    assign weights1[34][218] = 16'b0000000000011101;
    assign weights1[34][219] = 16'b0000000000101110;
    assign weights1[34][220] = 16'b0000000000001010;
    assign weights1[34][221] = 16'b1111111111101100;
    assign weights1[34][222] = 16'b1111111111101001;
    assign weights1[34][223] = 16'b1111111111101101;
    assign weights1[34][224] = 16'b0000000000000011;
    assign weights1[34][225] = 16'b1111111111111111;
    assign weights1[34][226] = 16'b0000000000000011;
    assign weights1[34][227] = 16'b1111111111111101;
    assign weights1[34][228] = 16'b1111111111110100;
    assign weights1[34][229] = 16'b1111111111100110;
    assign weights1[34][230] = 16'b1111111111100000;
    assign weights1[34][231] = 16'b1111111111110111;
    assign weights1[34][232] = 16'b1111111111100101;
    assign weights1[34][233] = 16'b0000000000000111;
    assign weights1[34][234] = 16'b0000000000100010;
    assign weights1[34][235] = 16'b0000000000001110;
    assign weights1[34][236] = 16'b0000000000101000;
    assign weights1[34][237] = 16'b0000000000001000;
    assign weights1[34][238] = 16'b1111111111101110;
    assign weights1[34][239] = 16'b1111111110101011;
    assign weights1[34][240] = 16'b1111111011111011;
    assign weights1[34][241] = 16'b1111111110100101;
    assign weights1[34][242] = 16'b0000000000111000;
    assign weights1[34][243] = 16'b0000000000100000;
    assign weights1[34][244] = 16'b0000000000011110;
    assign weights1[34][245] = 16'b1111111111100110;
    assign weights1[34][246] = 16'b0000000000100010;
    assign weights1[34][247] = 16'b0000000000100011;
    assign weights1[34][248] = 16'b1111111111101111;
    assign weights1[34][249] = 16'b1111111111111001;
    assign weights1[34][250] = 16'b1111111111001000;
    assign weights1[34][251] = 16'b1111111111011111;
    assign weights1[34][252] = 16'b0000000000000110;
    assign weights1[34][253] = 16'b1111111111111111;
    assign weights1[34][254] = 16'b0000000000010001;
    assign weights1[34][255] = 16'b0000000000000001;
    assign weights1[34][256] = 16'b1111111111110000;
    assign weights1[34][257] = 16'b1111111111111101;
    assign weights1[34][258] = 16'b1111111111101100;
    assign weights1[34][259] = 16'b1111111111110100;
    assign weights1[34][260] = 16'b0000000000000111;
    assign weights1[34][261] = 16'b1111111111111110;
    assign weights1[34][262] = 16'b0000000000000100;
    assign weights1[34][263] = 16'b0000000000010110;
    assign weights1[34][264] = 16'b0000000000011110;
    assign weights1[34][265] = 16'b0000000000100100;
    assign weights1[34][266] = 16'b1111111111101110;
    assign weights1[34][267] = 16'b1111111101101100;
    assign weights1[34][268] = 16'b1111111011110011;
    assign weights1[34][269] = 16'b1111111111111001;
    assign weights1[34][270] = 16'b0000000000101111;
    assign weights1[34][271] = 16'b0000000000000101;
    assign weights1[34][272] = 16'b0000000000100010;
    assign weights1[34][273] = 16'b0000000000001000;
    assign weights1[34][274] = 16'b0000000000010010;
    assign weights1[34][275] = 16'b0000000000000011;
    assign weights1[34][276] = 16'b1111111111110111;
    assign weights1[34][277] = 16'b1111111111011001;
    assign weights1[34][278] = 16'b1111111111010011;
    assign weights1[34][279] = 16'b1111111111100001;
    assign weights1[34][280] = 16'b0000000000000101;
    assign weights1[34][281] = 16'b0000000000000111;
    assign weights1[34][282] = 16'b0000000000000001;
    assign weights1[34][283] = 16'b1111111111111001;
    assign weights1[34][284] = 16'b1111111111110000;
    assign weights1[34][285] = 16'b1111111111110111;
    assign weights1[34][286] = 16'b1111111111101001;
    assign weights1[34][287] = 16'b0000000000000011;
    assign weights1[34][288] = 16'b0000000000001111;
    assign weights1[34][289] = 16'b0000000000010000;
    assign weights1[34][290] = 16'b0000000000001101;
    assign weights1[34][291] = 16'b0000000000011000;
    assign weights1[34][292] = 16'b0000000000100011;
    assign weights1[34][293] = 16'b0000000000100110;
    assign weights1[34][294] = 16'b1111111111111110;
    assign weights1[34][295] = 16'b1111111101010100;
    assign weights1[34][296] = 16'b1111111101011111;
    assign weights1[34][297] = 16'b0000000000001111;
    assign weights1[34][298] = 16'b0000000000010000;
    assign weights1[34][299] = 16'b0000000000010011;
    assign weights1[34][300] = 16'b0000000000010011;
    assign weights1[34][301] = 16'b0000000000001111;
    assign weights1[34][302] = 16'b0000000000000111;
    assign weights1[34][303] = 16'b0000000000000000;
    assign weights1[34][304] = 16'b1111111111110011;
    assign weights1[34][305] = 16'b1111111111011011;
    assign weights1[34][306] = 16'b1111111111010101;
    assign weights1[34][307] = 16'b1111111111100100;
    assign weights1[34][308] = 16'b0000000000000010;
    assign weights1[34][309] = 16'b0000000000001010;
    assign weights1[34][310] = 16'b1111111111111001;
    assign weights1[34][311] = 16'b1111111111110100;
    assign weights1[34][312] = 16'b1111111111011010;
    assign weights1[34][313] = 16'b1111111111110011;
    assign weights1[34][314] = 16'b1111111111110101;
    assign weights1[34][315] = 16'b0000000000000000;
    assign weights1[34][316] = 16'b1111111111110010;
    assign weights1[34][317] = 16'b0000000000000000;
    assign weights1[34][318] = 16'b0000000000010111;
    assign weights1[34][319] = 16'b0000000000001110;
    assign weights1[34][320] = 16'b0000000000110100;
    assign weights1[34][321] = 16'b0000000000010100;
    assign weights1[34][322] = 16'b1111111111010100;
    assign weights1[34][323] = 16'b1111111101111101;
    assign weights1[34][324] = 16'b1111111110100000;
    assign weights1[34][325] = 16'b1111111111110110;
    assign weights1[34][326] = 16'b0000000000101011;
    assign weights1[34][327] = 16'b0000000000001101;
    assign weights1[34][328] = 16'b0000000000000000;
    assign weights1[34][329] = 16'b0000000000010111;
    assign weights1[34][330] = 16'b0000000000001110;
    assign weights1[34][331] = 16'b0000000000001001;
    assign weights1[34][332] = 16'b1111111111100101;
    assign weights1[34][333] = 16'b1111111111011010;
    assign weights1[34][334] = 16'b1111111111011111;
    assign weights1[34][335] = 16'b1111111111100101;
    assign weights1[34][336] = 16'b0000000000000001;
    assign weights1[34][337] = 16'b0000000000010100;
    assign weights1[34][338] = 16'b0000000000001101;
    assign weights1[34][339] = 16'b0000000000000010;
    assign weights1[34][340] = 16'b1111111111101100;
    assign weights1[34][341] = 16'b1111111111101011;
    assign weights1[34][342] = 16'b1111111111110011;
    assign weights1[34][343] = 16'b1111111111100100;
    assign weights1[34][344] = 16'b0000000000000000;
    assign weights1[34][345] = 16'b0000000000000101;
    assign weights1[34][346] = 16'b0000000000001101;
    assign weights1[34][347] = 16'b0000000000010101;
    assign weights1[34][348] = 16'b0000000000011000;
    assign weights1[34][349] = 16'b0000000000101110;
    assign weights1[34][350] = 16'b1111111111110010;
    assign weights1[34][351] = 16'b1111111110101100;
    assign weights1[34][352] = 16'b1111111111001111;
    assign weights1[34][353] = 16'b1111111111111101;
    assign weights1[34][354] = 16'b0000000000010010;
    assign weights1[34][355] = 16'b0000000000100101;
    assign weights1[34][356] = 16'b0000000000010000;
    assign weights1[34][357] = 16'b0000000000010011;
    assign weights1[34][358] = 16'b0000000000001110;
    assign weights1[34][359] = 16'b1111111111111000;
    assign weights1[34][360] = 16'b1111111111100111;
    assign weights1[34][361] = 16'b1111111111100000;
    assign weights1[34][362] = 16'b1111111111101000;
    assign weights1[34][363] = 16'b1111111111110000;
    assign weights1[34][364] = 16'b1111111111111110;
    assign weights1[34][365] = 16'b0000000000010000;
    assign weights1[34][366] = 16'b0000000000000101;
    assign weights1[34][367] = 16'b0000000000001011;
    assign weights1[34][368] = 16'b0000000000000101;
    assign weights1[34][369] = 16'b1111111111101011;
    assign weights1[34][370] = 16'b0000000000010100;
    assign weights1[34][371] = 16'b1111111111110011;
    assign weights1[34][372] = 16'b0000000000000001;
    assign weights1[34][373] = 16'b1111111111110110;
    assign weights1[34][374] = 16'b0000000000001101;
    assign weights1[34][375] = 16'b0000000000001000;
    assign weights1[34][376] = 16'b0000000000011001;
    assign weights1[34][377] = 16'b1111111111111011;
    assign weights1[34][378] = 16'b1111111111100011;
    assign weights1[34][379] = 16'b1111111111011110;
    assign weights1[34][380] = 16'b1111111111011010;
    assign weights1[34][381] = 16'b0000000000001101;
    assign weights1[34][382] = 16'b0000000000010000;
    assign weights1[34][383] = 16'b0000000000100000;
    assign weights1[34][384] = 16'b0000000000011001;
    assign weights1[34][385] = 16'b0000000000001001;
    assign weights1[34][386] = 16'b0000000000000010;
    assign weights1[34][387] = 16'b1111111111100010;
    assign weights1[34][388] = 16'b1111111111110110;
    assign weights1[34][389] = 16'b1111111111011100;
    assign weights1[34][390] = 16'b1111111111101011;
    assign weights1[34][391] = 16'b1111111111110000;
    assign weights1[34][392] = 16'b1111111111111011;
    assign weights1[34][393] = 16'b0000000000000011;
    assign weights1[34][394] = 16'b0000000000001010;
    assign weights1[34][395] = 16'b0000000000001100;
    assign weights1[34][396] = 16'b0000000000001101;
    assign weights1[34][397] = 16'b1111111111110000;
    assign weights1[34][398] = 16'b0000000000001001;
    assign weights1[34][399] = 16'b1111111111110001;
    assign weights1[34][400] = 16'b0000000000000011;
    assign weights1[34][401] = 16'b0000000000010100;
    assign weights1[34][402] = 16'b1111111111111101;
    assign weights1[34][403] = 16'b0000000000010000;
    assign weights1[34][404] = 16'b0000000000001101;
    assign weights1[34][405] = 16'b0000000000000001;
    assign weights1[34][406] = 16'b1111111111101110;
    assign weights1[34][407] = 16'b1111111111011011;
    assign weights1[34][408] = 16'b1111111111111100;
    assign weights1[34][409] = 16'b0000000000010001;
    assign weights1[34][410] = 16'b0000000000001101;
    assign weights1[34][411] = 16'b0000000000010010;
    assign weights1[34][412] = 16'b0000000000000001;
    assign weights1[34][413] = 16'b0000000000010101;
    assign weights1[34][414] = 16'b1111111111111110;
    assign weights1[34][415] = 16'b1111111111110110;
    assign weights1[34][416] = 16'b1111111111110111;
    assign weights1[34][417] = 16'b1111111111110101;
    assign weights1[34][418] = 16'b1111111111100111;
    assign weights1[34][419] = 16'b1111111111110000;
    assign weights1[34][420] = 16'b0000000000001011;
    assign weights1[34][421] = 16'b0000000000001101;
    assign weights1[34][422] = 16'b0000000000011000;
    assign weights1[34][423] = 16'b0000000000001101;
    assign weights1[34][424] = 16'b1111111111111001;
    assign weights1[34][425] = 16'b0000000000000101;
    assign weights1[34][426] = 16'b1111111111110010;
    assign weights1[34][427] = 16'b0000000000000101;
    assign weights1[34][428] = 16'b0000000000000001;
    assign weights1[34][429] = 16'b1111111111111101;
    assign weights1[34][430] = 16'b0000000000001100;
    assign weights1[34][431] = 16'b0000000000000101;
    assign weights1[34][432] = 16'b1111111111111100;
    assign weights1[34][433] = 16'b1111111111111011;
    assign weights1[34][434] = 16'b1111111111101111;
    assign weights1[34][435] = 16'b1111111111101001;
    assign weights1[34][436] = 16'b0000000000000011;
    assign weights1[34][437] = 16'b0000000000010010;
    assign weights1[34][438] = 16'b0000000000001101;
    assign weights1[34][439] = 16'b0000000000011001;
    assign weights1[34][440] = 16'b0000000000001010;
    assign weights1[34][441] = 16'b1111111111111111;
    assign weights1[34][442] = 16'b1111111111111111;
    assign weights1[34][443] = 16'b1111111111111000;
    assign weights1[34][444] = 16'b1111111111100010;
    assign weights1[34][445] = 16'b1111111111111110;
    assign weights1[34][446] = 16'b1111111111111010;
    assign weights1[34][447] = 16'b1111111111110010;
    assign weights1[34][448] = 16'b0000000000000110;
    assign weights1[34][449] = 16'b0000000000001011;
    assign weights1[34][450] = 16'b0000000000001111;
    assign weights1[34][451] = 16'b0000000000000110;
    assign weights1[34][452] = 16'b1111111111111010;
    assign weights1[34][453] = 16'b1111111111111010;
    assign weights1[34][454] = 16'b0000000000000110;
    assign weights1[34][455] = 16'b1111111111111111;
    assign weights1[34][456] = 16'b1111111111100110;
    assign weights1[34][457] = 16'b1111111111111011;
    assign weights1[34][458] = 16'b1111111111111101;
    assign weights1[34][459] = 16'b0000000000000100;
    assign weights1[34][460] = 16'b1111111111110011;
    assign weights1[34][461] = 16'b1111111111111010;
    assign weights1[34][462] = 16'b0000000000000010;
    assign weights1[34][463] = 16'b0000000000000111;
    assign weights1[34][464] = 16'b0000000000000100;
    assign weights1[34][465] = 16'b0000000000001000;
    assign weights1[34][466] = 16'b1111111111111011;
    assign weights1[34][467] = 16'b1111111111110101;
    assign weights1[34][468] = 16'b1111111111111101;
    assign weights1[34][469] = 16'b0000000000000001;
    assign weights1[34][470] = 16'b0000000000000111;
    assign weights1[34][471] = 16'b1111111111100011;
    assign weights1[34][472] = 16'b1111111111110101;
    assign weights1[34][473] = 16'b1111111111111110;
    assign weights1[34][474] = 16'b1111111111111101;
    assign weights1[34][475] = 16'b1111111111111000;
    assign weights1[34][476] = 16'b0000000000000110;
    assign weights1[34][477] = 16'b0000000000000001;
    assign weights1[34][478] = 16'b0000000000010011;
    assign weights1[34][479] = 16'b0000000000000110;
    assign weights1[34][480] = 16'b1111111111110111;
    assign weights1[34][481] = 16'b0000000000000010;
    assign weights1[34][482] = 16'b0000000000001000;
    assign weights1[34][483] = 16'b1111111111111000;
    assign weights1[34][484] = 16'b1111111111100011;
    assign weights1[34][485] = 16'b1111111111110101;
    assign weights1[34][486] = 16'b1111111111111111;
    assign weights1[34][487] = 16'b1111111111100111;
    assign weights1[34][488] = 16'b1111111111111110;
    assign weights1[34][489] = 16'b1111111111110001;
    assign weights1[34][490] = 16'b1111111111101111;
    assign weights1[34][491] = 16'b1111111111111011;
    assign weights1[34][492] = 16'b1111111111111000;
    assign weights1[34][493] = 16'b0000000000010001;
    assign weights1[34][494] = 16'b0000000000000101;
    assign weights1[34][495] = 16'b1111111111111100;
    assign weights1[34][496] = 16'b1111111111111101;
    assign weights1[34][497] = 16'b0000000000001101;
    assign weights1[34][498] = 16'b0000000000000000;
    assign weights1[34][499] = 16'b1111111111111100;
    assign weights1[34][500] = 16'b0000000000001001;
    assign weights1[34][501] = 16'b0000000000001111;
    assign weights1[34][502] = 16'b1111111111111100;
    assign weights1[34][503] = 16'b0000000000000001;
    assign weights1[34][504] = 16'b1111111111110110;
    assign weights1[34][505] = 16'b1111111111111011;
    assign weights1[34][506] = 16'b1111111111111101;
    assign weights1[34][507] = 16'b0000000000000100;
    assign weights1[34][508] = 16'b0000000000001110;
    assign weights1[34][509] = 16'b0000000000000000;
    assign weights1[34][510] = 16'b1111111111110110;
    assign weights1[34][511] = 16'b0000000000001000;
    assign weights1[34][512] = 16'b1111111111110101;
    assign weights1[34][513] = 16'b0000000000001101;
    assign weights1[34][514] = 16'b1111111111111111;
    assign weights1[34][515] = 16'b0000000000000010;
    assign weights1[34][516] = 16'b1111111111111111;
    assign weights1[34][517] = 16'b0000000000000110;
    assign weights1[34][518] = 16'b1111111111110111;
    assign weights1[34][519] = 16'b0000000000001101;
    assign weights1[34][520] = 16'b0000000000010000;
    assign weights1[34][521] = 16'b1111111111110110;
    assign weights1[34][522] = 16'b1111111111111110;
    assign weights1[34][523] = 16'b1111111111110111;
    assign weights1[34][524] = 16'b1111111111101100;
    assign weights1[34][525] = 16'b0000000000000101;
    assign weights1[34][526] = 16'b1111111111111010;
    assign weights1[34][527] = 16'b0000000000001000;
    assign weights1[34][528] = 16'b1111111111111101;
    assign weights1[34][529] = 16'b0000000000010010;
    assign weights1[34][530] = 16'b1111111111111110;
    assign weights1[34][531] = 16'b0000000000000110;
    assign weights1[34][532] = 16'b1111111111111110;
    assign weights1[34][533] = 16'b1111111111111100;
    assign weights1[34][534] = 16'b1111111111110110;
    assign weights1[34][535] = 16'b1111111111101111;
    assign weights1[34][536] = 16'b0000000000000001;
    assign weights1[34][537] = 16'b0000000000010111;
    assign weights1[34][538] = 16'b1111111111111010;
    assign weights1[34][539] = 16'b1111111111101011;
    assign weights1[34][540] = 16'b1111111111111011;
    assign weights1[34][541] = 16'b1111111111110111;
    assign weights1[34][542] = 16'b1111111111101101;
    assign weights1[34][543] = 16'b1111111111110111;
    assign weights1[34][544] = 16'b1111111111101000;
    assign weights1[34][545] = 16'b1111111111110001;
    assign weights1[34][546] = 16'b0000000000000001;
    assign weights1[34][547] = 16'b0000000000000001;
    assign weights1[34][548] = 16'b1111111111101110;
    assign weights1[34][549] = 16'b1111111111110110;
    assign weights1[34][550] = 16'b1111111111111111;
    assign weights1[34][551] = 16'b1111111111111011;
    assign weights1[34][552] = 16'b0000000000000001;
    assign weights1[34][553] = 16'b1111111111110010;
    assign weights1[34][554] = 16'b0000000000010100;
    assign weights1[34][555] = 16'b1111111111111101;
    assign weights1[34][556] = 16'b1111111111111101;
    assign weights1[34][557] = 16'b0000000000000011;
    assign weights1[34][558] = 16'b0000000000001010;
    assign weights1[34][559] = 16'b0000000000000110;
    assign weights1[34][560] = 16'b1111111111111011;
    assign weights1[34][561] = 16'b1111111111111001;
    assign weights1[34][562] = 16'b1111111111101011;
    assign weights1[34][563] = 16'b1111111111110101;
    assign weights1[34][564] = 16'b1111111111111101;
    assign weights1[34][565] = 16'b1111111111110100;
    assign weights1[34][566] = 16'b1111111111111010;
    assign weights1[34][567] = 16'b1111111111111110;
    assign weights1[34][568] = 16'b1111111111110100;
    assign weights1[34][569] = 16'b1111111111110110;
    assign weights1[34][570] = 16'b0000000000010011;
    assign weights1[34][571] = 16'b0000000000000110;
    assign weights1[34][572] = 16'b1111111111111111;
    assign weights1[34][573] = 16'b0000000000000000;
    assign weights1[34][574] = 16'b0000000000000001;
    assign weights1[34][575] = 16'b0000000000000111;
    assign weights1[34][576] = 16'b0000000000010001;
    assign weights1[34][577] = 16'b0000000000001011;
    assign weights1[34][578] = 16'b1111111111111000;
    assign weights1[34][579] = 16'b1111111111111000;
    assign weights1[34][580] = 16'b1111111111110001;
    assign weights1[34][581] = 16'b0000000000001001;
    assign weights1[34][582] = 16'b0000000000001100;
    assign weights1[34][583] = 16'b0000000000001100;
    assign weights1[34][584] = 16'b0000000000001100;
    assign weights1[34][585] = 16'b0000000000000100;
    assign weights1[34][586] = 16'b0000000000000011;
    assign weights1[34][587] = 16'b0000000000000101;
    assign weights1[34][588] = 16'b1111111111111010;
    assign weights1[34][589] = 16'b1111111111111010;
    assign weights1[34][590] = 16'b1111111111101110;
    assign weights1[34][591] = 16'b1111111111100110;
    assign weights1[34][592] = 16'b1111111111111111;
    assign weights1[34][593] = 16'b1111111111111001;
    assign weights1[34][594] = 16'b1111111111100101;
    assign weights1[34][595] = 16'b0000000000000001;
    assign weights1[34][596] = 16'b1111111111101101;
    assign weights1[34][597] = 16'b0000000000010000;
    assign weights1[34][598] = 16'b0000000000000010;
    assign weights1[34][599] = 16'b1111111111111100;
    assign weights1[34][600] = 16'b1111111111111010;
    assign weights1[34][601] = 16'b0000000000000000;
    assign weights1[34][602] = 16'b1111111111101101;
    assign weights1[34][603] = 16'b1111111111111111;
    assign weights1[34][604] = 16'b1111111111110101;
    assign weights1[34][605] = 16'b0000000000000100;
    assign weights1[34][606] = 16'b0000000000000010;
    assign weights1[34][607] = 16'b0000000000010100;
    assign weights1[34][608] = 16'b0000000000000000;
    assign weights1[34][609] = 16'b0000000000000000;
    assign weights1[34][610] = 16'b1111111111111011;
    assign weights1[34][611] = 16'b1111111111111110;
    assign weights1[34][612] = 16'b1111111111111100;
    assign weights1[34][613] = 16'b1111111111111100;
    assign weights1[34][614] = 16'b0000000000000011;
    assign weights1[34][615] = 16'b0000000000000100;
    assign weights1[34][616] = 16'b0000000000000010;
    assign weights1[34][617] = 16'b1111111111111000;
    assign weights1[34][618] = 16'b1111111111111110;
    assign weights1[34][619] = 16'b1111111111110000;
    assign weights1[34][620] = 16'b0000000000000000;
    assign weights1[34][621] = 16'b1111111111110010;
    assign weights1[34][622] = 16'b0000000000000000;
    assign weights1[34][623] = 16'b0000000000000101;
    assign weights1[34][624] = 16'b1111111111111100;
    assign weights1[34][625] = 16'b0000000000001111;
    assign weights1[34][626] = 16'b1111111111111110;
    assign weights1[34][627] = 16'b0000000000000100;
    assign weights1[34][628] = 16'b0000000000000000;
    assign weights1[34][629] = 16'b0000000000000111;
    assign weights1[34][630] = 16'b1111111111110100;
    assign weights1[34][631] = 16'b1111111111111110;
    assign weights1[34][632] = 16'b1111111111110100;
    assign weights1[34][633] = 16'b1111111111110110;
    assign weights1[34][634] = 16'b0000000000000011;
    assign weights1[34][635] = 16'b1111111111100001;
    assign weights1[34][636] = 16'b0000000000100100;
    assign weights1[34][637] = 16'b0000000000001010;
    assign weights1[34][638] = 16'b0000000000001011;
    assign weights1[34][639] = 16'b0000000000000011;
    assign weights1[34][640] = 16'b1111111111110000;
    assign weights1[34][641] = 16'b1111111111110111;
    assign weights1[34][642] = 16'b0000000000000110;
    assign weights1[34][643] = 16'b0000000000000000;
    assign weights1[34][644] = 16'b1111111111111011;
    assign weights1[34][645] = 16'b1111111111111011;
    assign weights1[34][646] = 16'b0000000000001110;
    assign weights1[34][647] = 16'b1111111111111001;
    assign weights1[34][648] = 16'b0000000000000010;
    assign weights1[34][649] = 16'b0000000000000100;
    assign weights1[34][650] = 16'b0000000000001000;
    assign weights1[34][651] = 16'b0000000000001111;
    assign weights1[34][652] = 16'b1111111111110100;
    assign weights1[34][653] = 16'b0000000000010001;
    assign weights1[34][654] = 16'b1111111111111101;
    assign weights1[34][655] = 16'b1111111111111100;
    assign weights1[34][656] = 16'b1111111111111000;
    assign weights1[34][657] = 16'b1111111111101001;
    assign weights1[34][658] = 16'b0000000000000010;
    assign weights1[34][659] = 16'b1111111111110000;
    assign weights1[34][660] = 16'b1111111111111101;
    assign weights1[34][661] = 16'b0000000000000100;
    assign weights1[34][662] = 16'b1111111111101010;
    assign weights1[34][663] = 16'b0000000000001001;
    assign weights1[34][664] = 16'b0000000000000101;
    assign weights1[34][665] = 16'b1111111111111111;
    assign weights1[34][666] = 16'b0000000000000000;
    assign weights1[34][667] = 16'b0000000000000100;
    assign weights1[34][668] = 16'b0000000000010001;
    assign weights1[34][669] = 16'b0000000000010000;
    assign weights1[34][670] = 16'b0000000000000100;
    assign weights1[34][671] = 16'b0000000000000001;
    assign weights1[34][672] = 16'b0000000000000101;
    assign weights1[34][673] = 16'b1111111111111101;
    assign weights1[34][674] = 16'b0000000000001000;
    assign weights1[34][675] = 16'b0000000000000110;
    assign weights1[34][676] = 16'b1111111111111101;
    assign weights1[34][677] = 16'b0000000000000101;
    assign weights1[34][678] = 16'b1111111111111100;
    assign weights1[34][679] = 16'b0000000000010010;
    assign weights1[34][680] = 16'b1111111111111000;
    assign weights1[34][681] = 16'b1111111111110001;
    assign weights1[34][682] = 16'b1111111111111011;
    assign weights1[34][683] = 16'b1111111111111010;
    assign weights1[34][684] = 16'b0000000000000010;
    assign weights1[34][685] = 16'b0000000000010000;
    assign weights1[34][686] = 16'b0000000000000110;
    assign weights1[34][687] = 16'b1111111111111010;
    assign weights1[34][688] = 16'b1111111111111111;
    assign weights1[34][689] = 16'b0000000000000000;
    assign weights1[34][690] = 16'b1111111111100111;
    assign weights1[34][691] = 16'b1111111111111001;
    assign weights1[34][692] = 16'b1111111111110111;
    assign weights1[34][693] = 16'b1111111111110110;
    assign weights1[34][694] = 16'b0000000000000011;
    assign weights1[34][695] = 16'b0000000000000000;
    assign weights1[34][696] = 16'b1111111111111110;
    assign weights1[34][697] = 16'b0000000000001101;
    assign weights1[34][698] = 16'b0000000000001101;
    assign weights1[34][699] = 16'b0000000000000110;
    assign weights1[34][700] = 16'b0000000000000110;
    assign weights1[34][701] = 16'b0000000000000000;
    assign weights1[34][702] = 16'b1111111111111100;
    assign weights1[34][703] = 16'b1111111111111011;
    assign weights1[34][704] = 16'b0000000000000100;
    assign weights1[34][705] = 16'b1111111111111100;
    assign weights1[34][706] = 16'b0000000000000111;
    assign weights1[34][707] = 16'b1111111111111111;
    assign weights1[34][708] = 16'b0000000000000100;
    assign weights1[34][709] = 16'b0000000000001100;
    assign weights1[34][710] = 16'b0000000000001000;
    assign weights1[34][711] = 16'b0000000000000101;
    assign weights1[34][712] = 16'b0000000000000011;
    assign weights1[34][713] = 16'b0000000000000010;
    assign weights1[34][714] = 16'b1111111111101110;
    assign weights1[34][715] = 16'b0000000000001011;
    assign weights1[34][716] = 16'b1111111111110101;
    assign weights1[34][717] = 16'b1111111111111000;
    assign weights1[34][718] = 16'b0000000000000100;
    assign weights1[34][719] = 16'b0000000000000001;
    assign weights1[34][720] = 16'b1111111111101011;
    assign weights1[34][721] = 16'b1111111111101111;
    assign weights1[34][722] = 16'b1111111111110101;
    assign weights1[34][723] = 16'b0000000000000010;
    assign weights1[34][724] = 16'b1111111111110011;
    assign weights1[34][725] = 16'b0000000000000011;
    assign weights1[34][726] = 16'b0000000000001000;
    assign weights1[34][727] = 16'b0000000000000110;
    assign weights1[34][728] = 16'b0000000000000100;
    assign weights1[34][729] = 16'b0000000000000010;
    assign weights1[34][730] = 16'b0000000000000001;
    assign weights1[34][731] = 16'b0000000000000100;
    assign weights1[34][732] = 16'b0000000000000000;
    assign weights1[34][733] = 16'b0000000000001000;
    assign weights1[34][734] = 16'b0000000000001001;
    assign weights1[34][735] = 16'b0000000000001100;
    assign weights1[34][736] = 16'b0000000000000010;
    assign weights1[34][737] = 16'b0000000000001011;
    assign weights1[34][738] = 16'b1111111111111110;
    assign weights1[34][739] = 16'b1111111111110111;
    assign weights1[34][740] = 16'b1111111111111011;
    assign weights1[34][741] = 16'b1111111111110101;
    assign weights1[34][742] = 16'b1111111111110100;
    assign weights1[34][743] = 16'b1111111111111001;
    assign weights1[34][744] = 16'b1111111111111011;
    assign weights1[34][745] = 16'b1111111111111000;
    assign weights1[34][746] = 16'b0000000000001001;
    assign weights1[34][747] = 16'b0000000000000110;
    assign weights1[34][748] = 16'b0000000000011011;
    assign weights1[34][749] = 16'b0000000000011011;
    assign weights1[34][750] = 16'b0000000000010100;
    assign weights1[34][751] = 16'b0000000000000010;
    assign weights1[34][752] = 16'b1111111111110100;
    assign weights1[34][753] = 16'b1111111111111101;
    assign weights1[34][754] = 16'b1111111111111100;
    assign weights1[34][755] = 16'b0000000000000001;
    assign weights1[34][756] = 16'b0000000000000001;
    assign weights1[34][757] = 16'b0000000000000011;
    assign weights1[34][758] = 16'b1111111111111011;
    assign weights1[34][759] = 16'b0000000000000000;
    assign weights1[34][760] = 16'b1111111111101010;
    assign weights1[34][761] = 16'b1111111111111001;
    assign weights1[34][762] = 16'b0000000000010010;
    assign weights1[34][763] = 16'b0000000000001011;
    assign weights1[34][764] = 16'b1111111111111111;
    assign weights1[34][765] = 16'b0000000000000100;
    assign weights1[34][766] = 16'b0000000000000110;
    assign weights1[34][767] = 16'b0000000000001001;
    assign weights1[34][768] = 16'b0000000000000011;
    assign weights1[34][769] = 16'b0000000000001000;
    assign weights1[34][770] = 16'b0000000000000101;
    assign weights1[34][771] = 16'b0000000000001010;
    assign weights1[34][772] = 16'b0000000000001010;
    assign weights1[34][773] = 16'b0000000000001100;
    assign weights1[34][774] = 16'b0000000000000110;
    assign weights1[34][775] = 16'b0000000000001101;
    assign weights1[34][776] = 16'b0000000000010001;
    assign weights1[34][777] = 16'b0000000000001110;
    assign weights1[34][778] = 16'b0000000000010001;
    assign weights1[34][779] = 16'b0000000000000101;
    assign weights1[34][780] = 16'b1111111111111011;
    assign weights1[34][781] = 16'b1111111111111101;
    assign weights1[34][782] = 16'b1111111111111101;
    assign weights1[34][783] = 16'b0000000000000010;
    assign weights1[35][0] = 16'b0000000000000001;
    assign weights1[35][1] = 16'b0000000000000001;
    assign weights1[35][2] = 16'b0000000000000011;
    assign weights1[35][3] = 16'b0000000000001110;
    assign weights1[35][4] = 16'b0000000000010111;
    assign weights1[35][5] = 16'b0000000000010011;
    assign weights1[35][6] = 16'b0000000000100001;
    assign weights1[35][7] = 16'b0000000000011000;
    assign weights1[35][8] = 16'b0000000000011010;
    assign weights1[35][9] = 16'b0000000000100011;
    assign weights1[35][10] = 16'b0000000000011101;
    assign weights1[35][11] = 16'b0000000000000011;
    assign weights1[35][12] = 16'b0000000000100111;
    assign weights1[35][13] = 16'b0000000000011000;
    assign weights1[35][14] = 16'b0000000000010100;
    assign weights1[35][15] = 16'b0000000000000110;
    assign weights1[35][16] = 16'b0000000000001111;
    assign weights1[35][17] = 16'b0000000000010010;
    assign weights1[35][18] = 16'b0000000000010111;
    assign weights1[35][19] = 16'b0000000000001111;
    assign weights1[35][20] = 16'b0000000000000011;
    assign weights1[35][21] = 16'b0000000000001001;
    assign weights1[35][22] = 16'b0000000000001111;
    assign weights1[35][23] = 16'b0000000000001010;
    assign weights1[35][24] = 16'b0000000000000001;
    assign weights1[35][25] = 16'b0000000000000011;
    assign weights1[35][26] = 16'b1111111111111101;
    assign weights1[35][27] = 16'b1111111111111111;
    assign weights1[35][28] = 16'b0000000000000000;
    assign weights1[35][29] = 16'b0000000000000011;
    assign weights1[35][30] = 16'b0000000000010001;
    assign weights1[35][31] = 16'b0000000000011000;
    assign weights1[35][32] = 16'b0000000000011011;
    assign weights1[35][33] = 16'b0000000000010000;
    assign weights1[35][34] = 16'b0000000000011010;
    assign weights1[35][35] = 16'b0000000000010000;
    assign weights1[35][36] = 16'b1111111111111001;
    assign weights1[35][37] = 16'b0000000000001011;
    assign weights1[35][38] = 16'b1111111111111111;
    assign weights1[35][39] = 16'b1111111111101110;
    assign weights1[35][40] = 16'b0000000000000110;
    assign weights1[35][41] = 16'b0000000000001011;
    assign weights1[35][42] = 16'b1111111111111010;
    assign weights1[35][43] = 16'b0000000000001000;
    assign weights1[35][44] = 16'b0000000000001101;
    assign weights1[35][45] = 16'b0000000000000000;
    assign weights1[35][46] = 16'b1111111111111111;
    assign weights1[35][47] = 16'b0000000000001100;
    assign weights1[35][48] = 16'b1111111111110111;
    assign weights1[35][49] = 16'b0000000000001111;
    assign weights1[35][50] = 16'b0000000000001011;
    assign weights1[35][51] = 16'b1111111111111111;
    assign weights1[35][52] = 16'b1111111111111000;
    assign weights1[35][53] = 16'b0000000000001001;
    assign weights1[35][54] = 16'b0000000000000111;
    assign weights1[35][55] = 16'b0000000000000100;
    assign weights1[35][56] = 16'b1111111111111101;
    assign weights1[35][57] = 16'b0000000000001001;
    assign weights1[35][58] = 16'b0000000000001111;
    assign weights1[35][59] = 16'b0000000000001010;
    assign weights1[35][60] = 16'b0000000000001000;
    assign weights1[35][61] = 16'b0000000000010011;
    assign weights1[35][62] = 16'b0000000000011010;
    assign weights1[35][63] = 16'b0000000000000101;
    assign weights1[35][64] = 16'b1111111111111100;
    assign weights1[35][65] = 16'b0000000000001110;
    assign weights1[35][66] = 16'b0000000000000100;
    assign weights1[35][67] = 16'b1111111111111011;
    assign weights1[35][68] = 16'b1111111111110011;
    assign weights1[35][69] = 16'b0000000000000111;
    assign weights1[35][70] = 16'b1111111111111010;
    assign weights1[35][71] = 16'b1111111111110110;
    assign weights1[35][72] = 16'b1111111111111001;
    assign weights1[35][73] = 16'b1111111111101110;
    assign weights1[35][74] = 16'b0000000000010001;
    assign weights1[35][75] = 16'b0000000000000001;
    assign weights1[35][76] = 16'b0000000000000100;
    assign weights1[35][77] = 16'b0000000000001110;
    assign weights1[35][78] = 16'b1111111111111101;
    assign weights1[35][79] = 16'b1111111111101101;
    assign weights1[35][80] = 16'b0000000000000011;
    assign weights1[35][81] = 16'b1111111111111000;
    assign weights1[35][82] = 16'b1111111111111001;
    assign weights1[35][83] = 16'b0000000000001000;
    assign weights1[35][84] = 16'b1111111111111011;
    assign weights1[35][85] = 16'b0000000000000111;
    assign weights1[35][86] = 16'b0000000000000011;
    assign weights1[35][87] = 16'b0000000000000011;
    assign weights1[35][88] = 16'b0000000000011101;
    assign weights1[35][89] = 16'b0000000000000111;
    assign weights1[35][90] = 16'b0000000000000110;
    assign weights1[35][91] = 16'b0000000000001110;
    assign weights1[35][92] = 16'b1111111111110101;
    assign weights1[35][93] = 16'b1111111111111011;
    assign weights1[35][94] = 16'b1111111111111001;
    assign weights1[35][95] = 16'b1111111111101010;
    assign weights1[35][96] = 16'b1111111111110100;
    assign weights1[35][97] = 16'b1111111111101110;
    assign weights1[35][98] = 16'b1111111111111000;
    assign weights1[35][99] = 16'b1111111111110011;
    assign weights1[35][100] = 16'b1111111111111111;
    assign weights1[35][101] = 16'b0000000000000001;
    assign weights1[35][102] = 16'b1111111111110100;
    assign weights1[35][103] = 16'b0000000000000100;
    assign weights1[35][104] = 16'b1111111111111010;
    assign weights1[35][105] = 16'b1111111111111000;
    assign weights1[35][106] = 16'b1111111111111111;
    assign weights1[35][107] = 16'b0000000000000110;
    assign weights1[35][108] = 16'b1111111111111010;
    assign weights1[35][109] = 16'b0000000000001000;
    assign weights1[35][110] = 16'b1111111111111110;
    assign weights1[35][111] = 16'b1111111111111110;
    assign weights1[35][112] = 16'b1111111111111011;
    assign weights1[35][113] = 16'b0000000000000000;
    assign weights1[35][114] = 16'b1111111111111010;
    assign weights1[35][115] = 16'b1111111111111011;
    assign weights1[35][116] = 16'b0000000000000100;
    assign weights1[35][117] = 16'b0000000000000110;
    assign weights1[35][118] = 16'b1111111111111101;
    assign weights1[35][119] = 16'b1111111111110001;
    assign weights1[35][120] = 16'b1111111111110111;
    assign weights1[35][121] = 16'b0000000000001000;
    assign weights1[35][122] = 16'b1111111111110011;
    assign weights1[35][123] = 16'b1111111111110111;
    assign weights1[35][124] = 16'b1111111111111111;
    assign weights1[35][125] = 16'b1111111111111001;
    assign weights1[35][126] = 16'b1111111111110110;
    assign weights1[35][127] = 16'b1111111111110110;
    assign weights1[35][128] = 16'b1111111111110100;
    assign weights1[35][129] = 16'b0000000000000001;
    assign weights1[35][130] = 16'b1111111111111110;
    assign weights1[35][131] = 16'b1111111111110010;
    assign weights1[35][132] = 16'b1111111111111001;
    assign weights1[35][133] = 16'b1111111111111111;
    assign weights1[35][134] = 16'b1111111111101111;
    assign weights1[35][135] = 16'b1111111111111010;
    assign weights1[35][136] = 16'b1111111111111000;
    assign weights1[35][137] = 16'b0000000000000100;
    assign weights1[35][138] = 16'b0000000000000110;
    assign weights1[35][139] = 16'b1111111111110100;
    assign weights1[35][140] = 16'b1111111111110111;
    assign weights1[35][141] = 16'b1111111111111100;
    assign weights1[35][142] = 16'b1111111111111011;
    assign weights1[35][143] = 16'b1111111111110110;
    assign weights1[35][144] = 16'b1111111111111110;
    assign weights1[35][145] = 16'b1111111111111111;
    assign weights1[35][146] = 16'b0000000000001100;
    assign weights1[35][147] = 16'b1111111111110011;
    assign weights1[35][148] = 16'b1111111111110110;
    assign weights1[35][149] = 16'b1111111111111101;
    assign weights1[35][150] = 16'b1111111111111111;
    assign weights1[35][151] = 16'b1111111111110111;
    assign weights1[35][152] = 16'b1111111111111100;
    assign weights1[35][153] = 16'b1111111111110111;
    assign weights1[35][154] = 16'b1111111111110001;
    assign weights1[35][155] = 16'b1111111111111000;
    assign weights1[35][156] = 16'b1111111111110010;
    assign weights1[35][157] = 16'b1111111111110001;
    assign weights1[35][158] = 16'b1111111111100100;
    assign weights1[35][159] = 16'b1111111111110111;
    assign weights1[35][160] = 16'b1111111111111100;
    assign weights1[35][161] = 16'b1111111111100100;
    assign weights1[35][162] = 16'b1111111111111001;
    assign weights1[35][163] = 16'b1111111111111111;
    assign weights1[35][164] = 16'b0000000000000101;
    assign weights1[35][165] = 16'b0000000000001010;
    assign weights1[35][166] = 16'b1111111111111010;
    assign weights1[35][167] = 16'b1111111111111000;
    assign weights1[35][168] = 16'b1111111111111000;
    assign weights1[35][169] = 16'b0000000000000100;
    assign weights1[35][170] = 16'b1111111111111001;
    assign weights1[35][171] = 16'b1111111111110001;
    assign weights1[35][172] = 16'b0000000000001001;
    assign weights1[35][173] = 16'b1111111111110111;
    assign weights1[35][174] = 16'b1111111111110110;
    assign weights1[35][175] = 16'b1111111111111110;
    assign weights1[35][176] = 16'b0000000000000001;
    assign weights1[35][177] = 16'b1111111111111011;
    assign weights1[35][178] = 16'b1111111111111111;
    assign weights1[35][179] = 16'b1111111111110000;
    assign weights1[35][180] = 16'b1111111111111111;
    assign weights1[35][181] = 16'b1111111111111110;
    assign weights1[35][182] = 16'b1111111111111111;
    assign weights1[35][183] = 16'b1111111111111100;
    assign weights1[35][184] = 16'b1111111111110011;
    assign weights1[35][185] = 16'b1111111111111011;
    assign weights1[35][186] = 16'b0000000000000101;
    assign weights1[35][187] = 16'b1111111111101101;
    assign weights1[35][188] = 16'b1111111111110110;
    assign weights1[35][189] = 16'b0000000000000110;
    assign weights1[35][190] = 16'b0000000000001000;
    assign weights1[35][191] = 16'b1111111111111111;
    assign weights1[35][192] = 16'b1111111111100101;
    assign weights1[35][193] = 16'b1111111111110010;
    assign weights1[35][194] = 16'b1111111111111101;
    assign weights1[35][195] = 16'b1111111111110111;
    assign weights1[35][196] = 16'b1111111111111101;
    assign weights1[35][197] = 16'b0000000000000101;
    assign weights1[35][198] = 16'b1111111111111100;
    assign weights1[35][199] = 16'b0000000000000000;
    assign weights1[35][200] = 16'b0000000000000011;
    assign weights1[35][201] = 16'b0000000000000101;
    assign weights1[35][202] = 16'b0000000000000100;
    assign weights1[35][203] = 16'b0000000000000011;
    assign weights1[35][204] = 16'b1111111111111011;
    assign weights1[35][205] = 16'b0000000000000010;
    assign weights1[35][206] = 16'b1111111111110110;
    assign weights1[35][207] = 16'b0000000000000010;
    assign weights1[35][208] = 16'b1111111111111010;
    assign weights1[35][209] = 16'b1111111111110110;
    assign weights1[35][210] = 16'b0000000000001010;
    assign weights1[35][211] = 16'b1111111111111111;
    assign weights1[35][212] = 16'b0000000000000010;
    assign weights1[35][213] = 16'b1111111111111111;
    assign weights1[35][214] = 16'b0000000000000011;
    assign weights1[35][215] = 16'b0000000000000101;
    assign weights1[35][216] = 16'b0000000000001110;
    assign weights1[35][217] = 16'b1111111111110101;
    assign weights1[35][218] = 16'b1111111111110000;
    assign weights1[35][219] = 16'b1111111111111010;
    assign weights1[35][220] = 16'b1111111111111010;
    assign weights1[35][221] = 16'b0000000000000001;
    assign weights1[35][222] = 16'b1111111111111011;
    assign weights1[35][223] = 16'b1111111111101100;
    assign weights1[35][224] = 16'b1111111111110010;
    assign weights1[35][225] = 16'b0000000000000000;
    assign weights1[35][226] = 16'b1111111111110101;
    assign weights1[35][227] = 16'b1111111111110101;
    assign weights1[35][228] = 16'b0000000000000100;
    assign weights1[35][229] = 16'b1111111111111000;
    assign weights1[35][230] = 16'b1111111111110101;
    assign weights1[35][231] = 16'b1111111111111001;
    assign weights1[35][232] = 16'b1111111111111001;
    assign weights1[35][233] = 16'b0000000000001101;
    assign weights1[35][234] = 16'b1111111111111000;
    assign weights1[35][235] = 16'b0000000000001010;
    assign weights1[35][236] = 16'b0000000000000001;
    assign weights1[35][237] = 16'b0000000000000011;
    assign weights1[35][238] = 16'b0000000000000000;
    assign weights1[35][239] = 16'b0000000000000111;
    assign weights1[35][240] = 16'b1111111111111110;
    assign weights1[35][241] = 16'b0000000000000010;
    assign weights1[35][242] = 16'b0000000000001001;
    assign weights1[35][243] = 16'b1111111111111101;
    assign weights1[35][244] = 16'b1111111111110010;
    assign weights1[35][245] = 16'b1111111111110001;
    assign weights1[35][246] = 16'b1111111111101101;
    assign weights1[35][247] = 16'b0000000000000100;
    assign weights1[35][248] = 16'b0000000000000001;
    assign weights1[35][249] = 16'b0000000000001111;
    assign weights1[35][250] = 16'b1111111111110011;
    assign weights1[35][251] = 16'b1111111111110111;
    assign weights1[35][252] = 16'b1111111111111001;
    assign weights1[35][253] = 16'b1111111111110100;
    assign weights1[35][254] = 16'b0000000000000000;
    assign weights1[35][255] = 16'b1111111111110110;
    assign weights1[35][256] = 16'b1111111111111111;
    assign weights1[35][257] = 16'b0000000000001000;
    assign weights1[35][258] = 16'b1111111111101100;
    assign weights1[35][259] = 16'b1111111111111101;
    assign weights1[35][260] = 16'b1111111111111111;
    assign weights1[35][261] = 16'b0000000000001001;
    assign weights1[35][262] = 16'b0000000000010000;
    assign weights1[35][263] = 16'b1111111111111010;
    assign weights1[35][264] = 16'b0000000000010000;
    assign weights1[35][265] = 16'b0000000000001001;
    assign weights1[35][266] = 16'b0000000000001111;
    assign weights1[35][267] = 16'b0000000000001000;
    assign weights1[35][268] = 16'b1111111111111111;
    assign weights1[35][269] = 16'b1111111111110001;
    assign weights1[35][270] = 16'b0000000000000101;
    assign weights1[35][271] = 16'b0000000000000011;
    assign weights1[35][272] = 16'b0000000000001100;
    assign weights1[35][273] = 16'b1111111111111101;
    assign weights1[35][274] = 16'b0000000000010010;
    assign weights1[35][275] = 16'b1111111111111011;
    assign weights1[35][276] = 16'b0000000000001001;
    assign weights1[35][277] = 16'b0000000000000000;
    assign weights1[35][278] = 16'b1111111111101011;
    assign weights1[35][279] = 16'b0000000000000001;
    assign weights1[35][280] = 16'b1111111111111011;
    assign weights1[35][281] = 16'b0000000000000000;
    assign weights1[35][282] = 16'b0000000000001000;
    assign weights1[35][283] = 16'b1111111111111001;
    assign weights1[35][284] = 16'b1111111111111101;
    assign weights1[35][285] = 16'b1111111111111110;
    assign weights1[35][286] = 16'b0000000000000011;
    assign weights1[35][287] = 16'b0000000000001100;
    assign weights1[35][288] = 16'b0000000000000010;
    assign weights1[35][289] = 16'b0000000000000011;
    assign weights1[35][290] = 16'b0000000000010011;
    assign weights1[35][291] = 16'b0000000000001011;
    assign weights1[35][292] = 16'b0000000000001010;
    assign weights1[35][293] = 16'b1111111111111100;
    assign weights1[35][294] = 16'b1111111111111100;
    assign weights1[35][295] = 16'b1111111111111110;
    assign weights1[35][296] = 16'b0000000000000110;
    assign weights1[35][297] = 16'b0000000000001000;
    assign weights1[35][298] = 16'b1111111111111110;
    assign weights1[35][299] = 16'b0000000000001010;
    assign weights1[35][300] = 16'b1111111111111101;
    assign weights1[35][301] = 16'b0000000000000001;
    assign weights1[35][302] = 16'b0000000000010000;
    assign weights1[35][303] = 16'b0000000000001001;
    assign weights1[35][304] = 16'b1111111111101111;
    assign weights1[35][305] = 16'b0000000000001101;
    assign weights1[35][306] = 16'b0000000000000010;
    assign weights1[35][307] = 16'b0000000000001101;
    assign weights1[35][308] = 16'b1111111111111101;
    assign weights1[35][309] = 16'b0000000000001001;
    assign weights1[35][310] = 16'b0000000000001111;
    assign weights1[35][311] = 16'b0000000000011110;
    assign weights1[35][312] = 16'b0000000000001001;
    assign weights1[35][313] = 16'b1111111111111000;
    assign weights1[35][314] = 16'b1111111111111101;
    assign weights1[35][315] = 16'b1111111111111110;
    assign weights1[35][316] = 16'b0000000000001011;
    assign weights1[35][317] = 16'b0000000000001011;
    assign weights1[35][318] = 16'b0000000000001001;
    assign weights1[35][319] = 16'b1111111111111011;
    assign weights1[35][320] = 16'b0000000000000001;
    assign weights1[35][321] = 16'b1111111111111001;
    assign weights1[35][322] = 16'b0000000000001100;
    assign weights1[35][323] = 16'b0000000000000010;
    assign weights1[35][324] = 16'b0000000000000001;
    assign weights1[35][325] = 16'b0000000000000101;
    assign weights1[35][326] = 16'b0000000000001011;
    assign weights1[35][327] = 16'b0000000000001000;
    assign weights1[35][328] = 16'b0000000000000111;
    assign weights1[35][329] = 16'b0000000000011010;
    assign weights1[35][330] = 16'b0000000000000000;
    assign weights1[35][331] = 16'b0000000000011000;
    assign weights1[35][332] = 16'b0000000000001100;
    assign weights1[35][333] = 16'b0000000000010010;
    assign weights1[35][334] = 16'b0000000000000010;
    assign weights1[35][335] = 16'b0000000000001001;
    assign weights1[35][336] = 16'b0000000000000111;
    assign weights1[35][337] = 16'b0000000000001111;
    assign weights1[35][338] = 16'b0000000000011111;
    assign weights1[35][339] = 16'b1111111111111110;
    assign weights1[35][340] = 16'b0000000000000100;
    assign weights1[35][341] = 16'b0000000000010100;
    assign weights1[35][342] = 16'b0000000000001011;
    assign weights1[35][343] = 16'b0000000000000010;
    assign weights1[35][344] = 16'b1111111111110000;
    assign weights1[35][345] = 16'b0000000000000100;
    assign weights1[35][346] = 16'b1111111111111011;
    assign weights1[35][347] = 16'b0000000000010101;
    assign weights1[35][348] = 16'b0000000000011000;
    assign weights1[35][349] = 16'b0000000000000110;
    assign weights1[35][350] = 16'b0000000000000010;
    assign weights1[35][351] = 16'b0000000000001011;
    assign weights1[35][352] = 16'b1111111111111110;
    assign weights1[35][353] = 16'b0000000000000101;
    assign weights1[35][354] = 16'b0000000000000010;
    assign weights1[35][355] = 16'b1111111111111111;
    assign weights1[35][356] = 16'b0000000000000111;
    assign weights1[35][357] = 16'b0000000000000010;
    assign weights1[35][358] = 16'b0000000000001000;
    assign weights1[35][359] = 16'b0000000000011010;
    assign weights1[35][360] = 16'b1111111111111111;
    assign weights1[35][361] = 16'b0000000000001001;
    assign weights1[35][362] = 16'b0000000000010000;
    assign weights1[35][363] = 16'b0000000000010101;
    assign weights1[35][364] = 16'b0000000000001101;
    assign weights1[35][365] = 16'b0000000000001110;
    assign weights1[35][366] = 16'b0000000000010000;
    assign weights1[35][367] = 16'b0000000000010010;
    assign weights1[35][368] = 16'b0000000000000111;
    assign weights1[35][369] = 16'b0000000000001100;
    assign weights1[35][370] = 16'b1111111111111001;
    assign weights1[35][371] = 16'b0000000000000001;
    assign weights1[35][372] = 16'b0000000000011010;
    assign weights1[35][373] = 16'b1111111111111100;
    assign weights1[35][374] = 16'b0000000000000101;
    assign weights1[35][375] = 16'b1111111111111101;
    assign weights1[35][376] = 16'b0000000000000010;
    assign weights1[35][377] = 16'b0000000000000111;
    assign weights1[35][378] = 16'b0000000000001000;
    assign weights1[35][379] = 16'b0000000000001000;
    assign weights1[35][380] = 16'b0000000000000101;
    assign weights1[35][381] = 16'b0000000000001101;
    assign weights1[35][382] = 16'b0000000000001100;
    assign weights1[35][383] = 16'b0000000000010111;
    assign weights1[35][384] = 16'b1111111111110110;
    assign weights1[35][385] = 16'b0000000000010010;
    assign weights1[35][386] = 16'b0000000000011000;
    assign weights1[35][387] = 16'b0000000000001011;
    assign weights1[35][388] = 16'b0000000000010000;
    assign weights1[35][389] = 16'b0000000000001011;
    assign weights1[35][390] = 16'b0000000000001010;
    assign weights1[35][391] = 16'b0000000000001011;
    assign weights1[35][392] = 16'b0000000000001010;
    assign weights1[35][393] = 16'b0000000000001000;
    assign weights1[35][394] = 16'b0000000000001100;
    assign weights1[35][395] = 16'b0000000000011111;
    assign weights1[35][396] = 16'b0000000000010000;
    assign weights1[35][397] = 16'b0000000000011011;
    assign weights1[35][398] = 16'b0000000000010011;
    assign weights1[35][399] = 16'b0000000000001110;
    assign weights1[35][400] = 16'b0000000000010000;
    assign weights1[35][401] = 16'b0000000000001010;
    assign weights1[35][402] = 16'b0000000000001010;
    assign weights1[35][403] = 16'b1111111111111010;
    assign weights1[35][404] = 16'b0000000000000111;
    assign weights1[35][405] = 16'b0000000000001100;
    assign weights1[35][406] = 16'b0000000000001110;
    assign weights1[35][407] = 16'b1111111111111011;
    assign weights1[35][408] = 16'b0000000000001110;
    assign weights1[35][409] = 16'b1111111111111111;
    assign weights1[35][410] = 16'b0000000000000110;
    assign weights1[35][411] = 16'b0000000000010010;
    assign weights1[35][412] = 16'b0000000000000110;
    assign weights1[35][413] = 16'b0000000000000011;
    assign weights1[35][414] = 16'b0000000000010011;
    assign weights1[35][415] = 16'b0000000000100001;
    assign weights1[35][416] = 16'b0000000000010000;
    assign weights1[35][417] = 16'b0000000000001010;
    assign weights1[35][418] = 16'b1111111111111100;
    assign weights1[35][419] = 16'b0000000000000011;
    assign weights1[35][420] = 16'b0000000000000000;
    assign weights1[35][421] = 16'b0000000000001110;
    assign weights1[35][422] = 16'b0000000000001101;
    assign weights1[35][423] = 16'b0000000000010010;
    assign weights1[35][424] = 16'b0000000000001011;
    assign weights1[35][425] = 16'b0000000000000111;
    assign weights1[35][426] = 16'b1111111111101011;
    assign weights1[35][427] = 16'b0000000000010101;
    assign weights1[35][428] = 16'b0000000000000100;
    assign weights1[35][429] = 16'b0000000000000111;
    assign weights1[35][430] = 16'b0000000000010000;
    assign weights1[35][431] = 16'b0000000000000000;
    assign weights1[35][432] = 16'b0000000000000111;
    assign weights1[35][433] = 16'b0000000000011100;
    assign weights1[35][434] = 16'b1111111111111110;
    assign weights1[35][435] = 16'b0000000000001011;
    assign weights1[35][436] = 16'b0000000000010100;
    assign weights1[35][437] = 16'b0000000000010000;
    assign weights1[35][438] = 16'b0000000000100000;
    assign weights1[35][439] = 16'b0000000000001110;
    assign weights1[35][440] = 16'b0000000000011101;
    assign weights1[35][441] = 16'b0000000000000111;
    assign weights1[35][442] = 16'b0000000000001110;
    assign weights1[35][443] = 16'b0000000000001101;
    assign weights1[35][444] = 16'b0000000000001101;
    assign weights1[35][445] = 16'b0000000000000110;
    assign weights1[35][446] = 16'b1111111111110001;
    assign weights1[35][447] = 16'b0000000000000010;
    assign weights1[35][448] = 16'b0000000000000011;
    assign weights1[35][449] = 16'b1111111111111101;
    assign weights1[35][450] = 16'b1111111111111001;
    assign weights1[35][451] = 16'b0000000000000110;
    assign weights1[35][452] = 16'b0000000000010111;
    assign weights1[35][453] = 16'b0000000000011001;
    assign weights1[35][454] = 16'b0000000000001111;
    assign weights1[35][455] = 16'b0000000000011000;
    assign weights1[35][456] = 16'b0000000000001110;
    assign weights1[35][457] = 16'b0000000000001100;
    assign weights1[35][458] = 16'b0000000000000111;
    assign weights1[35][459] = 16'b0000000000010000;
    assign weights1[35][460] = 16'b0000000000010110;
    assign weights1[35][461] = 16'b0000000000001101;
    assign weights1[35][462] = 16'b0000000000001110;
    assign weights1[35][463] = 16'b0000000000010101;
    assign weights1[35][464] = 16'b0000000000010111;
    assign weights1[35][465] = 16'b0000000000010101;
    assign weights1[35][466] = 16'b0000000000000000;
    assign weights1[35][467] = 16'b0000000000010111;
    assign weights1[35][468] = 16'b0000000000010011;
    assign weights1[35][469] = 16'b0000000000010110;
    assign weights1[35][470] = 16'b1111111111111110;
    assign weights1[35][471] = 16'b0000000000001000;
    assign weights1[35][472] = 16'b0000000000000101;
    assign weights1[35][473] = 16'b0000000000001001;
    assign weights1[35][474] = 16'b1111111111101101;
    assign weights1[35][475] = 16'b1111111111101101;
    assign weights1[35][476] = 16'b0000000000000001;
    assign weights1[35][477] = 16'b1111111111111100;
    assign weights1[35][478] = 16'b1111111111111001;
    assign weights1[35][479] = 16'b0000000000000001;
    assign weights1[35][480] = 16'b0000000000000100;
    assign weights1[35][481] = 16'b1111111111101010;
    assign weights1[35][482] = 16'b0000000000010101;
    assign weights1[35][483] = 16'b0000000000001110;
    assign weights1[35][484] = 16'b1111111111111101;
    assign weights1[35][485] = 16'b0000000000000110;
    assign weights1[35][486] = 16'b0000000000000000;
    assign weights1[35][487] = 16'b0000000000000000;
    assign weights1[35][488] = 16'b0000000000001100;
    assign weights1[35][489] = 16'b1111111111111111;
    assign weights1[35][490] = 16'b0000000000000110;
    assign weights1[35][491] = 16'b0000000000000001;
    assign weights1[35][492] = 16'b0000000000011010;
    assign weights1[35][493] = 16'b0000000000001010;
    assign weights1[35][494] = 16'b0000000000001011;
    assign weights1[35][495] = 16'b0000000000010110;
    assign weights1[35][496] = 16'b0000000000010110;
    assign weights1[35][497] = 16'b0000000000010111;
    assign weights1[35][498] = 16'b0000000000010001;
    assign weights1[35][499] = 16'b0000000000001000;
    assign weights1[35][500] = 16'b1111111111101100;
    assign weights1[35][501] = 16'b1111111111100111;
    assign weights1[35][502] = 16'b1111111111101000;
    assign weights1[35][503] = 16'b1111111111011000;
    assign weights1[35][504] = 16'b1111111111111101;
    assign weights1[35][505] = 16'b1111111111101111;
    assign weights1[35][506] = 16'b1111111111101010;
    assign weights1[35][507] = 16'b0000000000000001;
    assign weights1[35][508] = 16'b0000000000000011;
    assign weights1[35][509] = 16'b1111111111111001;
    assign weights1[35][510] = 16'b1111111111110011;
    assign weights1[35][511] = 16'b1111111111111010;
    assign weights1[35][512] = 16'b0000000000011010;
    assign weights1[35][513] = 16'b1111111111111111;
    assign weights1[35][514] = 16'b0000000000001011;
    assign weights1[35][515] = 16'b0000000000000101;
    assign weights1[35][516] = 16'b1111111111111000;
    assign weights1[35][517] = 16'b0000000000001011;
    assign weights1[35][518] = 16'b1111111111111001;
    assign weights1[35][519] = 16'b0000000000000100;
    assign weights1[35][520] = 16'b1111111111110111;
    assign weights1[35][521] = 16'b0000000000010000;
    assign weights1[35][522] = 16'b0000000000100001;
    assign weights1[35][523] = 16'b0000000000011010;
    assign weights1[35][524] = 16'b0000000000001111;
    assign weights1[35][525] = 16'b0000000000001101;
    assign weights1[35][526] = 16'b1111111111101001;
    assign weights1[35][527] = 16'b1111111111101100;
    assign weights1[35][528] = 16'b1111111111100010;
    assign weights1[35][529] = 16'b1111111111001100;
    assign weights1[35][530] = 16'b1111111110111110;
    assign weights1[35][531] = 16'b1111111111001011;
    assign weights1[35][532] = 16'b1111111111111000;
    assign weights1[35][533] = 16'b1111111111101010;
    assign weights1[35][534] = 16'b1111111111101011;
    assign weights1[35][535] = 16'b1111111111110111;
    assign weights1[35][536] = 16'b1111111111101001;
    assign weights1[35][537] = 16'b1111111111111011;
    assign weights1[35][538] = 16'b1111111111101010;
    assign weights1[35][539] = 16'b1111111111101100;
    assign weights1[35][540] = 16'b1111111111110100;
    assign weights1[35][541] = 16'b1111111111100001;
    assign weights1[35][542] = 16'b1111111111011011;
    assign weights1[35][543] = 16'b1111111111110001;
    assign weights1[35][544] = 16'b1111111111110101;
    assign weights1[35][545] = 16'b1111111111111100;
    assign weights1[35][546] = 16'b1111111111111101;
    assign weights1[35][547] = 16'b0000000000000101;
    assign weights1[35][548] = 16'b1111111111110001;
    assign weights1[35][549] = 16'b1111111111101001;
    assign weights1[35][550] = 16'b1111111111101101;
    assign weights1[35][551] = 16'b1111111111101101;
    assign weights1[35][552] = 16'b1111111111011100;
    assign weights1[35][553] = 16'b1111111111001010;
    assign weights1[35][554] = 16'b1111111110111111;
    assign weights1[35][555] = 16'b1111111110101110;
    assign weights1[35][556] = 16'b1111111110111010;
    assign weights1[35][557] = 16'b1111111110111101;
    assign weights1[35][558] = 16'b1111111110111101;
    assign weights1[35][559] = 16'b1111111111001110;
    assign weights1[35][560] = 16'b1111111111110010;
    assign weights1[35][561] = 16'b1111111111100110;
    assign weights1[35][562] = 16'b1111111111100101;
    assign weights1[35][563] = 16'b1111111111010101;
    assign weights1[35][564] = 16'b1111111111010011;
    assign weights1[35][565] = 16'b1111111111100000;
    assign weights1[35][566] = 16'b1111111111010011;
    assign weights1[35][567] = 16'b1111111111000110;
    assign weights1[35][568] = 16'b1111111111100001;
    assign weights1[35][569] = 16'b1111111111010010;
    assign weights1[35][570] = 16'b1111111111001111;
    assign weights1[35][571] = 16'b1111111111011100;
    assign weights1[35][572] = 16'b1111111111011111;
    assign weights1[35][573] = 16'b1111111111001001;
    assign weights1[35][574] = 16'b1111111111010011;
    assign weights1[35][575] = 16'b1111111111001010;
    assign weights1[35][576] = 16'b1111111110111000;
    assign weights1[35][577] = 16'b1111111110011100;
    assign weights1[35][578] = 16'b1111111101111011;
    assign weights1[35][579] = 16'b1111111101111111;
    assign weights1[35][580] = 16'b1111111101101010;
    assign weights1[35][581] = 16'b1111111101011100;
    assign weights1[35][582] = 16'b1111111110010000;
    assign weights1[35][583] = 16'b1111111110100010;
    assign weights1[35][584] = 16'b1111111110110000;
    assign weights1[35][585] = 16'b1111111110100110;
    assign weights1[35][586] = 16'b1111111111001101;
    assign weights1[35][587] = 16'b1111111111010001;
    assign weights1[35][588] = 16'b1111111111110111;
    assign weights1[35][589] = 16'b1111111111100100;
    assign weights1[35][590] = 16'b1111111111011100;
    assign weights1[35][591] = 16'b1111111111010100;
    assign weights1[35][592] = 16'b1111111111000010;
    assign weights1[35][593] = 16'b1111111110110011;
    assign weights1[35][594] = 16'b1111111110100011;
    assign weights1[35][595] = 16'b1111111110011111;
    assign weights1[35][596] = 16'b1111111110011100;
    assign weights1[35][597] = 16'b1111111101111011;
    assign weights1[35][598] = 16'b1111111110001001;
    assign weights1[35][599] = 16'b1111111101110011;
    assign weights1[35][600] = 16'b1111111101110001;
    assign weights1[35][601] = 16'b1111111101101111;
    assign weights1[35][602] = 16'b1111111101100111;
    assign weights1[35][603] = 16'b1111111101100001;
    assign weights1[35][604] = 16'b1111111101100011;
    assign weights1[35][605] = 16'b1111111101011111;
    assign weights1[35][606] = 16'b1111111110000000;
    assign weights1[35][607] = 16'b1111111101111100;
    assign weights1[35][608] = 16'b1111111110010100;
    assign weights1[35][609] = 16'b1111111110101000;
    assign weights1[35][610] = 16'b1111111110101100;
    assign weights1[35][611] = 16'b1111111111000000;
    assign weights1[35][612] = 16'b1111111111010110;
    assign weights1[35][613] = 16'b1111111111010011;
    assign weights1[35][614] = 16'b1111111111011011;
    assign weights1[35][615] = 16'b1111111111100110;
    assign weights1[35][616] = 16'b1111111111110110;
    assign weights1[35][617] = 16'b1111111111101111;
    assign weights1[35][618] = 16'b1111111111100101;
    assign weights1[35][619] = 16'b1111111111100000;
    assign weights1[35][620] = 16'b1111111111011011;
    assign weights1[35][621] = 16'b1111111111011100;
    assign weights1[35][622] = 16'b1111111111001010;
    assign weights1[35][623] = 16'b1111111111000011;
    assign weights1[35][624] = 16'b1111111111000000;
    assign weights1[35][625] = 16'b1111111110111000;
    assign weights1[35][626] = 16'b1111111111000000;
    assign weights1[35][627] = 16'b1111111110100111;
    assign weights1[35][628] = 16'b1111111110111011;
    assign weights1[35][629] = 16'b1111111110100011;
    assign weights1[35][630] = 16'b1111111110101000;
    assign weights1[35][631] = 16'b1111111110011100;
    assign weights1[35][632] = 16'b1111111110101010;
    assign weights1[35][633] = 16'b1111111110100101;
    assign weights1[35][634] = 16'b1111111110110001;
    assign weights1[35][635] = 16'b1111111110101010;
    assign weights1[35][636] = 16'b1111111111000010;
    assign weights1[35][637] = 16'b1111111111000010;
    assign weights1[35][638] = 16'b1111111111010011;
    assign weights1[35][639] = 16'b1111111111010000;
    assign weights1[35][640] = 16'b1111111111100100;
    assign weights1[35][641] = 16'b1111111111101100;
    assign weights1[35][642] = 16'b1111111111101111;
    assign weights1[35][643] = 16'b1111111111101010;
    assign weights1[35][644] = 16'b0000000000000000;
    assign weights1[35][645] = 16'b1111111111111001;
    assign weights1[35][646] = 16'b1111111111111001;
    assign weights1[35][647] = 16'b1111111111110101;
    assign weights1[35][648] = 16'b1111111111110001;
    assign weights1[35][649] = 16'b1111111111101111;
    assign weights1[35][650] = 16'b1111111111101010;
    assign weights1[35][651] = 16'b1111111111100101;
    assign weights1[35][652] = 16'b1111111111100110;
    assign weights1[35][653] = 16'b1111111111010101;
    assign weights1[35][654] = 16'b1111111111100101;
    assign weights1[35][655] = 16'b1111111111010000;
    assign weights1[35][656] = 16'b1111111111010101;
    assign weights1[35][657] = 16'b1111111111001101;
    assign weights1[35][658] = 16'b1111111111001001;
    assign weights1[35][659] = 16'b1111111110111010;
    assign weights1[35][660] = 16'b1111111111001010;
    assign weights1[35][661] = 16'b1111111111000111;
    assign weights1[35][662] = 16'b1111111111001011;
    assign weights1[35][663] = 16'b1111111110111011;
    assign weights1[35][664] = 16'b1111111111001111;
    assign weights1[35][665] = 16'b1111111111010111;
    assign weights1[35][666] = 16'b1111111111011010;
    assign weights1[35][667] = 16'b1111111111101110;
    assign weights1[35][668] = 16'b1111111111101100;
    assign weights1[35][669] = 16'b1111111111110010;
    assign weights1[35][670] = 16'b1111111111110111;
    assign weights1[35][671] = 16'b1111111111110100;
    assign weights1[35][672] = 16'b0000000000000011;
    assign weights1[35][673] = 16'b0000000000000000;
    assign weights1[35][674] = 16'b1111111111111010;
    assign weights1[35][675] = 16'b1111111111111011;
    assign weights1[35][676] = 16'b1111111111111110;
    assign weights1[35][677] = 16'b0000000000000100;
    assign weights1[35][678] = 16'b0000000000000001;
    assign weights1[35][679] = 16'b1111111111110100;
    assign weights1[35][680] = 16'b1111111111111111;
    assign weights1[35][681] = 16'b1111111111110110;
    assign weights1[35][682] = 16'b1111111111010001;
    assign weights1[35][683] = 16'b1111111111100001;
    assign weights1[35][684] = 16'b1111111111101000;
    assign weights1[35][685] = 16'b1111111111001111;
    assign weights1[35][686] = 16'b1111111111011100;
    assign weights1[35][687] = 16'b1111111111101010;
    assign weights1[35][688] = 16'b1111111111100000;
    assign weights1[35][689] = 16'b1111111111011101;
    assign weights1[35][690] = 16'b1111111111100010;
    assign weights1[35][691] = 16'b1111111111011000;
    assign weights1[35][692] = 16'b1111111111010110;
    assign weights1[35][693] = 16'b1111111111010110;
    assign weights1[35][694] = 16'b1111111111101111;
    assign weights1[35][695] = 16'b1111111111110000;
    assign weights1[35][696] = 16'b1111111111111001;
    assign weights1[35][697] = 16'b1111111111110101;
    assign weights1[35][698] = 16'b1111111111111001;
    assign weights1[35][699] = 16'b1111111111111011;
    assign weights1[35][700] = 16'b0000000000000011;
    assign weights1[35][701] = 16'b1111111111111110;
    assign weights1[35][702] = 16'b1111111111111011;
    assign weights1[35][703] = 16'b0000000000000001;
    assign weights1[35][704] = 16'b1111111111111110;
    assign weights1[35][705] = 16'b0000000000000011;
    assign weights1[35][706] = 16'b0000000000000010;
    assign weights1[35][707] = 16'b0000000000000000;
    assign weights1[35][708] = 16'b1111111111111011;
    assign weights1[35][709] = 16'b1111111111101110;
    assign weights1[35][710] = 16'b1111111111101011;
    assign weights1[35][711] = 16'b1111111111110100;
    assign weights1[35][712] = 16'b1111111111101101;
    assign weights1[35][713] = 16'b1111111111101000;
    assign weights1[35][714] = 16'b1111111111100111;
    assign weights1[35][715] = 16'b1111111111110111;
    assign weights1[35][716] = 16'b1111111111100111;
    assign weights1[35][717] = 16'b1111111111100110;
    assign weights1[35][718] = 16'b1111111111110110;
    assign weights1[35][719] = 16'b1111111111011101;
    assign weights1[35][720] = 16'b1111111111100101;
    assign weights1[35][721] = 16'b1111111111111000;
    assign weights1[35][722] = 16'b1111111111111001;
    assign weights1[35][723] = 16'b1111111111110010;
    assign weights1[35][724] = 16'b1111111111111000;
    assign weights1[35][725] = 16'b1111111111111010;
    assign weights1[35][726] = 16'b1111111111111111;
    assign weights1[35][727] = 16'b1111111111111101;
    assign weights1[35][728] = 16'b0000000000000001;
    assign weights1[35][729] = 16'b0000000000000001;
    assign weights1[35][730] = 16'b0000000000000001;
    assign weights1[35][731] = 16'b0000000000000010;
    assign weights1[35][732] = 16'b1111111111111111;
    assign weights1[35][733] = 16'b1111111111111010;
    assign weights1[35][734] = 16'b1111111111111100;
    assign weights1[35][735] = 16'b1111111111111111;
    assign weights1[35][736] = 16'b1111111111101111;
    assign weights1[35][737] = 16'b1111111111111000;
    assign weights1[35][738] = 16'b1111111111111010;
    assign weights1[35][739] = 16'b1111111111110100;
    assign weights1[35][740] = 16'b1111111111110111;
    assign weights1[35][741] = 16'b1111111111110011;
    assign weights1[35][742] = 16'b1111111111111010;
    assign weights1[35][743] = 16'b1111111111111110;
    assign weights1[35][744] = 16'b1111111111101110;
    assign weights1[35][745] = 16'b1111111111111000;
    assign weights1[35][746] = 16'b1111111111111010;
    assign weights1[35][747] = 16'b1111111111110000;
    assign weights1[35][748] = 16'b1111111111101000;
    assign weights1[35][749] = 16'b1111111111111100;
    assign weights1[35][750] = 16'b1111111111111100;
    assign weights1[35][751] = 16'b1111111111111011;
    assign weights1[35][752] = 16'b1111111111111010;
    assign weights1[35][753] = 16'b1111111111111011;
    assign weights1[35][754] = 16'b1111111111111111;
    assign weights1[35][755] = 16'b0000000000000000;
    assign weights1[35][756] = 16'b0000000000000000;
    assign weights1[35][757] = 16'b0000000000000000;
    assign weights1[35][758] = 16'b0000000000000001;
    assign weights1[35][759] = 16'b0000000000000001;
    assign weights1[35][760] = 16'b1111111111111100;
    assign weights1[35][761] = 16'b1111111111111101;
    assign weights1[35][762] = 16'b0000000000000000;
    assign weights1[35][763] = 16'b1111111111110010;
    assign weights1[35][764] = 16'b1111111111110010;
    assign weights1[35][765] = 16'b1111111111111100;
    assign weights1[35][766] = 16'b1111111111110111;
    assign weights1[35][767] = 16'b1111111111111001;
    assign weights1[35][768] = 16'b1111111111111100;
    assign weights1[35][769] = 16'b1111111111111111;
    assign weights1[35][770] = 16'b1111111111111010;
    assign weights1[35][771] = 16'b1111111111110111;
    assign weights1[35][772] = 16'b1111111111111001;
    assign weights1[35][773] = 16'b0000000000000000;
    assign weights1[35][774] = 16'b1111111111111111;
    assign weights1[35][775] = 16'b0000000000000000;
    assign weights1[35][776] = 16'b0000000000000000;
    assign weights1[35][777] = 16'b0000000000000000;
    assign weights1[35][778] = 16'b0000000000000000;
    assign weights1[35][779] = 16'b1111111111111110;
    assign weights1[35][780] = 16'b1111111111111100;
    assign weights1[35][781] = 16'b1111111111111110;
    assign weights1[35][782] = 16'b0000000000000001;
    assign weights1[35][783] = 16'b0000000000000000;
    assign weights1[36][0] = 16'b0000000000000000;
    assign weights1[36][1] = 16'b0000000000000000;
    assign weights1[36][2] = 16'b0000000000000000;
    assign weights1[36][3] = 16'b0000000000000010;
    assign weights1[36][4] = 16'b0000000000000000;
    assign weights1[36][5] = 16'b1111111111111101;
    assign weights1[36][6] = 16'b1111111111111011;
    assign weights1[36][7] = 16'b1111111111111111;
    assign weights1[36][8] = 16'b1111111111111101;
    assign weights1[36][9] = 16'b1111111111111101;
    assign weights1[36][10] = 16'b1111111111111010;
    assign weights1[36][11] = 16'b0000000000000010;
    assign weights1[36][12] = 16'b1111111111111110;
    assign weights1[36][13] = 16'b1111111111111010;
    assign weights1[36][14] = 16'b1111111111111101;
    assign weights1[36][15] = 16'b1111111111111011;
    assign weights1[36][16] = 16'b1111111111110110;
    assign weights1[36][17] = 16'b1111111111110011;
    assign weights1[36][18] = 16'b1111111111101101;
    assign weights1[36][19] = 16'b1111111111101101;
    assign weights1[36][20] = 16'b1111111111110001;
    assign weights1[36][21] = 16'b1111111111111010;
    assign weights1[36][22] = 16'b0000000000000000;
    assign weights1[36][23] = 16'b0000000000000000;
    assign weights1[36][24] = 16'b0000000000000001;
    assign weights1[36][25] = 16'b0000000000000000;
    assign weights1[36][26] = 16'b0000000000000000;
    assign weights1[36][27] = 16'b0000000000000000;
    assign weights1[36][28] = 16'b0000000000000000;
    assign weights1[36][29] = 16'b0000000000000000;
    assign weights1[36][30] = 16'b1111111111111100;
    assign weights1[36][31] = 16'b1111111111111101;
    assign weights1[36][32] = 16'b1111111111111100;
    assign weights1[36][33] = 16'b1111111111110111;
    assign weights1[36][34] = 16'b1111111111111010;
    assign weights1[36][35] = 16'b1111111111111111;
    assign weights1[36][36] = 16'b1111111111111011;
    assign weights1[36][37] = 16'b1111111111111101;
    assign weights1[36][38] = 16'b1111111111111100;
    assign weights1[36][39] = 16'b0000000000000011;
    assign weights1[36][40] = 16'b1111111111111101;
    assign weights1[36][41] = 16'b1111111111111100;
    assign weights1[36][42] = 16'b0000000000000000;
    assign weights1[36][43] = 16'b1111111111111010;
    assign weights1[36][44] = 16'b1111111111111101;
    assign weights1[36][45] = 16'b1111111111100011;
    assign weights1[36][46] = 16'b1111111111111100;
    assign weights1[36][47] = 16'b1111111111101110;
    assign weights1[36][48] = 16'b1111111111111101;
    assign weights1[36][49] = 16'b1111111111111110;
    assign weights1[36][50] = 16'b1111111111111101;
    assign weights1[36][51] = 16'b0000000000000000;
    assign weights1[36][52] = 16'b1111111111111110;
    assign weights1[36][53] = 16'b0000000000000011;
    assign weights1[36][54] = 16'b1111111111111101;
    assign weights1[36][55] = 16'b0000000000000000;
    assign weights1[36][56] = 16'b0000000000000001;
    assign weights1[36][57] = 16'b1111111111111100;
    assign weights1[36][58] = 16'b1111111111111001;
    assign weights1[36][59] = 16'b1111111111111000;
    assign weights1[36][60] = 16'b1111111111110010;
    assign weights1[36][61] = 16'b1111111111110001;
    assign weights1[36][62] = 16'b1111111111110100;
    assign weights1[36][63] = 16'b1111111111111110;
    assign weights1[36][64] = 16'b1111111111110111;
    assign weights1[36][65] = 16'b1111111111111100;
    assign weights1[36][66] = 16'b0000000000001111;
    assign weights1[36][67] = 16'b0000000000000001;
    assign weights1[36][68] = 16'b1111111111111110;
    assign weights1[36][69] = 16'b0000000000000111;
    assign weights1[36][70] = 16'b0000000000000110;
    assign weights1[36][71] = 16'b1111111111111111;
    assign weights1[36][72] = 16'b0000000000000000;
    assign weights1[36][73] = 16'b0000000000001001;
    assign weights1[36][74] = 16'b0000000000000100;
    assign weights1[36][75] = 16'b0000000000001011;
    assign weights1[36][76] = 16'b1111111111111100;
    assign weights1[36][77] = 16'b1111111111111100;
    assign weights1[36][78] = 16'b1111111111110110;
    assign weights1[36][79] = 16'b1111111111110010;
    assign weights1[36][80] = 16'b1111111111111011;
    assign weights1[36][81] = 16'b0000000000000011;
    assign weights1[36][82] = 16'b0000000000000000;
    assign weights1[36][83] = 16'b1111111111111011;
    assign weights1[36][84] = 16'b0000000000000001;
    assign weights1[36][85] = 16'b0000000000000000;
    assign weights1[36][86] = 16'b1111111111111011;
    assign weights1[36][87] = 16'b1111111111110110;
    assign weights1[36][88] = 16'b1111111111110001;
    assign weights1[36][89] = 16'b1111111111110100;
    assign weights1[36][90] = 16'b1111111111110001;
    assign weights1[36][91] = 16'b1111111111111000;
    assign weights1[36][92] = 16'b1111111111111001;
    assign weights1[36][93] = 16'b1111111111111001;
    assign weights1[36][94] = 16'b1111111111111111;
    assign weights1[36][95] = 16'b1111111111111100;
    assign weights1[36][96] = 16'b0000000000000110;
    assign weights1[36][97] = 16'b0000000000000011;
    assign weights1[36][98] = 16'b0000000000000110;
    assign weights1[36][99] = 16'b1111111111111001;
    assign weights1[36][100] = 16'b1111111111110011;
    assign weights1[36][101] = 16'b1111111111111110;
    assign weights1[36][102] = 16'b0000000000000111;
    assign weights1[36][103] = 16'b0000000000001001;
    assign weights1[36][104] = 16'b0000000000001000;
    assign weights1[36][105] = 16'b1111111111111001;
    assign weights1[36][106] = 16'b1111111111110001;
    assign weights1[36][107] = 16'b1111111111110011;
    assign weights1[36][108] = 16'b1111111111110110;
    assign weights1[36][109] = 16'b0000000000000101;
    assign weights1[36][110] = 16'b0000000000000010;
    assign weights1[36][111] = 16'b1111111111111110;
    assign weights1[36][112] = 16'b1111111111111110;
    assign weights1[36][113] = 16'b1111111111111100;
    assign weights1[36][114] = 16'b1111111111110101;
    assign weights1[36][115] = 16'b1111111111101011;
    assign weights1[36][116] = 16'b1111111111101111;
    assign weights1[36][117] = 16'b1111111111100110;
    assign weights1[36][118] = 16'b1111111111110101;
    assign weights1[36][119] = 16'b1111111111101101;
    assign weights1[36][120] = 16'b1111111111111100;
    assign weights1[36][121] = 16'b1111111111111111;
    assign weights1[36][122] = 16'b0000000000000001;
    assign weights1[36][123] = 16'b1111111111111000;
    assign weights1[36][124] = 16'b1111111111110011;
    assign weights1[36][125] = 16'b1111111111111010;
    assign weights1[36][126] = 16'b1111111111111111;
    assign weights1[36][127] = 16'b0000000000000001;
    assign weights1[36][128] = 16'b0000000000000001;
    assign weights1[36][129] = 16'b0000000000000110;
    assign weights1[36][130] = 16'b1111111111111001;
    assign weights1[36][131] = 16'b1111111111110111;
    assign weights1[36][132] = 16'b1111111111110110;
    assign weights1[36][133] = 16'b1111111111110101;
    assign weights1[36][134] = 16'b1111111111110111;
    assign weights1[36][135] = 16'b1111111111110010;
    assign weights1[36][136] = 16'b1111111111101110;
    assign weights1[36][137] = 16'b0000000000001001;
    assign weights1[36][138] = 16'b0000000000000001;
    assign weights1[36][139] = 16'b0000000000000011;
    assign weights1[36][140] = 16'b1111111111111101;
    assign weights1[36][141] = 16'b1111111111111100;
    assign weights1[36][142] = 16'b1111111111110111;
    assign weights1[36][143] = 16'b1111111111101111;
    assign weights1[36][144] = 16'b1111111111100110;
    assign weights1[36][145] = 16'b1111111111110100;
    assign weights1[36][146] = 16'b1111111111110111;
    assign weights1[36][147] = 16'b0000000000000011;
    assign weights1[36][148] = 16'b1111111111110101;
    assign weights1[36][149] = 16'b1111111111111000;
    assign weights1[36][150] = 16'b1111111111100010;
    assign weights1[36][151] = 16'b1111111111110110;
    assign weights1[36][152] = 16'b1111111111111110;
    assign weights1[36][153] = 16'b1111111111011010;
    assign weights1[36][154] = 16'b0000000000010010;
    assign weights1[36][155] = 16'b0000000000000001;
    assign weights1[36][156] = 16'b1111111111111000;
    assign weights1[36][157] = 16'b1111111111101000;
    assign weights1[36][158] = 16'b1111111111111001;
    assign weights1[36][159] = 16'b1111111111111001;
    assign weights1[36][160] = 16'b0000000000000111;
    assign weights1[36][161] = 16'b1111111111111110;
    assign weights1[36][162] = 16'b0000000000010110;
    assign weights1[36][163] = 16'b1111111111110001;
    assign weights1[36][164] = 16'b1111111111110111;
    assign weights1[36][165] = 16'b0000000000000011;
    assign weights1[36][166] = 16'b1111111111111000;
    assign weights1[36][167] = 16'b0000000000000000;
    assign weights1[36][168] = 16'b1111111111111110;
    assign weights1[36][169] = 16'b1111111111111111;
    assign weights1[36][170] = 16'b1111111111111011;
    assign weights1[36][171] = 16'b1111111111110011;
    assign weights1[36][172] = 16'b1111111111100101;
    assign weights1[36][173] = 16'b1111111111101010;
    assign weights1[36][174] = 16'b0000000000000000;
    assign weights1[36][175] = 16'b1111111111110000;
    assign weights1[36][176] = 16'b0000000000001100;
    assign weights1[36][177] = 16'b1111111111111100;
    assign weights1[36][178] = 16'b1111111111110111;
    assign weights1[36][179] = 16'b1111111111110000;
    assign weights1[36][180] = 16'b1111111111101111;
    assign weights1[36][181] = 16'b1111111111111101;
    assign weights1[36][182] = 16'b1111111111101111;
    assign weights1[36][183] = 16'b0000000000000000;
    assign weights1[36][184] = 16'b1111111111111100;
    assign weights1[36][185] = 16'b0000000000000001;
    assign weights1[36][186] = 16'b0000000000001000;
    assign weights1[36][187] = 16'b0000000000000010;
    assign weights1[36][188] = 16'b0000000000001000;
    assign weights1[36][189] = 16'b1111111111111101;
    assign weights1[36][190] = 16'b1111111111111111;
    assign weights1[36][191] = 16'b1111111111110011;
    assign weights1[36][192] = 16'b0000000000001101;
    assign weights1[36][193] = 16'b0000000000000111;
    assign weights1[36][194] = 16'b1111111111111101;
    assign weights1[36][195] = 16'b0000000000000000;
    assign weights1[36][196] = 16'b1111111111111110;
    assign weights1[36][197] = 16'b1111111111110111;
    assign weights1[36][198] = 16'b1111111111111010;
    assign weights1[36][199] = 16'b1111111111110001;
    assign weights1[36][200] = 16'b1111111111101001;
    assign weights1[36][201] = 16'b1111111111110001;
    assign weights1[36][202] = 16'b1111111111110111;
    assign weights1[36][203] = 16'b0000000000001100;
    assign weights1[36][204] = 16'b0000000000001101;
    assign weights1[36][205] = 16'b0000000000000001;
    assign weights1[36][206] = 16'b0000000000001000;
    assign weights1[36][207] = 16'b1111111111110101;
    assign weights1[36][208] = 16'b1111111111110100;
    assign weights1[36][209] = 16'b0000000000000000;
    assign weights1[36][210] = 16'b1111111111110010;
    assign weights1[36][211] = 16'b0000000000010010;
    assign weights1[36][212] = 16'b0000000000010100;
    assign weights1[36][213] = 16'b0000000000010111;
    assign weights1[36][214] = 16'b1111111111111101;
    assign weights1[36][215] = 16'b0000000000000110;
    assign weights1[36][216] = 16'b0000000000000111;
    assign weights1[36][217] = 16'b1111111111110010;
    assign weights1[36][218] = 16'b1111111111111010;
    assign weights1[36][219] = 16'b0000000000000110;
    assign weights1[36][220] = 16'b1111111111110101;
    assign weights1[36][221] = 16'b0000000000001010;
    assign weights1[36][222] = 16'b1111111111101111;
    assign weights1[36][223] = 16'b1111111111111110;
    assign weights1[36][224] = 16'b1111111111111001;
    assign weights1[36][225] = 16'b1111111111110010;
    assign weights1[36][226] = 16'b1111111111111101;
    assign weights1[36][227] = 16'b1111111111110010;
    assign weights1[36][228] = 16'b1111111111111110;
    assign weights1[36][229] = 16'b1111111111111000;
    assign weights1[36][230] = 16'b1111111111111100;
    assign weights1[36][231] = 16'b0000000000000001;
    assign weights1[36][232] = 16'b0000000000000001;
    assign weights1[36][233] = 16'b0000000000000100;
    assign weights1[36][234] = 16'b0000000000001011;
    assign weights1[36][235] = 16'b0000000000001100;
    assign weights1[36][236] = 16'b1111111111110101;
    assign weights1[36][237] = 16'b0000000000001011;
    assign weights1[36][238] = 16'b1111111111110101;
    assign weights1[36][239] = 16'b1111111111111101;
    assign weights1[36][240] = 16'b1111111111111111;
    assign weights1[36][241] = 16'b1111111111101011;
    assign weights1[36][242] = 16'b0000000000000010;
    assign weights1[36][243] = 16'b0000000000100001;
    assign weights1[36][244] = 16'b0000000000000010;
    assign weights1[36][245] = 16'b1111111111101001;
    assign weights1[36][246] = 16'b1111111111110000;
    assign weights1[36][247] = 16'b0000000000000100;
    assign weights1[36][248] = 16'b0000000000000100;
    assign weights1[36][249] = 16'b1111111111110001;
    assign weights1[36][250] = 16'b0000000000001010;
    assign weights1[36][251] = 16'b0000000000001110;
    assign weights1[36][252] = 16'b1111111111110100;
    assign weights1[36][253] = 16'b0000000000000000;
    assign weights1[36][254] = 16'b0000000000000101;
    assign weights1[36][255] = 16'b1111111111110111;
    assign weights1[36][256] = 16'b1111111111101001;
    assign weights1[36][257] = 16'b1111111111100110;
    assign weights1[36][258] = 16'b1111111111110110;
    assign weights1[36][259] = 16'b1111111111110000;
    assign weights1[36][260] = 16'b1111111111111000;
    assign weights1[36][261] = 16'b0000000000001111;
    assign weights1[36][262] = 16'b0000000000000101;
    assign weights1[36][263] = 16'b0000000000000011;
    assign weights1[36][264] = 16'b0000000000000001;
    assign weights1[36][265] = 16'b1111111111101011;
    assign weights1[36][266] = 16'b1111111111101100;
    assign weights1[36][267] = 16'b1111111111111110;
    assign weights1[36][268] = 16'b0000000000001111;
    assign weights1[36][269] = 16'b0000000000010011;
    assign weights1[36][270] = 16'b0000000000001100;
    assign weights1[36][271] = 16'b0000000000001001;
    assign weights1[36][272] = 16'b0000000000011000;
    assign weights1[36][273] = 16'b0000000000011100;
    assign weights1[36][274] = 16'b1111111111111011;
    assign weights1[36][275] = 16'b0000000000010100;
    assign weights1[36][276] = 16'b1111111111111110;
    assign weights1[36][277] = 16'b1111111111111010;
    assign weights1[36][278] = 16'b0000000000000001;
    assign weights1[36][279] = 16'b0000000000000000;
    assign weights1[36][280] = 16'b1111111111111011;
    assign weights1[36][281] = 16'b0000000000000111;
    assign weights1[36][282] = 16'b1111111111111011;
    assign weights1[36][283] = 16'b1111111111110101;
    assign weights1[36][284] = 16'b1111111111110000;
    assign weights1[36][285] = 16'b1111111111110101;
    assign weights1[36][286] = 16'b1111111111101001;
    assign weights1[36][287] = 16'b1111111111111100;
    assign weights1[36][288] = 16'b1111111111110000;
    assign weights1[36][289] = 16'b1111111111110110;
    assign weights1[36][290] = 16'b1111111111111111;
    assign weights1[36][291] = 16'b0000000000010011;
    assign weights1[36][292] = 16'b1111111111101001;
    assign weights1[36][293] = 16'b1111111111011001;
    assign weights1[36][294] = 16'b0000000000000011;
    assign weights1[36][295] = 16'b0000000000000000;
    assign weights1[36][296] = 16'b0000000000000010;
    assign weights1[36][297] = 16'b0000000000001110;
    assign weights1[36][298] = 16'b0000000000000111;
    assign weights1[36][299] = 16'b0000000000000110;
    assign weights1[36][300] = 16'b0000000000001100;
    assign weights1[36][301] = 16'b0000000000010011;
    assign weights1[36][302] = 16'b0000000000010111;
    assign weights1[36][303] = 16'b0000000000011101;
    assign weights1[36][304] = 16'b0000000000010100;
    assign weights1[36][305] = 16'b0000000000001110;
    assign weights1[36][306] = 16'b0000000000001011;
    assign weights1[36][307] = 16'b0000000000001100;
    assign weights1[36][308] = 16'b1111111111111101;
    assign weights1[36][309] = 16'b1111111111111101;
    assign weights1[36][310] = 16'b0000000000000000;
    assign weights1[36][311] = 16'b1111111111101100;
    assign weights1[36][312] = 16'b1111111111100011;
    assign weights1[36][313] = 16'b1111111111100110;
    assign weights1[36][314] = 16'b0000000000001001;
    assign weights1[36][315] = 16'b1111111111110111;
    assign weights1[36][316] = 16'b0000000000000111;
    assign weights1[36][317] = 16'b0000000000010110;
    assign weights1[36][318] = 16'b0000000000010111;
    assign weights1[36][319] = 16'b0000000000001000;
    assign weights1[36][320] = 16'b0000000000000001;
    assign weights1[36][321] = 16'b1111111111101011;
    assign weights1[36][322] = 16'b1111111111110101;
    assign weights1[36][323] = 16'b1111111111100101;
    assign weights1[36][324] = 16'b0000000000000000;
    assign weights1[36][325] = 16'b0000000000000101;
    assign weights1[36][326] = 16'b0000000000000110;
    assign weights1[36][327] = 16'b0000000000001110;
    assign weights1[36][328] = 16'b0000000000000100;
    assign weights1[36][329] = 16'b0000000000000111;
    assign weights1[36][330] = 16'b0000000000011100;
    assign weights1[36][331] = 16'b0000000000100011;
    assign weights1[36][332] = 16'b0000000000100110;
    assign weights1[36][333] = 16'b0000000000011000;
    assign weights1[36][334] = 16'b0000000000011000;
    assign weights1[36][335] = 16'b0000000000010000;
    assign weights1[36][336] = 16'b1111111111111111;
    assign weights1[36][337] = 16'b0000000000001011;
    assign weights1[36][338] = 16'b1111111111111100;
    assign weights1[36][339] = 16'b1111111111111000;
    assign weights1[36][340] = 16'b1111111111110010;
    assign weights1[36][341] = 16'b1111111111100011;
    assign weights1[36][342] = 16'b1111111111110001;
    assign weights1[36][343] = 16'b1111111111111100;
    assign weights1[36][344] = 16'b0000000000000111;
    assign weights1[36][345] = 16'b0000000000001000;
    assign weights1[36][346] = 16'b0000000000010111;
    assign weights1[36][347] = 16'b0000000000001000;
    assign weights1[36][348] = 16'b0000000000001010;
    assign weights1[36][349] = 16'b1111111111110110;
    assign weights1[36][350] = 16'b1111111111001101;
    assign weights1[36][351] = 16'b1111111111101101;
    assign weights1[36][352] = 16'b1111111111101010;
    assign weights1[36][353] = 16'b0000000000000100;
    assign weights1[36][354] = 16'b0000000000000101;
    assign weights1[36][355] = 16'b0000000000011101;
    assign weights1[36][356] = 16'b0000000000010101;
    assign weights1[36][357] = 16'b0000000000000000;
    assign weights1[36][358] = 16'b0000000000000101;
    assign weights1[36][359] = 16'b0000000000011110;
    assign weights1[36][360] = 16'b0000000000100011;
    assign weights1[36][361] = 16'b0000000000001111;
    assign weights1[36][362] = 16'b0000000000010110;
    assign weights1[36][363] = 16'b0000000000001001;
    assign weights1[36][364] = 16'b1111111111111100;
    assign weights1[36][365] = 16'b0000000000001100;
    assign weights1[36][366] = 16'b0000000000010000;
    assign weights1[36][367] = 16'b0000000000000010;
    assign weights1[36][368] = 16'b1111111111110011;
    assign weights1[36][369] = 16'b1111111111111110;
    assign weights1[36][370] = 16'b1111111111110101;
    assign weights1[36][371] = 16'b1111111111100110;
    assign weights1[36][372] = 16'b0000000000001100;
    assign weights1[36][373] = 16'b0000000000001010;
    assign weights1[36][374] = 16'b0000000000100001;
    assign weights1[36][375] = 16'b0000000000101000;
    assign weights1[36][376] = 16'b1111111111111111;
    assign weights1[36][377] = 16'b1111111111010000;
    assign weights1[36][378] = 16'b1111111111001101;
    assign weights1[36][379] = 16'b1111111111011000;
    assign weights1[36][380] = 16'b1111111111110101;
    assign weights1[36][381] = 16'b0000000000011001;
    assign weights1[36][382] = 16'b0000000000100001;
    assign weights1[36][383] = 16'b0000000000010000;
    assign weights1[36][384] = 16'b0000000000100001;
    assign weights1[36][385] = 16'b0000000000110000;
    assign weights1[36][386] = 16'b0000000000110111;
    assign weights1[36][387] = 16'b0000000000111010;
    assign weights1[36][388] = 16'b0000000000011110;
    assign weights1[36][389] = 16'b0000000000001100;
    assign weights1[36][390] = 16'b0000000000001000;
    assign weights1[36][391] = 16'b1111111111111000;
    assign weights1[36][392] = 16'b0000000000001001;
    assign weights1[36][393] = 16'b0000000000000111;
    assign weights1[36][394] = 16'b0000000000010001;
    assign weights1[36][395] = 16'b0000000000000100;
    assign weights1[36][396] = 16'b1111111111111100;
    assign weights1[36][397] = 16'b1111111111110010;
    assign weights1[36][398] = 16'b1111111111110110;
    assign weights1[36][399] = 16'b0000000000001100;
    assign weights1[36][400] = 16'b0000000000010000;
    assign weights1[36][401] = 16'b0000000000011001;
    assign weights1[36][402] = 16'b0000000000011010;
    assign weights1[36][403] = 16'b0000000000001100;
    assign weights1[36][404] = 16'b1111111111110110;
    assign weights1[36][405] = 16'b1111111111101001;
    assign weights1[36][406] = 16'b1111111110100110;
    assign weights1[36][407] = 16'b1111111110110110;
    assign weights1[36][408] = 16'b1111111111101000;
    assign weights1[36][409] = 16'b1111111111101100;
    assign weights1[36][410] = 16'b1111111111111001;
    assign weights1[36][411] = 16'b0000000000100010;
    assign weights1[36][412] = 16'b0000000000100111;
    assign weights1[36][413] = 16'b0000000000110001;
    assign weights1[36][414] = 16'b0000000000010110;
    assign weights1[36][415] = 16'b0000000000011111;
    assign weights1[36][416] = 16'b0000000000001101;
    assign weights1[36][417] = 16'b1111111111111100;
    assign weights1[36][418] = 16'b1111111111110001;
    assign weights1[36][419] = 16'b1111111111101110;
    assign weights1[36][420] = 16'b0000000000010010;
    assign weights1[36][421] = 16'b0000000000000100;
    assign weights1[36][422] = 16'b0000000000010000;
    assign weights1[36][423] = 16'b0000000000010111;
    assign weights1[36][424] = 16'b0000000000000111;
    assign weights1[36][425] = 16'b0000000000001110;
    assign weights1[36][426] = 16'b1111111111110101;
    assign weights1[36][427] = 16'b0000000000000111;
    assign weights1[36][428] = 16'b1111111111111001;
    assign weights1[36][429] = 16'b0000000000010111;
    assign weights1[36][430] = 16'b0000000000010100;
    assign weights1[36][431] = 16'b0000000000100010;
    assign weights1[36][432] = 16'b0000000000001010;
    assign weights1[36][433] = 16'b1111111111110100;
    assign weights1[36][434] = 16'b1111111110111100;
    assign weights1[36][435] = 16'b1111111110010010;
    assign weights1[36][436] = 16'b1111111111001000;
    assign weights1[36][437] = 16'b1111111111011000;
    assign weights1[36][438] = 16'b0000000000000110;
    assign weights1[36][439] = 16'b1111111111111010;
    assign weights1[36][440] = 16'b0000000000001000;
    assign weights1[36][441] = 16'b0000000000001011;
    assign weights1[36][442] = 16'b1111111111110000;
    assign weights1[36][443] = 16'b0000000000000110;
    assign weights1[36][444] = 16'b1111111111101011;
    assign weights1[36][445] = 16'b1111111111101101;
    assign weights1[36][446] = 16'b1111111111101101;
    assign weights1[36][447] = 16'b1111111111100101;
    assign weights1[36][448] = 16'b0000000000000101;
    assign weights1[36][449] = 16'b1111111111111010;
    assign weights1[36][450] = 16'b0000000000011001;
    assign weights1[36][451] = 16'b0000000000010011;
    assign weights1[36][452] = 16'b0000000000000010;
    assign weights1[36][453] = 16'b0000000000000011;
    assign weights1[36][454] = 16'b0000000000001111;
    assign weights1[36][455] = 16'b0000000000010011;
    assign weights1[36][456] = 16'b0000000000000110;
    assign weights1[36][457] = 16'b0000000000001101;
    assign weights1[36][458] = 16'b0000000000011100;
    assign weights1[36][459] = 16'b0000000000010110;
    assign weights1[36][460] = 16'b0000000000011011;
    assign weights1[36][461] = 16'b0000000000000101;
    assign weights1[36][462] = 16'b1111111111001111;
    assign weights1[36][463] = 16'b1111111110000111;
    assign weights1[36][464] = 16'b1111111110001111;
    assign weights1[36][465] = 16'b1111111110100000;
    assign weights1[36][466] = 16'b1111111110100111;
    assign weights1[36][467] = 16'b1111111110111100;
    assign weights1[36][468] = 16'b1111111110111101;
    assign weights1[36][469] = 16'b1111111110111000;
    assign weights1[36][470] = 16'b1111111111001011;
    assign weights1[36][471] = 16'b1111111111001111;
    assign weights1[36][472] = 16'b1111111111011010;
    assign weights1[36][473] = 16'b1111111111010101;
    assign weights1[36][474] = 16'b1111111111100100;
    assign weights1[36][475] = 16'b1111111111100110;
    assign weights1[36][476] = 16'b0000000000000100;
    assign weights1[36][477] = 16'b0000000000001100;
    assign weights1[36][478] = 16'b0000000000011010;
    assign weights1[36][479] = 16'b0000000000010001;
    assign weights1[36][480] = 16'b0000000000010001;
    assign weights1[36][481] = 16'b0000000000011010;
    assign weights1[36][482] = 16'b0000000000001011;
    assign weights1[36][483] = 16'b0000000000001110;
    assign weights1[36][484] = 16'b0000000000010111;
    assign weights1[36][485] = 16'b0000000000010000;
    assign weights1[36][486] = 16'b0000000000010110;
    assign weights1[36][487] = 16'b0000000000011011;
    assign weights1[36][488] = 16'b0000000000000110;
    assign weights1[36][489] = 16'b0000000000010010;
    assign weights1[36][490] = 16'b1111111111100101;
    assign weights1[36][491] = 16'b1111111110010100;
    assign weights1[36][492] = 16'b1111111101110110;
    assign weights1[36][493] = 16'b1111111101101111;
    assign weights1[36][494] = 16'b1111111101111111;
    assign weights1[36][495] = 16'b1111111110011001;
    assign weights1[36][496] = 16'b1111111110100001;
    assign weights1[36][497] = 16'b1111111110101010;
    assign weights1[36][498] = 16'b1111111111000111;
    assign weights1[36][499] = 16'b1111111111001010;
    assign weights1[36][500] = 16'b1111111111001101;
    assign weights1[36][501] = 16'b1111111111010001;
    assign weights1[36][502] = 16'b1111111111100001;
    assign weights1[36][503] = 16'b1111111111100111;
    assign weights1[36][504] = 16'b1111111111111000;
    assign weights1[36][505] = 16'b0000000000010111;
    assign weights1[36][506] = 16'b0000000000100100;
    assign weights1[36][507] = 16'b0000000000001011;
    assign weights1[36][508] = 16'b0000000000000000;
    assign weights1[36][509] = 16'b0000000000010011;
    assign weights1[36][510] = 16'b0000000000000101;
    assign weights1[36][511] = 16'b1111111111111110;
    assign weights1[36][512] = 16'b0000000000000110;
    assign weights1[36][513] = 16'b0000000000001100;
    assign weights1[36][514] = 16'b0000000000001100;
    assign weights1[36][515] = 16'b0000000000011001;
    assign weights1[36][516] = 16'b0000000000010001;
    assign weights1[36][517] = 16'b0000000000011001;
    assign weights1[36][518] = 16'b1111111111101010;
    assign weights1[36][519] = 16'b1111111111001000;
    assign weights1[36][520] = 16'b1111111101110111;
    assign weights1[36][521] = 16'b1111111101001110;
    assign weights1[36][522] = 16'b1111111110000001;
    assign weights1[36][523] = 16'b1111111110011100;
    assign weights1[36][524] = 16'b1111111110101010;
    assign weights1[36][525] = 16'b1111111111001000;
    assign weights1[36][526] = 16'b1111111111000100;
    assign weights1[36][527] = 16'b1111111111010010;
    assign weights1[36][528] = 16'b1111111111010001;
    assign weights1[36][529] = 16'b1111111111011011;
    assign weights1[36][530] = 16'b1111111111100001;
    assign weights1[36][531] = 16'b1111111111101000;
    assign weights1[36][532] = 16'b1111111111111001;
    assign weights1[36][533] = 16'b0000000000000000;
    assign weights1[36][534] = 16'b0000000000000100;
    assign weights1[36][535] = 16'b0000000000000100;
    assign weights1[36][536] = 16'b1111111111111100;
    assign weights1[36][537] = 16'b1111111111111110;
    assign weights1[36][538] = 16'b0000000000001010;
    assign weights1[36][539] = 16'b0000000000010001;
    assign weights1[36][540] = 16'b0000000000010011;
    assign weights1[36][541] = 16'b0000000000000110;
    assign weights1[36][542] = 16'b0000000000010000;
    assign weights1[36][543] = 16'b0000000000001111;
    assign weights1[36][544] = 16'b0000000000010000;
    assign weights1[36][545] = 16'b0000000000100101;
    assign weights1[36][546] = 16'b0000000000100010;
    assign weights1[36][547] = 16'b0000000000001001;
    assign weights1[36][548] = 16'b1111111110101111;
    assign weights1[36][549] = 16'b1111111101110101;
    assign weights1[36][550] = 16'b1111111110000010;
    assign weights1[36][551] = 16'b1111111110011110;
    assign weights1[36][552] = 16'b1111111110110010;
    assign weights1[36][553] = 16'b1111111111000001;
    assign weights1[36][554] = 16'b1111111111001011;
    assign weights1[36][555] = 16'b1111111111010000;
    assign weights1[36][556] = 16'b1111111111010110;
    assign weights1[36][557] = 16'b1111111111011101;
    assign weights1[36][558] = 16'b1111111111100101;
    assign weights1[36][559] = 16'b1111111111101101;
    assign weights1[36][560] = 16'b1111111111111100;
    assign weights1[36][561] = 16'b0000000000000011;
    assign weights1[36][562] = 16'b1111111111111111;
    assign weights1[36][563] = 16'b0000000000011001;
    assign weights1[36][564] = 16'b0000000000010010;
    assign weights1[36][565] = 16'b0000000000001011;
    assign weights1[36][566] = 16'b1111111111110101;
    assign weights1[36][567] = 16'b0000000000011010;
    assign weights1[36][568] = 16'b0000000000000011;
    assign weights1[36][569] = 16'b0000000000001100;
    assign weights1[36][570] = 16'b0000000000001111;
    assign weights1[36][571] = 16'b0000000000001000;
    assign weights1[36][572] = 16'b0000000000100011;
    assign weights1[36][573] = 16'b0000000000011111;
    assign weights1[36][574] = 16'b0000000000101101;
    assign weights1[36][575] = 16'b0000000000101110;
    assign weights1[36][576] = 16'b1111111111110100;
    assign weights1[36][577] = 16'b1111111110011101;
    assign weights1[36][578] = 16'b1111111110001011;
    assign weights1[36][579] = 16'b1111111110011100;
    assign weights1[36][580] = 16'b1111111110111001;
    assign weights1[36][581] = 16'b1111111111001000;
    assign weights1[36][582] = 16'b1111111111010100;
    assign weights1[36][583] = 16'b1111111111011010;
    assign weights1[36][584] = 16'b1111111111011101;
    assign weights1[36][585] = 16'b1111111111011111;
    assign weights1[36][586] = 16'b1111111111100110;
    assign weights1[36][587] = 16'b1111111111101011;
    assign weights1[36][588] = 16'b1111111111110111;
    assign weights1[36][589] = 16'b0000000000001101;
    assign weights1[36][590] = 16'b0000000000010100;
    assign weights1[36][591] = 16'b0000000000001100;
    assign weights1[36][592] = 16'b1111111111110101;
    assign weights1[36][593] = 16'b0000000000011101;
    assign weights1[36][594] = 16'b0000000000001101;
    assign weights1[36][595] = 16'b0000000000011101;
    assign weights1[36][596] = 16'b0000000000001111;
    assign weights1[36][597] = 16'b0000000000010000;
    assign weights1[36][598] = 16'b0000000000001101;
    assign weights1[36][599] = 16'b0000000000001001;
    assign weights1[36][600] = 16'b0000000000010001;
    assign weights1[36][601] = 16'b0000000000011010;
    assign weights1[36][602] = 16'b0000000000010001;
    assign weights1[36][603] = 16'b0000000000111000;
    assign weights1[36][604] = 16'b0000000000000100;
    assign weights1[36][605] = 16'b1111111110111000;
    assign weights1[36][606] = 16'b1111111110011010;
    assign weights1[36][607] = 16'b1111111110100010;
    assign weights1[36][608] = 16'b1111111110111110;
    assign weights1[36][609] = 16'b1111111111001111;
    assign weights1[36][610] = 16'b1111111111010111;
    assign weights1[36][611] = 16'b1111111111011010;
    assign weights1[36][612] = 16'b1111111111100001;
    assign weights1[36][613] = 16'b1111111111100011;
    assign weights1[36][614] = 16'b1111111111101110;
    assign weights1[36][615] = 16'b1111111111100110;
    assign weights1[36][616] = 16'b1111111111111001;
    assign weights1[36][617] = 16'b0000000000000101;
    assign weights1[36][618] = 16'b0000000000010011;
    assign weights1[36][619] = 16'b0000000000010001;
    assign weights1[36][620] = 16'b0000000000001000;
    assign weights1[36][621] = 16'b0000000000000100;
    assign weights1[36][622] = 16'b0000000000010100;
    assign weights1[36][623] = 16'b0000000000001101;
    assign weights1[36][624] = 16'b1111111111110100;
    assign weights1[36][625] = 16'b0000000000001001;
    assign weights1[36][626] = 16'b0000000000000101;
    assign weights1[36][627] = 16'b0000000000000111;
    assign weights1[36][628] = 16'b0000000000011001;
    assign weights1[36][629] = 16'b0000000000000010;
    assign weights1[36][630] = 16'b0000000000010111;
    assign weights1[36][631] = 16'b0000000000100101;
    assign weights1[36][632] = 16'b0000000000101010;
    assign weights1[36][633] = 16'b1111111111010111;
    assign weights1[36][634] = 16'b1111111110111000;
    assign weights1[36][635] = 16'b1111111110101101;
    assign weights1[36][636] = 16'b1111111111001010;
    assign weights1[36][637] = 16'b1111111111010000;
    assign weights1[36][638] = 16'b1111111111011010;
    assign weights1[36][639] = 16'b1111111111011110;
    assign weights1[36][640] = 16'b1111111111100100;
    assign weights1[36][641] = 16'b1111111111100101;
    assign weights1[36][642] = 16'b1111111111100110;
    assign weights1[36][643] = 16'b1111111111101101;
    assign weights1[36][644] = 16'b1111111111111101;
    assign weights1[36][645] = 16'b0000000000010000;
    assign weights1[36][646] = 16'b0000000000001100;
    assign weights1[36][647] = 16'b0000000000001011;
    assign weights1[36][648] = 16'b0000000000010001;
    assign weights1[36][649] = 16'b0000000000010111;
    assign weights1[36][650] = 16'b1111111111111101;
    assign weights1[36][651] = 16'b0000000000001001;
    assign weights1[36][652] = 16'b1111111111111010;
    assign weights1[36][653] = 16'b0000000000010110;
    assign weights1[36][654] = 16'b0000000000010110;
    assign weights1[36][655] = 16'b0000000000010000;
    assign weights1[36][656] = 16'b0000000000000011;
    assign weights1[36][657] = 16'b0000000000000111;
    assign weights1[36][658] = 16'b0000000000011110;
    assign weights1[36][659] = 16'b0000000000010100;
    assign weights1[36][660] = 16'b0000000000101001;
    assign weights1[36][661] = 16'b1111111111011000;
    assign weights1[36][662] = 16'b1111111110111001;
    assign weights1[36][663] = 16'b1111111110111001;
    assign weights1[36][664] = 16'b1111111111001100;
    assign weights1[36][665] = 16'b1111111111001111;
    assign weights1[36][666] = 16'b1111111111011011;
    assign weights1[36][667] = 16'b1111111111100000;
    assign weights1[36][668] = 16'b1111111111100001;
    assign weights1[36][669] = 16'b1111111111100101;
    assign weights1[36][670] = 16'b1111111111101011;
    assign weights1[36][671] = 16'b1111111111110000;
    assign weights1[36][672] = 16'b1111111111111000;
    assign weights1[36][673] = 16'b0000000000000101;
    assign weights1[36][674] = 16'b0000000000010001;
    assign weights1[36][675] = 16'b0000000000010100;
    assign weights1[36][676] = 16'b0000000000010101;
    assign weights1[36][677] = 16'b0000000000011011;
    assign weights1[36][678] = 16'b0000000000001000;
    assign weights1[36][679] = 16'b0000000000010100;
    assign weights1[36][680] = 16'b0000000000000101;
    assign weights1[36][681] = 16'b0000000000001001;
    assign weights1[36][682] = 16'b0000000000011101;
    assign weights1[36][683] = 16'b0000000000010111;
    assign weights1[36][684] = 16'b0000000000010110;
    assign weights1[36][685] = 16'b0000000000010110;
    assign weights1[36][686] = 16'b0000000000100000;
    assign weights1[36][687] = 16'b0000000000111101;
    assign weights1[36][688] = 16'b0000000000011111;
    assign weights1[36][689] = 16'b1111111111110110;
    assign weights1[36][690] = 16'b1111111111010001;
    assign weights1[36][691] = 16'b1111111111001000;
    assign weights1[36][692] = 16'b1111111111010010;
    assign weights1[36][693] = 16'b1111111111100000;
    assign weights1[36][694] = 16'b1111111111100101;
    assign weights1[36][695] = 16'b1111111111100011;
    assign weights1[36][696] = 16'b1111111111100100;
    assign weights1[36][697] = 16'b1111111111101010;
    assign weights1[36][698] = 16'b1111111111110000;
    assign weights1[36][699] = 16'b1111111111111001;
    assign weights1[36][700] = 16'b0000000000000011;
    assign weights1[36][701] = 16'b0000000000001001;
    assign weights1[36][702] = 16'b0000000000001001;
    assign weights1[36][703] = 16'b0000000000001100;
    assign weights1[36][704] = 16'b0000000000000111;
    assign weights1[36][705] = 16'b0000000000010001;
    assign weights1[36][706] = 16'b0000000000000000;
    assign weights1[36][707] = 16'b0000000000001010;
    assign weights1[36][708] = 16'b0000000000010000;
    assign weights1[36][709] = 16'b1111111111111101;
    assign weights1[36][710] = 16'b0000000000011110;
    assign weights1[36][711] = 16'b0000000000010001;
    assign weights1[36][712] = 16'b0000000000001101;
    assign weights1[36][713] = 16'b0000000000010000;
    assign weights1[36][714] = 16'b0000000000010000;
    assign weights1[36][715] = 16'b0000000000001010;
    assign weights1[36][716] = 16'b0000000000000001;
    assign weights1[36][717] = 16'b1111111111100011;
    assign weights1[36][718] = 16'b1111111111001100;
    assign weights1[36][719] = 16'b1111111111001010;
    assign weights1[36][720] = 16'b1111111111011010;
    assign weights1[36][721] = 16'b1111111111100011;
    assign weights1[36][722] = 16'b1111111111100000;
    assign weights1[36][723] = 16'b1111111111011111;
    assign weights1[36][724] = 16'b1111111111101101;
    assign weights1[36][725] = 16'b1111111111110101;
    assign weights1[36][726] = 16'b1111111111111010;
    assign weights1[36][727] = 16'b1111111111111111;
    assign weights1[36][728] = 16'b0000000000000010;
    assign weights1[36][729] = 16'b0000000000001000;
    assign weights1[36][730] = 16'b0000000000010010;
    assign weights1[36][731] = 16'b0000000000001011;
    assign weights1[36][732] = 16'b1111111111111101;
    assign weights1[36][733] = 16'b0000000000010000;
    assign weights1[36][734] = 16'b0000000000000101;
    assign weights1[36][735] = 16'b0000000000001111;
    assign weights1[36][736] = 16'b0000000000011000;
    assign weights1[36][737] = 16'b0000000000010000;
    assign weights1[36][738] = 16'b0000000000011111;
    assign weights1[36][739] = 16'b0000000000000101;
    assign weights1[36][740] = 16'b0000000000010110;
    assign weights1[36][741] = 16'b0000000000011011;
    assign weights1[36][742] = 16'b0000000000001111;
    assign weights1[36][743] = 16'b0000000000010001;
    assign weights1[36][744] = 16'b1111111111111111;
    assign weights1[36][745] = 16'b1111111111011110;
    assign weights1[36][746] = 16'b1111111111100000;
    assign weights1[36][747] = 16'b1111111111010010;
    assign weights1[36][748] = 16'b1111111111011100;
    assign weights1[36][749] = 16'b1111111111011111;
    assign weights1[36][750] = 16'b1111111111100101;
    assign weights1[36][751] = 16'b1111111111101101;
    assign weights1[36][752] = 16'b1111111111110011;
    assign weights1[36][753] = 16'b1111111111111000;
    assign weights1[36][754] = 16'b1111111111111101;
    assign weights1[36][755] = 16'b0000000000000000;
    assign weights1[36][756] = 16'b0000000000000010;
    assign weights1[36][757] = 16'b0000000000000000;
    assign weights1[36][758] = 16'b0000000000000111;
    assign weights1[36][759] = 16'b0000000000001010;
    assign weights1[36][760] = 16'b0000000000001110;
    assign weights1[36][761] = 16'b0000000000001111;
    assign weights1[36][762] = 16'b0000000000011001;
    assign weights1[36][763] = 16'b0000000000011010;
    assign weights1[36][764] = 16'b0000000000010110;
    assign weights1[36][765] = 16'b0000000000011001;
    assign weights1[36][766] = 16'b0000000000011011;
    assign weights1[36][767] = 16'b0000000000100100;
    assign weights1[36][768] = 16'b0000000000100001;
    assign weights1[36][769] = 16'b0000000000010111;
    assign weights1[36][770] = 16'b0000000000000011;
    assign weights1[36][771] = 16'b1111111111111100;
    assign weights1[36][772] = 16'b1111111111110001;
    assign weights1[36][773] = 16'b1111111111100101;
    assign weights1[36][774] = 16'b1111111111100000;
    assign weights1[36][775] = 16'b1111111111011111;
    assign weights1[36][776] = 16'b1111111111100100;
    assign weights1[36][777] = 16'b1111111111100111;
    assign weights1[36][778] = 16'b1111111111101111;
    assign weights1[36][779] = 16'b1111111111110111;
    assign weights1[36][780] = 16'b1111111111111001;
    assign weights1[36][781] = 16'b1111111111111110;
    assign weights1[36][782] = 16'b0000000000000000;
    assign weights1[36][783] = 16'b0000000000000000;
    assign weights1[37][0] = 16'b0000000000000000;
    assign weights1[37][1] = 16'b0000000000000001;
    assign weights1[37][2] = 16'b0000000000000001;
    assign weights1[37][3] = 16'b1111111111111110;
    assign weights1[37][4] = 16'b1111111111111010;
    assign weights1[37][5] = 16'b1111111111111011;
    assign weights1[37][6] = 16'b1111111111111100;
    assign weights1[37][7] = 16'b1111111111111110;
    assign weights1[37][8] = 16'b1111111111111111;
    assign weights1[37][9] = 16'b1111111111110001;
    assign weights1[37][10] = 16'b1111111111101110;
    assign weights1[37][11] = 16'b1111111111110111;
    assign weights1[37][12] = 16'b1111111111110110;
    assign weights1[37][13] = 16'b0000000000000100;
    assign weights1[37][14] = 16'b0000000000000011;
    assign weights1[37][15] = 16'b0000000000000101;
    assign weights1[37][16] = 16'b1111111111111111;
    assign weights1[37][17] = 16'b1111111111110000;
    assign weights1[37][18] = 16'b1111111111111010;
    assign weights1[37][19] = 16'b1111111111111100;
    assign weights1[37][20] = 16'b0000000000000000;
    assign weights1[37][21] = 16'b1111111111111101;
    assign weights1[37][22] = 16'b1111111111111000;
    assign weights1[37][23] = 16'b1111111111110101;
    assign weights1[37][24] = 16'b1111111111111110;
    assign weights1[37][25] = 16'b0000000000000111;
    assign weights1[37][26] = 16'b0000000000000010;
    assign weights1[37][27] = 16'b1111111111111110;
    assign weights1[37][28] = 16'b1111111111111111;
    assign weights1[37][29] = 16'b0000000000000001;
    assign weights1[37][30] = 16'b0000000000000000;
    assign weights1[37][31] = 16'b1111111111111111;
    assign weights1[37][32] = 16'b1111111111111101;
    assign weights1[37][33] = 16'b1111111111110111;
    assign weights1[37][34] = 16'b1111111111111001;
    assign weights1[37][35] = 16'b1111111111111111;
    assign weights1[37][36] = 16'b1111111111111111;
    assign weights1[37][37] = 16'b1111111111110011;
    assign weights1[37][38] = 16'b1111111111111011;
    assign weights1[37][39] = 16'b1111111111110010;
    assign weights1[37][40] = 16'b0000000000000001;
    assign weights1[37][41] = 16'b0000000000000110;
    assign weights1[37][42] = 16'b0000000000000100;
    assign weights1[37][43] = 16'b1111111111111001;
    assign weights1[37][44] = 16'b1111111111111110;
    assign weights1[37][45] = 16'b1111111111111000;
    assign weights1[37][46] = 16'b1111111111110101;
    assign weights1[37][47] = 16'b0000000000000010;
    assign weights1[37][48] = 16'b0000000000000110;
    assign weights1[37][49] = 16'b0000000000000101;
    assign weights1[37][50] = 16'b1111111111110101;
    assign weights1[37][51] = 16'b1111111111110111;
    assign weights1[37][52] = 16'b0000000000000010;
    assign weights1[37][53] = 16'b0000000000001001;
    assign weights1[37][54] = 16'b0000000000000000;
    assign weights1[37][55] = 16'b0000000000000001;
    assign weights1[37][56] = 16'b0000000000000000;
    assign weights1[37][57] = 16'b1111111111111101;
    assign weights1[37][58] = 16'b1111111111111110;
    assign weights1[37][59] = 16'b0000000000000111;
    assign weights1[37][60] = 16'b1111111111111001;
    assign weights1[37][61] = 16'b0000000000000000;
    assign weights1[37][62] = 16'b1111111111101100;
    assign weights1[37][63] = 16'b1111111111110010;
    assign weights1[37][64] = 16'b1111111111111111;
    assign weights1[37][65] = 16'b0000000000001000;
    assign weights1[37][66] = 16'b1111111111111110;
    assign weights1[37][67] = 16'b0000000000000010;
    assign weights1[37][68] = 16'b1111111111110101;
    assign weights1[37][69] = 16'b0000000000000110;
    assign weights1[37][70] = 16'b1111111111110110;
    assign weights1[37][71] = 16'b0000000000001001;
    assign weights1[37][72] = 16'b0000000000000000;
    assign weights1[37][73] = 16'b1111111111111000;
    assign weights1[37][74] = 16'b1111111111111101;
    assign weights1[37][75] = 16'b1111111111110101;
    assign weights1[37][76] = 16'b0000000000000100;
    assign weights1[37][77] = 16'b1111111111110101;
    assign weights1[37][78] = 16'b1111111111101110;
    assign weights1[37][79] = 16'b0000000000000010;
    assign weights1[37][80] = 16'b0000000000000001;
    assign weights1[37][81] = 16'b0000000000000001;
    assign weights1[37][82] = 16'b0000000000001001;
    assign weights1[37][83] = 16'b1111111111111110;
    assign weights1[37][84] = 16'b1111111111111111;
    assign weights1[37][85] = 16'b1111111111111100;
    assign weights1[37][86] = 16'b0000000000000000;
    assign weights1[37][87] = 16'b0000000000000000;
    assign weights1[37][88] = 16'b1111111111110110;
    assign weights1[37][89] = 16'b1111111111111010;
    assign weights1[37][90] = 16'b1111111111111110;
    assign weights1[37][91] = 16'b1111111111111000;
    assign weights1[37][92] = 16'b1111111111111100;
    assign weights1[37][93] = 16'b0000000000000000;
    assign weights1[37][94] = 16'b0000000000001111;
    assign weights1[37][95] = 16'b1111111111111101;
    assign weights1[37][96] = 16'b0000000000000110;
    assign weights1[37][97] = 16'b1111111111110110;
    assign weights1[37][98] = 16'b0000000000000111;
    assign weights1[37][99] = 16'b0000000000000111;
    assign weights1[37][100] = 16'b1111111111110011;
    assign weights1[37][101] = 16'b0000000000000100;
    assign weights1[37][102] = 16'b1111111111111101;
    assign weights1[37][103] = 16'b0000000000001001;
    assign weights1[37][104] = 16'b1111111111111011;
    assign weights1[37][105] = 16'b1111111111111100;
    assign weights1[37][106] = 16'b0000000000000010;
    assign weights1[37][107] = 16'b0000000000001000;
    assign weights1[37][108] = 16'b0000000000000111;
    assign weights1[37][109] = 16'b1111111111111010;
    assign weights1[37][110] = 16'b0000000000000001;
    assign weights1[37][111] = 16'b1111111111111110;
    assign weights1[37][112] = 16'b1111111111111110;
    assign weights1[37][113] = 16'b1111111111111011;
    assign weights1[37][114] = 16'b1111111111111110;
    assign weights1[37][115] = 16'b1111111111111110;
    assign weights1[37][116] = 16'b0000000000000011;
    assign weights1[37][117] = 16'b0000000000000001;
    assign weights1[37][118] = 16'b0000000000000101;
    assign weights1[37][119] = 16'b1111111111111011;
    assign weights1[37][120] = 16'b0000000000000100;
    assign weights1[37][121] = 16'b1111111111111110;
    assign weights1[37][122] = 16'b1111111111111101;
    assign weights1[37][123] = 16'b1111111111111101;
    assign weights1[37][124] = 16'b0000000000000100;
    assign weights1[37][125] = 16'b0000000000000011;
    assign weights1[37][126] = 16'b0000000000001000;
    assign weights1[37][127] = 16'b0000000000000110;
    assign weights1[37][128] = 16'b0000000000001011;
    assign weights1[37][129] = 16'b1111111111101101;
    assign weights1[37][130] = 16'b0000000000000010;
    assign weights1[37][131] = 16'b0000000000000000;
    assign weights1[37][132] = 16'b0000000000001110;
    assign weights1[37][133] = 16'b0000000000000011;
    assign weights1[37][134] = 16'b1111111111110011;
    assign weights1[37][135] = 16'b1111111111111101;
    assign weights1[37][136] = 16'b1111111111110110;
    assign weights1[37][137] = 16'b1111111111111110;
    assign weights1[37][138] = 16'b1111111111111100;
    assign weights1[37][139] = 16'b1111111111110100;
    assign weights1[37][140] = 16'b0000000000000010;
    assign weights1[37][141] = 16'b0000000000000000;
    assign weights1[37][142] = 16'b1111111111111101;
    assign weights1[37][143] = 16'b1111111111110101;
    assign weights1[37][144] = 16'b1111111111111001;
    assign weights1[37][145] = 16'b0000000000000000;
    assign weights1[37][146] = 16'b0000000000000000;
    assign weights1[37][147] = 16'b1111111111110011;
    assign weights1[37][148] = 16'b1111111111111010;
    assign weights1[37][149] = 16'b1111111111111110;
    assign weights1[37][150] = 16'b1111111111111100;
    assign weights1[37][151] = 16'b1111111111111111;
    assign weights1[37][152] = 16'b1111111111110000;
    assign weights1[37][153] = 16'b1111111111110010;
    assign weights1[37][154] = 16'b0000000000001011;
    assign weights1[37][155] = 16'b0000000000000100;
    assign weights1[37][156] = 16'b1111111111111111;
    assign weights1[37][157] = 16'b1111111111111010;
    assign weights1[37][158] = 16'b1111111111110110;
    assign weights1[37][159] = 16'b0000000000001001;
    assign weights1[37][160] = 16'b1111111111110100;
    assign weights1[37][161] = 16'b0000000000011010;
    assign weights1[37][162] = 16'b0000000000000001;
    assign weights1[37][163] = 16'b0000000000001011;
    assign weights1[37][164] = 16'b0000000000000100;
    assign weights1[37][165] = 16'b0000000000000010;
    assign weights1[37][166] = 16'b1111111111111111;
    assign weights1[37][167] = 16'b0000000000000100;
    assign weights1[37][168] = 16'b0000000000000111;
    assign weights1[37][169] = 16'b0000000000000010;
    assign weights1[37][170] = 16'b0000000000001011;
    assign weights1[37][171] = 16'b0000000000000011;
    assign weights1[37][172] = 16'b0000000000000101;
    assign weights1[37][173] = 16'b1111111111111010;
    assign weights1[37][174] = 16'b1111111111110010;
    assign weights1[37][175] = 16'b1111111111111101;
    assign weights1[37][176] = 16'b1111111111111101;
    assign weights1[37][177] = 16'b1111111111111100;
    assign weights1[37][178] = 16'b0000000000000000;
    assign weights1[37][179] = 16'b1111111111111000;
    assign weights1[37][180] = 16'b0000000000000101;
    assign weights1[37][181] = 16'b1111111111110011;
    assign weights1[37][182] = 16'b1111111111101111;
    assign weights1[37][183] = 16'b1111111111111101;
    assign weights1[37][184] = 16'b1111111111111110;
    assign weights1[37][185] = 16'b0000000000000100;
    assign weights1[37][186] = 16'b1111111111111011;
    assign weights1[37][187] = 16'b1111111111110111;
    assign weights1[37][188] = 16'b1111111111111000;
    assign weights1[37][189] = 16'b0000000000001011;
    assign weights1[37][190] = 16'b0000000000000011;
    assign weights1[37][191] = 16'b1111111111111110;
    assign weights1[37][192] = 16'b1111111111101110;
    assign weights1[37][193] = 16'b1111111111111011;
    assign weights1[37][194] = 16'b1111111111111111;
    assign weights1[37][195] = 16'b0000000000000110;
    assign weights1[37][196] = 16'b0000000000001011;
    assign weights1[37][197] = 16'b0000000000010001;
    assign weights1[37][198] = 16'b0000000000001100;
    assign weights1[37][199] = 16'b0000000000000011;
    assign weights1[37][200] = 16'b0000000000000101;
    assign weights1[37][201] = 16'b1111111111110101;
    assign weights1[37][202] = 16'b0000000000001110;
    assign weights1[37][203] = 16'b1111111111111100;
    assign weights1[37][204] = 16'b1111111111111100;
    assign weights1[37][205] = 16'b0000000000000000;
    assign weights1[37][206] = 16'b1111111111101000;
    assign weights1[37][207] = 16'b0000000000000010;
    assign weights1[37][208] = 16'b0000000000000011;
    assign weights1[37][209] = 16'b0000000000000010;
    assign weights1[37][210] = 16'b0000000000010100;
    assign weights1[37][211] = 16'b1111111111110000;
    assign weights1[37][212] = 16'b0000000000000100;
    assign weights1[37][213] = 16'b0000000000000111;
    assign weights1[37][214] = 16'b0000000000000010;
    assign weights1[37][215] = 16'b0000000000000011;
    assign weights1[37][216] = 16'b0000000000000011;
    assign weights1[37][217] = 16'b1111111111111100;
    assign weights1[37][218] = 16'b0000000000000101;
    assign weights1[37][219] = 16'b0000000000000001;
    assign weights1[37][220] = 16'b1111111111111011;
    assign weights1[37][221] = 16'b0000000000000001;
    assign weights1[37][222] = 16'b0000000000001001;
    assign weights1[37][223] = 16'b0000000000001001;
    assign weights1[37][224] = 16'b0000000000001100;
    assign weights1[37][225] = 16'b0000000000010110;
    assign weights1[37][226] = 16'b0000000000000000;
    assign weights1[37][227] = 16'b0000000000010001;
    assign weights1[37][228] = 16'b1111111111111010;
    assign weights1[37][229] = 16'b1111111111111110;
    assign weights1[37][230] = 16'b0000000000000000;
    assign weights1[37][231] = 16'b0000000000000001;
    assign weights1[37][232] = 16'b1111111111110101;
    assign weights1[37][233] = 16'b1111111111110111;
    assign weights1[37][234] = 16'b1111111111111101;
    assign weights1[37][235] = 16'b1111111111110011;
    assign weights1[37][236] = 16'b0000000000001000;
    assign weights1[37][237] = 16'b1111111111111001;
    assign weights1[37][238] = 16'b1111111111111010;
    assign weights1[37][239] = 16'b1111111111111100;
    assign weights1[37][240] = 16'b0000000000000000;
    assign weights1[37][241] = 16'b1111111111111001;
    assign weights1[37][242] = 16'b0000000000001101;
    assign weights1[37][243] = 16'b0000000000001111;
    assign weights1[37][244] = 16'b0000000000001000;
    assign weights1[37][245] = 16'b1111111111110111;
    assign weights1[37][246] = 16'b1111111111111000;
    assign weights1[37][247] = 16'b1111111111111110;
    assign weights1[37][248] = 16'b0000000000000101;
    assign weights1[37][249] = 16'b0000000000010001;
    assign weights1[37][250] = 16'b1111111111101111;
    assign weights1[37][251] = 16'b1111111111110111;
    assign weights1[37][252] = 16'b0000000000001110;
    assign weights1[37][253] = 16'b0000000000001101;
    assign weights1[37][254] = 16'b1111111111111000;
    assign weights1[37][255] = 16'b0000000000000000;
    assign weights1[37][256] = 16'b1111111111111010;
    assign weights1[37][257] = 16'b1111111111111011;
    assign weights1[37][258] = 16'b0000000000000100;
    assign weights1[37][259] = 16'b0000000000000010;
    assign weights1[37][260] = 16'b0000000000001100;
    assign weights1[37][261] = 16'b0000000000001000;
    assign weights1[37][262] = 16'b1111111111110000;
    assign weights1[37][263] = 16'b1111111111111001;
    assign weights1[37][264] = 16'b1111111111110101;
    assign weights1[37][265] = 16'b1111111111111000;
    assign weights1[37][266] = 16'b0000000000001111;
    assign weights1[37][267] = 16'b1111111111111010;
    assign weights1[37][268] = 16'b1111111111111000;
    assign weights1[37][269] = 16'b0000000000001011;
    assign weights1[37][270] = 16'b1111111111111010;
    assign weights1[37][271] = 16'b0000000000000000;
    assign weights1[37][272] = 16'b1111111111110110;
    assign weights1[37][273] = 16'b0000000000001001;
    assign weights1[37][274] = 16'b0000000000001010;
    assign weights1[37][275] = 16'b1111111111111110;
    assign weights1[37][276] = 16'b1111111111111110;
    assign weights1[37][277] = 16'b1111111111111001;
    assign weights1[37][278] = 16'b0000000000000100;
    assign weights1[37][279] = 16'b0000000000000000;
    assign weights1[37][280] = 16'b0000000000000110;
    assign weights1[37][281] = 16'b1111111111111100;
    assign weights1[37][282] = 16'b1111111111110011;
    assign weights1[37][283] = 16'b0000000000000011;
    assign weights1[37][284] = 16'b1111111111111000;
    assign weights1[37][285] = 16'b1111111111111001;
    assign weights1[37][286] = 16'b1111111111110001;
    assign weights1[37][287] = 16'b0000000000000000;
    assign weights1[37][288] = 16'b1111111111111000;
    assign weights1[37][289] = 16'b1111111111111111;
    assign weights1[37][290] = 16'b0000000000001011;
    assign weights1[37][291] = 16'b1111111111110001;
    assign weights1[37][292] = 16'b0000000000001101;
    assign weights1[37][293] = 16'b1111111111101101;
    assign weights1[37][294] = 16'b1111111111110111;
    assign weights1[37][295] = 16'b1111111111111000;
    assign weights1[37][296] = 16'b1111111111111110;
    assign weights1[37][297] = 16'b1111111111111011;
    assign weights1[37][298] = 16'b0000000000000110;
    assign weights1[37][299] = 16'b0000000000000101;
    assign weights1[37][300] = 16'b0000000000000111;
    assign weights1[37][301] = 16'b0000000000000001;
    assign weights1[37][302] = 16'b1111111111110011;
    assign weights1[37][303] = 16'b0000000000001111;
    assign weights1[37][304] = 16'b1111111111111111;
    assign weights1[37][305] = 16'b0000000000010100;
    assign weights1[37][306] = 16'b1111111111110100;
    assign weights1[37][307] = 16'b1111111111111011;
    assign weights1[37][308] = 16'b0000000000000111;
    assign weights1[37][309] = 16'b0000000000000111;
    assign weights1[37][310] = 16'b1111111111111110;
    assign weights1[37][311] = 16'b0000000000010011;
    assign weights1[37][312] = 16'b0000000000011011;
    assign weights1[37][313] = 16'b1111111111111111;
    assign weights1[37][314] = 16'b0000000000001001;
    assign weights1[37][315] = 16'b0000000000000111;
    assign weights1[37][316] = 16'b0000000000000011;
    assign weights1[37][317] = 16'b0000000000000101;
    assign weights1[37][318] = 16'b0000000000001000;
    assign weights1[37][319] = 16'b1111111111110110;
    assign weights1[37][320] = 16'b0000000000000111;
    assign weights1[37][321] = 16'b1111111111111101;
    assign weights1[37][322] = 16'b0000000000000101;
    assign weights1[37][323] = 16'b1111111111111110;
    assign weights1[37][324] = 16'b1111111111111101;
    assign weights1[37][325] = 16'b0000000000000001;
    assign weights1[37][326] = 16'b0000000000000000;
    assign weights1[37][327] = 16'b0000000000000111;
    assign weights1[37][328] = 16'b1111111111111010;
    assign weights1[37][329] = 16'b0000000000000111;
    assign weights1[37][330] = 16'b0000000000001000;
    assign weights1[37][331] = 16'b1111111111111001;
    assign weights1[37][332] = 16'b0000000000000001;
    assign weights1[37][333] = 16'b1111111111110000;
    assign weights1[37][334] = 16'b1111111111111000;
    assign weights1[37][335] = 16'b0000000000000100;
    assign weights1[37][336] = 16'b0000000000001000;
    assign weights1[37][337] = 16'b1111111111110111;
    assign weights1[37][338] = 16'b0000000000000010;
    assign weights1[37][339] = 16'b0000000000001100;
    assign weights1[37][340] = 16'b1111111111111101;
    assign weights1[37][341] = 16'b0000000000001011;
    assign weights1[37][342] = 16'b0000000000000101;
    assign weights1[37][343] = 16'b0000000000001011;
    assign weights1[37][344] = 16'b0000000000001011;
    assign weights1[37][345] = 16'b1111111111111011;
    assign weights1[37][346] = 16'b1111111111110101;
    assign weights1[37][347] = 16'b0000000000001010;
    assign weights1[37][348] = 16'b1111111111110101;
    assign weights1[37][349] = 16'b0000000000000111;
    assign weights1[37][350] = 16'b1111111111110000;
    assign weights1[37][351] = 16'b0000000000000100;
    assign weights1[37][352] = 16'b1111111111111111;
    assign weights1[37][353] = 16'b0000000000000110;
    assign weights1[37][354] = 16'b0000000000000000;
    assign weights1[37][355] = 16'b1111111111110110;
    assign weights1[37][356] = 16'b0000000000001110;
    assign weights1[37][357] = 16'b0000000000000110;
    assign weights1[37][358] = 16'b0000000000000000;
    assign weights1[37][359] = 16'b0000000000000011;
    assign weights1[37][360] = 16'b1111111111101110;
    assign weights1[37][361] = 16'b1111111111111100;
    assign weights1[37][362] = 16'b1111111111110110;
    assign weights1[37][363] = 16'b1111111111111110;
    assign weights1[37][364] = 16'b1111111111111101;
    assign weights1[37][365] = 16'b1111111111111000;
    assign weights1[37][366] = 16'b0000000000001010;
    assign weights1[37][367] = 16'b0000000000000011;
    assign weights1[37][368] = 16'b1111111111110101;
    assign weights1[37][369] = 16'b1111111111111001;
    assign weights1[37][370] = 16'b0000000000000011;
    assign weights1[37][371] = 16'b0000000000000000;
    assign weights1[37][372] = 16'b1111111111110111;
    assign weights1[37][373] = 16'b0000000000001101;
    assign weights1[37][374] = 16'b0000000000001001;
    assign weights1[37][375] = 16'b0000000000001001;
    assign weights1[37][376] = 16'b1111111111110010;
    assign weights1[37][377] = 16'b1111111111111010;
    assign weights1[37][378] = 16'b0000000000000011;
    assign weights1[37][379] = 16'b1111111111101101;
    assign weights1[37][380] = 16'b1111111111111110;
    assign weights1[37][381] = 16'b0000000000000100;
    assign weights1[37][382] = 16'b1111111111111111;
    assign weights1[37][383] = 16'b0000000000000110;
    assign weights1[37][384] = 16'b0000000000010010;
    assign weights1[37][385] = 16'b1111111111111001;
    assign weights1[37][386] = 16'b1111111111111010;
    assign weights1[37][387] = 16'b1111111111110100;
    assign weights1[37][388] = 16'b0000000000001001;
    assign weights1[37][389] = 16'b1111111111111000;
    assign weights1[37][390] = 16'b0000000000000100;
    assign weights1[37][391] = 16'b1111111111111100;
    assign weights1[37][392] = 16'b1111111111110100;
    assign weights1[37][393] = 16'b1111111111101111;
    assign weights1[37][394] = 16'b1111111111111110;
    assign weights1[37][395] = 16'b1111111111101110;
    assign weights1[37][396] = 16'b1111111111110101;
    assign weights1[37][397] = 16'b0000000000001000;
    assign weights1[37][398] = 16'b1111111111111000;
    assign weights1[37][399] = 16'b0000000000001000;
    assign weights1[37][400] = 16'b0000000000001000;
    assign weights1[37][401] = 16'b1111111111111110;
    assign weights1[37][402] = 16'b1111111111111100;
    assign weights1[37][403] = 16'b0000000000000010;
    assign weights1[37][404] = 16'b0000000000001011;
    assign weights1[37][405] = 16'b0000000000000000;
    assign weights1[37][406] = 16'b0000000000000001;
    assign weights1[37][407] = 16'b1111111111110100;
    assign weights1[37][408] = 16'b0000000000000011;
    assign weights1[37][409] = 16'b1111111111111010;
    assign weights1[37][410] = 16'b0000000000010001;
    assign weights1[37][411] = 16'b0000000000000001;
    assign weights1[37][412] = 16'b0000000000001000;
    assign weights1[37][413] = 16'b1111111111111110;
    assign weights1[37][414] = 16'b0000000000001100;
    assign weights1[37][415] = 16'b0000000000001000;
    assign weights1[37][416] = 16'b1111111111111011;
    assign weights1[37][417] = 16'b0000000000000001;
    assign weights1[37][418] = 16'b0000000000000110;
    assign weights1[37][419] = 16'b0000000000000110;
    assign weights1[37][420] = 16'b1111111111110011;
    assign weights1[37][421] = 16'b1111111111110101;
    assign weights1[37][422] = 16'b1111111111111000;
    assign weights1[37][423] = 16'b1111111111110110;
    assign weights1[37][424] = 16'b0000000000000101;
    assign weights1[37][425] = 16'b0000000000001010;
    assign weights1[37][426] = 16'b0000000000000011;
    assign weights1[37][427] = 16'b0000000000011001;
    assign weights1[37][428] = 16'b0000000000001011;
    assign weights1[37][429] = 16'b0000000000001110;
    assign weights1[37][430] = 16'b1111111111101110;
    assign weights1[37][431] = 16'b0000000000001010;
    assign weights1[37][432] = 16'b1111111111110100;
    assign weights1[37][433] = 16'b1111111111111001;
    assign weights1[37][434] = 16'b0000000000000011;
    assign weights1[37][435] = 16'b0000000000000010;
    assign weights1[37][436] = 16'b1111111111110000;
    assign weights1[37][437] = 16'b0000000000000000;
    assign weights1[37][438] = 16'b0000000000000010;
    assign weights1[37][439] = 16'b0000000000000111;
    assign weights1[37][440] = 16'b0000000000010000;
    assign weights1[37][441] = 16'b0000000000000100;
    assign weights1[37][442] = 16'b0000000000001001;
    assign weights1[37][443] = 16'b1111111111110001;
    assign weights1[37][444] = 16'b1111111111111110;
    assign weights1[37][445] = 16'b0000000000001000;
    assign weights1[37][446] = 16'b0000000000000000;
    assign weights1[37][447] = 16'b0000000000000101;
    assign weights1[37][448] = 16'b1111111111110011;
    assign weights1[37][449] = 16'b1111111111110110;
    assign weights1[37][450] = 16'b0000000000000000;
    assign weights1[37][451] = 16'b1111111111110100;
    assign weights1[37][452] = 16'b1111111111111111;
    assign weights1[37][453] = 16'b0000000000011000;
    assign weights1[37][454] = 16'b0000000000010110;
    assign weights1[37][455] = 16'b0000000000000110;
    assign weights1[37][456] = 16'b0000000000001100;
    assign weights1[37][457] = 16'b1111111111110111;
    assign weights1[37][458] = 16'b1111111111101001;
    assign weights1[37][459] = 16'b1111111111110001;
    assign weights1[37][460] = 16'b0000000000000000;
    assign weights1[37][461] = 16'b1111111111111100;
    assign weights1[37][462] = 16'b1111111111101011;
    assign weights1[37][463] = 16'b1111111111100000;
    assign weights1[37][464] = 16'b1111111111110111;
    assign weights1[37][465] = 16'b1111111111110011;
    assign weights1[37][466] = 16'b0000000000011010;
    assign weights1[37][467] = 16'b0000000000011010;
    assign weights1[37][468] = 16'b0000000000001011;
    assign weights1[37][469] = 16'b0000000000001010;
    assign weights1[37][470] = 16'b0000000000001100;
    assign weights1[37][471] = 16'b1111111111111110;
    assign weights1[37][472] = 16'b1111111111101001;
    assign weights1[37][473] = 16'b1111111111111111;
    assign weights1[37][474] = 16'b0000000000000010;
    assign weights1[37][475] = 16'b1111111111111111;
    assign weights1[37][476] = 16'b1111111111111101;
    assign weights1[37][477] = 16'b0000000000000111;
    assign weights1[37][478] = 16'b0000000000001110;
    assign weights1[37][479] = 16'b0000000000000010;
    assign weights1[37][480] = 16'b0000000000000110;
    assign weights1[37][481] = 16'b0000000000011001;
    assign weights1[37][482] = 16'b0000000000001011;
    assign weights1[37][483] = 16'b1111111111111011;
    assign weights1[37][484] = 16'b1111111111111001;
    assign weights1[37][485] = 16'b1111111111011100;
    assign weights1[37][486] = 16'b1111111111101110;
    assign weights1[37][487] = 16'b0000000000000011;
    assign weights1[37][488] = 16'b0000000000010111;
    assign weights1[37][489] = 16'b0000000000001001;
    assign weights1[37][490] = 16'b1111111111111111;
    assign weights1[37][491] = 16'b1111111111101111;
    assign weights1[37][492] = 16'b1111111111011011;
    assign weights1[37][493] = 16'b1111111111100101;
    assign weights1[37][494] = 16'b0000000000000010;
    assign weights1[37][495] = 16'b0000000000010011;
    assign weights1[37][496] = 16'b0000000000010000;
    assign weights1[37][497] = 16'b0000000000001110;
    assign weights1[37][498] = 16'b1111111111111000;
    assign weights1[37][499] = 16'b1111111111101011;
    assign weights1[37][500] = 16'b1111111111101001;
    assign weights1[37][501] = 16'b1111111111011011;
    assign weights1[37][502] = 16'b1111111111110010;
    assign weights1[37][503] = 16'b1111111111111100;
    assign weights1[37][504] = 16'b0000000000001010;
    assign weights1[37][505] = 16'b0000000000010000;
    assign weights1[37][506] = 16'b0000000000010100;
    assign weights1[37][507] = 16'b0000000000010010;
    assign weights1[37][508] = 16'b0000000000101011;
    assign weights1[37][509] = 16'b0000000000100111;
    assign weights1[37][510] = 16'b1111111111111101;
    assign weights1[37][511] = 16'b0000000000010101;
    assign weights1[37][512] = 16'b1111111111101110;
    assign weights1[37][513] = 16'b1111111111001101;
    assign weights1[37][514] = 16'b1111111111110111;
    assign weights1[37][515] = 16'b1111111111110101;
    assign weights1[37][516] = 16'b0000000000100111;
    assign weights1[37][517] = 16'b0000000000100000;
    assign weights1[37][518] = 16'b1111111111110101;
    assign weights1[37][519] = 16'b1111111111100110;
    assign weights1[37][520] = 16'b1111111111011010;
    assign weights1[37][521] = 16'b1111111111010111;
    assign weights1[37][522] = 16'b0000000000001110;
    assign weights1[37][523] = 16'b0000000000101100;
    assign weights1[37][524] = 16'b0000000000000110;
    assign weights1[37][525] = 16'b0000000000100110;
    assign weights1[37][526] = 16'b0000000000010000;
    assign weights1[37][527] = 16'b1111111111111111;
    assign weights1[37][528] = 16'b1111111111100001;
    assign weights1[37][529] = 16'b1111111111100111;
    assign weights1[37][530] = 16'b1111111111100101;
    assign weights1[37][531] = 16'b1111111111111100;
    assign weights1[37][532] = 16'b0000000000010001;
    assign weights1[37][533] = 16'b0000000000010010;
    assign weights1[37][534] = 16'b0000000000011110;
    assign weights1[37][535] = 16'b0000000000101001;
    assign weights1[37][536] = 16'b0000000000101110;
    assign weights1[37][537] = 16'b0000000000100101;
    assign weights1[37][538] = 16'b1111111111111001;
    assign weights1[37][539] = 16'b1111111111011000;
    assign weights1[37][540] = 16'b1111111111011100;
    assign weights1[37][541] = 16'b1111111111011011;
    assign weights1[37][542] = 16'b1111111111110110;
    assign weights1[37][543] = 16'b0000000000001111;
    assign weights1[37][544] = 16'b0000000000100001;
    assign weights1[37][545] = 16'b0000000000011100;
    assign weights1[37][546] = 16'b1111111111110100;
    assign weights1[37][547] = 16'b1111111111011011;
    assign weights1[37][548] = 16'b1111111110111111;
    assign weights1[37][549] = 16'b1111111111001010;
    assign weights1[37][550] = 16'b0000000000001101;
    assign weights1[37][551] = 16'b0000000000100101;
    assign weights1[37][552] = 16'b0000000000000111;
    assign weights1[37][553] = 16'b0000000000101100;
    assign weights1[37][554] = 16'b0000000000001101;
    assign weights1[37][555] = 16'b0000000000001001;
    assign weights1[37][556] = 16'b0000000000000111;
    assign weights1[37][557] = 16'b1111111111010110;
    assign weights1[37][558] = 16'b1111111111100111;
    assign weights1[37][559] = 16'b1111111111110001;
    assign weights1[37][560] = 16'b0000000000001100;
    assign weights1[37][561] = 16'b0000000000011001;
    assign weights1[37][562] = 16'b0000000000100000;
    assign weights1[37][563] = 16'b0000000000011100;
    assign weights1[37][564] = 16'b0000000000010010;
    assign weights1[37][565] = 16'b0000000000000000;
    assign weights1[37][566] = 16'b1111111111101110;
    assign weights1[37][567] = 16'b1111111111001100;
    assign weights1[37][568] = 16'b1111111110110111;
    assign weights1[37][569] = 16'b1111111111010001;
    assign weights1[37][570] = 16'b1111111111101000;
    assign weights1[37][571] = 16'b0000000000100000;
    assign weights1[37][572] = 16'b0000000000111111;
    assign weights1[37][573] = 16'b0000000000001000;
    assign weights1[37][574] = 16'b1111111111111000;
    assign weights1[37][575] = 16'b1111111111000111;
    assign weights1[37][576] = 16'b1111111111000110;
    assign weights1[37][577] = 16'b1111111110110100;
    assign weights1[37][578] = 16'b0000000000001010;
    assign weights1[37][579] = 16'b0000000001000100;
    assign weights1[37][580] = 16'b0000000000010011;
    assign weights1[37][581] = 16'b0000000000010000;
    assign weights1[37][582] = 16'b0000000000100100;
    assign weights1[37][583] = 16'b0000000000010000;
    assign weights1[37][584] = 16'b1111111111111111;
    assign weights1[37][585] = 16'b1111111111011010;
    assign weights1[37][586] = 16'b1111111111101100;
    assign weights1[37][587] = 16'b1111111111101110;
    assign weights1[37][588] = 16'b0000000000000111;
    assign weights1[37][589] = 16'b0000000000001100;
    assign weights1[37][590] = 16'b0000000000011000;
    assign weights1[37][591] = 16'b0000000000000010;
    assign weights1[37][592] = 16'b0000000000000000;
    assign weights1[37][593] = 16'b1111111111011011;
    assign weights1[37][594] = 16'b1111111111001100;
    assign weights1[37][595] = 16'b1111111110011001;
    assign weights1[37][596] = 16'b1111111110010110;
    assign weights1[37][597] = 16'b1111111111111101;
    assign weights1[37][598] = 16'b0000000000011101;
    assign weights1[37][599] = 16'b0000000000110100;
    assign weights1[37][600] = 16'b0000000001010100;
    assign weights1[37][601] = 16'b0000000000000000;
    assign weights1[37][602] = 16'b1111111111011110;
    assign weights1[37][603] = 16'b1111111111010000;
    assign weights1[37][604] = 16'b1111111110000110;
    assign weights1[37][605] = 16'b1111111110010111;
    assign weights1[37][606] = 16'b0000000000101101;
    assign weights1[37][607] = 16'b0000000001001110;
    assign weights1[37][608] = 16'b0000000000011110;
    assign weights1[37][609] = 16'b0000000000001110;
    assign weights1[37][610] = 16'b0000000000010111;
    assign weights1[37][611] = 16'b0000000000001001;
    assign weights1[37][612] = 16'b0000000000011001;
    assign weights1[37][613] = 16'b1111111111011111;
    assign weights1[37][614] = 16'b1111111111111001;
    assign weights1[37][615] = 16'b1111111111101110;
    assign weights1[37][616] = 16'b1111111111111110;
    assign weights1[37][617] = 16'b1111111111111111;
    assign weights1[37][618] = 16'b1111111111111011;
    assign weights1[37][619] = 16'b1111111111010111;
    assign weights1[37][620] = 16'b1111111110111110;
    assign weights1[37][621] = 16'b1111111110110000;
    assign weights1[37][622] = 16'b1111111110000010;
    assign weights1[37][623] = 16'b1111111101011101;
    assign weights1[37][624] = 16'b1111111111011100;
    assign weights1[37][625] = 16'b1111111111111110;
    assign weights1[37][626] = 16'b0000000000110100;
    assign weights1[37][627] = 16'b0000000000110100;
    assign weights1[37][628] = 16'b0000000000111111;
    assign weights1[37][629] = 16'b1111111111110110;
    assign weights1[37][630] = 16'b1111111111001011;
    assign weights1[37][631] = 16'b1111111110110000;
    assign weights1[37][632] = 16'b1111111101001010;
    assign weights1[37][633] = 16'b1111111101110110;
    assign weights1[37][634] = 16'b0000000000100100;
    assign weights1[37][635] = 16'b0000000001100100;
    assign weights1[37][636] = 16'b0000000000010111;
    assign weights1[37][637] = 16'b0000000000100111;
    assign weights1[37][638] = 16'b0000000000100011;
    assign weights1[37][639] = 16'b0000000000001110;
    assign weights1[37][640] = 16'b1111111111110110;
    assign weights1[37][641] = 16'b1111111111111001;
    assign weights1[37][642] = 16'b1111111111101101;
    assign weights1[37][643] = 16'b1111111111111001;
    assign weights1[37][644] = 16'b1111111111111000;
    assign weights1[37][645] = 16'b1111111111101010;
    assign weights1[37][646] = 16'b1111111111011100;
    assign weights1[37][647] = 16'b1111111111001011;
    assign weights1[37][648] = 16'b1111111110111000;
    assign weights1[37][649] = 16'b1111111110010101;
    assign weights1[37][650] = 16'b1111111101110110;
    assign weights1[37][651] = 16'b1111111110100101;
    assign weights1[37][652] = 16'b0000000000000000;
    assign weights1[37][653] = 16'b0000000000011101;
    assign weights1[37][654] = 16'b0000000000100101;
    assign weights1[37][655] = 16'b0000000000111001;
    assign weights1[37][656] = 16'b0000000000110111;
    assign weights1[37][657] = 16'b0000000000001101;
    assign weights1[37][658] = 16'b1111111110110010;
    assign weights1[37][659] = 16'b1111111101111011;
    assign weights1[37][660] = 16'b1111111101001101;
    assign weights1[37][661] = 16'b1111111110100100;
    assign weights1[37][662] = 16'b0000000001000111;
    assign weights1[37][663] = 16'b0000000001000111;
    assign weights1[37][664] = 16'b0000000000011110;
    assign weights1[37][665] = 16'b0000000000101111;
    assign weights1[37][666] = 16'b0000000000001010;
    assign weights1[37][667] = 16'b0000000000000110;
    assign weights1[37][668] = 16'b0000000000010001;
    assign weights1[37][669] = 16'b0000000000000011;
    assign weights1[37][670] = 16'b1111111111110110;
    assign weights1[37][671] = 16'b1111111111111100;
    assign weights1[37][672] = 16'b1111111111110101;
    assign weights1[37][673] = 16'b1111111111100111;
    assign weights1[37][674] = 16'b1111111111011001;
    assign weights1[37][675] = 16'b1111111111000011;
    assign weights1[37][676] = 16'b1111111110101100;
    assign weights1[37][677] = 16'b1111111110000110;
    assign weights1[37][678] = 16'b1111111110100110;
    assign weights1[37][679] = 16'b1111111111101100;
    assign weights1[37][680] = 16'b0000000001000111;
    assign weights1[37][681] = 16'b0000000000101010;
    assign weights1[37][682] = 16'b0000000000010010;
    assign weights1[37][683] = 16'b0000000000100011;
    assign weights1[37][684] = 16'b0000000000100101;
    assign weights1[37][685] = 16'b1111111110110010;
    assign weights1[37][686] = 16'b1111111110100100;
    assign weights1[37][687] = 16'b1111111101100101;
    assign weights1[37][688] = 16'b1111111101010001;
    assign weights1[37][689] = 16'b1111111110101011;
    assign weights1[37][690] = 16'b0000000000010110;
    assign weights1[37][691] = 16'b0000000000111001;
    assign weights1[37][692] = 16'b0000000000011100;
    assign weights1[37][693] = 16'b1111111111111010;
    assign weights1[37][694] = 16'b0000000000011101;
    assign weights1[37][695] = 16'b0000000000101011;
    assign weights1[37][696] = 16'b0000000000011101;
    assign weights1[37][697] = 16'b0000000000000110;
    assign weights1[37][698] = 16'b1111111111111100;
    assign weights1[37][699] = 16'b1111111111111010;
    assign weights1[37][700] = 16'b1111111111111100;
    assign weights1[37][701] = 16'b1111111111101101;
    assign weights1[37][702] = 16'b1111111111100010;
    assign weights1[37][703] = 16'b1111111111000001;
    assign weights1[37][704] = 16'b1111111110100011;
    assign weights1[37][705] = 16'b1111111110100011;
    assign weights1[37][706] = 16'b1111111111011001;
    assign weights1[37][707] = 16'b1111111111111101;
    assign weights1[37][708] = 16'b0000000000111100;
    assign weights1[37][709] = 16'b0000000001000111;
    assign weights1[37][710] = 16'b0000000000101011;
    assign weights1[37][711] = 16'b0000000000111111;
    assign weights1[37][712] = 16'b0000000000011101;
    assign weights1[37][713] = 16'b1111111111000000;
    assign weights1[37][714] = 16'b1111111110010001;
    assign weights1[37][715] = 16'b1111111101010100;
    assign weights1[37][716] = 16'b1111111100101110;
    assign weights1[37][717] = 16'b1111111110111011;
    assign weights1[37][718] = 16'b0000000000000000;
    assign weights1[37][719] = 16'b0000000000111111;
    assign weights1[37][720] = 16'b0000000000101100;
    assign weights1[37][721] = 16'b0000000000011000;
    assign weights1[37][722] = 16'b0000000000011001;
    assign weights1[37][723] = 16'b0000000000100101;
    assign weights1[37][724] = 16'b0000000000011000;
    assign weights1[37][725] = 16'b0000000000001000;
    assign weights1[37][726] = 16'b1111111111111011;
    assign weights1[37][727] = 16'b1111111111111011;
    assign weights1[37][728] = 16'b1111111111111011;
    assign weights1[37][729] = 16'b1111111111110001;
    assign weights1[37][730] = 16'b1111111111100001;
    assign weights1[37][731] = 16'b1111111111001101;
    assign weights1[37][732] = 16'b1111111111001000;
    assign weights1[37][733] = 16'b1111111111001110;
    assign weights1[37][734] = 16'b1111111111111001;
    assign weights1[37][735] = 16'b0000000000100101;
    assign weights1[37][736] = 16'b0000000000011100;
    assign weights1[37][737] = 16'b0000000000001111;
    assign weights1[37][738] = 16'b0000000000011110;
    assign weights1[37][739] = 16'b0000000000010011;
    assign weights1[37][740] = 16'b1111111111100111;
    assign weights1[37][741] = 16'b1111111111010010;
    assign weights1[37][742] = 16'b1111111110000101;
    assign weights1[37][743] = 16'b1111111101101011;
    assign weights1[37][744] = 16'b1111111101110001;
    assign weights1[37][745] = 16'b1111111111000110;
    assign weights1[37][746] = 16'b1111111111111010;
    assign weights1[37][747] = 16'b0000000000001100;
    assign weights1[37][748] = 16'b0000000000010010;
    assign weights1[37][749] = 16'b0000000000001110;
    assign weights1[37][750] = 16'b0000000000011010;
    assign weights1[37][751] = 16'b0000000000100011;
    assign weights1[37][752] = 16'b0000000000010110;
    assign weights1[37][753] = 16'b0000000000001111;
    assign weights1[37][754] = 16'b0000000000000111;
    assign weights1[37][755] = 16'b0000000000000000;
    assign weights1[37][756] = 16'b1111111111111110;
    assign weights1[37][757] = 16'b1111111111110110;
    assign weights1[37][758] = 16'b1111111111101011;
    assign weights1[37][759] = 16'b1111111111100101;
    assign weights1[37][760] = 16'b1111111111110000;
    assign weights1[37][761] = 16'b1111111111111001;
    assign weights1[37][762] = 16'b0000000000100000;
    assign weights1[37][763] = 16'b0000000000101100;
    assign weights1[37][764] = 16'b0000000000101000;
    assign weights1[37][765] = 16'b0000000000101010;
    assign weights1[37][766] = 16'b1111111111111011;
    assign weights1[37][767] = 16'b1111111111110011;
    assign weights1[37][768] = 16'b1111111111010111;
    assign weights1[37][769] = 16'b1111111110100101;
    assign weights1[37][770] = 16'b1111111101101100;
    assign weights1[37][771] = 16'b1111111101001101;
    assign weights1[37][772] = 16'b1111111101011101;
    assign weights1[37][773] = 16'b1111111110100001;
    assign weights1[37][774] = 16'b1111111111010011;
    assign weights1[37][775] = 16'b1111111111101110;
    assign weights1[37][776] = 16'b0000000000001100;
    assign weights1[37][777] = 16'b0000000000011011;
    assign weights1[37][778] = 16'b0000000000011110;
    assign weights1[37][779] = 16'b0000000000100100;
    assign weights1[37][780] = 16'b0000000000100111;
    assign weights1[37][781] = 16'b0000000000001101;
    assign weights1[37][782] = 16'b0000000000001001;
    assign weights1[37][783] = 16'b0000000000000011;
    assign weights1[38][0] = 16'b0000000000000000;
    assign weights1[38][1] = 16'b0000000000000000;
    assign weights1[38][2] = 16'b0000000000000000;
    assign weights1[38][3] = 16'b0000000000000000;
    assign weights1[38][4] = 16'b1111111111111111;
    assign weights1[38][5] = 16'b1111111111111111;
    assign weights1[38][6] = 16'b0000000000000000;
    assign weights1[38][7] = 16'b1111111111111111;
    assign weights1[38][8] = 16'b0000000000000010;
    assign weights1[38][9] = 16'b0000000000000001;
    assign weights1[38][10] = 16'b1111111111111111;
    assign weights1[38][11] = 16'b0000000000000100;
    assign weights1[38][12] = 16'b0000000000001100;
    assign weights1[38][13] = 16'b0000000000001010;
    assign weights1[38][14] = 16'b0000000000010110;
    assign weights1[38][15] = 16'b0000000000011011;
    assign weights1[38][16] = 16'b0000000000010111;
    assign weights1[38][17] = 16'b0000000000001001;
    assign weights1[38][18] = 16'b0000000000001000;
    assign weights1[38][19] = 16'b0000000000001100;
    assign weights1[38][20] = 16'b0000000000001001;
    assign weights1[38][21] = 16'b1111111111111110;
    assign weights1[38][22] = 16'b1111111111111010;
    assign weights1[38][23] = 16'b1111111111111111;
    assign weights1[38][24] = 16'b1111111111111101;
    assign weights1[38][25] = 16'b1111111111111111;
    assign weights1[38][26] = 16'b1111111111111111;
    assign weights1[38][27] = 16'b0000000000000000;
    assign weights1[38][28] = 16'b0000000000000000;
    assign weights1[38][29] = 16'b0000000000000000;
    assign weights1[38][30] = 16'b0000000000000000;
    assign weights1[38][31] = 16'b1111111111111110;
    assign weights1[38][32] = 16'b1111111111111111;
    assign weights1[38][33] = 16'b1111111111111100;
    assign weights1[38][34] = 16'b0000000000000000;
    assign weights1[38][35] = 16'b1111111111111110;
    assign weights1[38][36] = 16'b1111111111111110;
    assign weights1[38][37] = 16'b1111111111111100;
    assign weights1[38][38] = 16'b0000000000000000;
    assign weights1[38][39] = 16'b0000000000001000;
    assign weights1[38][40] = 16'b0000000000001100;
    assign weights1[38][41] = 16'b0000000000001111;
    assign weights1[38][42] = 16'b0000000000001011;
    assign weights1[38][43] = 16'b0000000000011000;
    assign weights1[38][44] = 16'b0000000000010010;
    assign weights1[38][45] = 16'b0000000000001010;
    assign weights1[38][46] = 16'b0000000000001000;
    assign weights1[38][47] = 16'b0000000000000101;
    assign weights1[38][48] = 16'b0000000000001001;
    assign weights1[38][49] = 16'b0000000000000100;
    assign weights1[38][50] = 16'b0000000000000011;
    assign weights1[38][51] = 16'b1111111111111110;
    assign weights1[38][52] = 16'b1111111111111010;
    assign weights1[38][53] = 16'b1111111111111100;
    assign weights1[38][54] = 16'b1111111111111111;
    assign weights1[38][55] = 16'b0000000000000000;
    assign weights1[38][56] = 16'b0000000000000000;
    assign weights1[38][57] = 16'b0000000000000000;
    assign weights1[38][58] = 16'b1111111111111110;
    assign weights1[38][59] = 16'b1111111111111011;
    assign weights1[38][60] = 16'b1111111111111101;
    assign weights1[38][61] = 16'b1111111111111101;
    assign weights1[38][62] = 16'b1111111111111100;
    assign weights1[38][63] = 16'b1111111111111101;
    assign weights1[38][64] = 16'b1111111111111001;
    assign weights1[38][65] = 16'b1111111111110101;
    assign weights1[38][66] = 16'b1111111111110110;
    assign weights1[38][67] = 16'b0000000000000000;
    assign weights1[38][68] = 16'b0000000000000111;
    assign weights1[38][69] = 16'b0000000000010100;
    assign weights1[38][70] = 16'b0000000000011000;
    assign weights1[38][71] = 16'b0000000000011100;
    assign weights1[38][72] = 16'b0000000000010000;
    assign weights1[38][73] = 16'b0000000000001010;
    assign weights1[38][74] = 16'b0000000000001011;
    assign weights1[38][75] = 16'b0000000000000100;
    assign weights1[38][76] = 16'b0000000000000000;
    assign weights1[38][77] = 16'b1111111111111010;
    assign weights1[38][78] = 16'b1111111111101110;
    assign weights1[38][79] = 16'b1111111111101110;
    assign weights1[38][80] = 16'b1111111111110010;
    assign weights1[38][81] = 16'b1111111111111011;
    assign weights1[38][82] = 16'b1111111111111110;
    assign weights1[38][83] = 16'b1111111111111111;
    assign weights1[38][84] = 16'b0000000000000000;
    assign weights1[38][85] = 16'b0000000000000000;
    assign weights1[38][86] = 16'b1111111111111101;
    assign weights1[38][87] = 16'b1111111111111101;
    assign weights1[38][88] = 16'b1111111111111010;
    assign weights1[38][89] = 16'b1111111111111101;
    assign weights1[38][90] = 16'b1111111111110110;
    assign weights1[38][91] = 16'b1111111111110100;
    assign weights1[38][92] = 16'b1111111111110100;
    assign weights1[38][93] = 16'b1111111111101101;
    assign weights1[38][94] = 16'b1111111111101010;
    assign weights1[38][95] = 16'b1111111111111000;
    assign weights1[38][96] = 16'b1111111111111111;
    assign weights1[38][97] = 16'b0000000000001011;
    assign weights1[38][98] = 16'b0000000000001011;
    assign weights1[38][99] = 16'b0000000000001101;
    assign weights1[38][100] = 16'b0000000000001001;
    assign weights1[38][101] = 16'b0000000000000011;
    assign weights1[38][102] = 16'b0000000000000011;
    assign weights1[38][103] = 16'b1111111111111100;
    assign weights1[38][104] = 16'b1111111111111101;
    assign weights1[38][105] = 16'b1111111111111100;
    assign weights1[38][106] = 16'b1111111111100111;
    assign weights1[38][107] = 16'b1111111111100110;
    assign weights1[38][108] = 16'b1111111111101111;
    assign weights1[38][109] = 16'b1111111111110101;
    assign weights1[38][110] = 16'b1111111111111010;
    assign weights1[38][111] = 16'b1111111111111111;
    assign weights1[38][112] = 16'b0000000000000000;
    assign weights1[38][113] = 16'b0000000000000001;
    assign weights1[38][114] = 16'b1111111111111110;
    assign weights1[38][115] = 16'b1111111111111000;
    assign weights1[38][116] = 16'b1111111111111011;
    assign weights1[38][117] = 16'b1111111111111000;
    assign weights1[38][118] = 16'b1111111111101110;
    assign weights1[38][119] = 16'b1111111111101001;
    assign weights1[38][120] = 16'b1111111111101010;
    assign weights1[38][121] = 16'b1111111111100111;
    assign weights1[38][122] = 16'b1111111111101011;
    assign weights1[38][123] = 16'b1111111111110100;
    assign weights1[38][124] = 16'b1111111111111101;
    assign weights1[38][125] = 16'b1111111111111100;
    assign weights1[38][126] = 16'b0000000000001000;
    assign weights1[38][127] = 16'b1111111111111111;
    assign weights1[38][128] = 16'b1111111111110111;
    assign weights1[38][129] = 16'b0000000000000100;
    assign weights1[38][130] = 16'b1111111111111010;
    assign weights1[38][131] = 16'b1111111111110100;
    assign weights1[38][132] = 16'b1111111111101101;
    assign weights1[38][133] = 16'b1111111111101001;
    assign weights1[38][134] = 16'b1111111111101011;
    assign weights1[38][135] = 16'b1111111111101001;
    assign weights1[38][136] = 16'b1111111111101100;
    assign weights1[38][137] = 16'b1111111111110111;
    assign weights1[38][138] = 16'b1111111111111001;
    assign weights1[38][139] = 16'b1111111111111110;
    assign weights1[38][140] = 16'b0000000000000001;
    assign weights1[38][141] = 16'b0000000000000010;
    assign weights1[38][142] = 16'b1111111111111101;
    assign weights1[38][143] = 16'b1111111111111100;
    assign weights1[38][144] = 16'b1111111111110110;
    assign weights1[38][145] = 16'b1111111111111100;
    assign weights1[38][146] = 16'b1111111111111000;
    assign weights1[38][147] = 16'b1111111111110111;
    assign weights1[38][148] = 16'b1111111111101100;
    assign weights1[38][149] = 16'b1111111111100110;
    assign weights1[38][150] = 16'b1111111111101000;
    assign weights1[38][151] = 16'b1111111111110100;
    assign weights1[38][152] = 16'b1111111111110011;
    assign weights1[38][153] = 16'b0000000000000001;
    assign weights1[38][154] = 16'b1111111111111100;
    assign weights1[38][155] = 16'b0000000000000111;
    assign weights1[38][156] = 16'b0000000000000101;
    assign weights1[38][157] = 16'b0000000000001011;
    assign weights1[38][158] = 16'b0000000000000001;
    assign weights1[38][159] = 16'b1111111111110101;
    assign weights1[38][160] = 16'b1111111111110101;
    assign weights1[38][161] = 16'b1111111111101100;
    assign weights1[38][162] = 16'b1111111111011001;
    assign weights1[38][163] = 16'b1111111111100011;
    assign weights1[38][164] = 16'b1111111111110010;
    assign weights1[38][165] = 16'b1111111111110101;
    assign weights1[38][166] = 16'b1111111111111100;
    assign weights1[38][167] = 16'b0000000000000000;
    assign weights1[38][168] = 16'b0000000000000000;
    assign weights1[38][169] = 16'b0000000000000000;
    assign weights1[38][170] = 16'b0000000000000001;
    assign weights1[38][171] = 16'b1111111111111101;
    assign weights1[38][172] = 16'b1111111111111001;
    assign weights1[38][173] = 16'b1111111111111101;
    assign weights1[38][174] = 16'b1111111111110100;
    assign weights1[38][175] = 16'b1111111111110000;
    assign weights1[38][176] = 16'b1111111111101101;
    assign weights1[38][177] = 16'b1111111111101110;
    assign weights1[38][178] = 16'b1111111111101010;
    assign weights1[38][179] = 16'b1111111111100111;
    assign weights1[38][180] = 16'b1111111111101111;
    assign weights1[38][181] = 16'b1111111111110100;
    assign weights1[38][182] = 16'b1111111111111111;
    assign weights1[38][183] = 16'b0000000000001011;
    assign weights1[38][184] = 16'b0000000000010110;
    assign weights1[38][185] = 16'b0000000000000111;
    assign weights1[38][186] = 16'b1111111111111000;
    assign weights1[38][187] = 16'b1111111111110010;
    assign weights1[38][188] = 16'b1111111111101100;
    assign weights1[38][189] = 16'b1111111111100011;
    assign weights1[38][190] = 16'b1111111111011011;
    assign weights1[38][191] = 16'b1111111111101000;
    assign weights1[38][192] = 16'b1111111111101100;
    assign weights1[38][193] = 16'b1111111111110111;
    assign weights1[38][194] = 16'b1111111111111100;
    assign weights1[38][195] = 16'b1111111111111111;
    assign weights1[38][196] = 16'b0000000000000001;
    assign weights1[38][197] = 16'b0000000000000000;
    assign weights1[38][198] = 16'b0000000000000000;
    assign weights1[38][199] = 16'b1111111111111101;
    assign weights1[38][200] = 16'b0000000000000000;
    assign weights1[38][201] = 16'b1111111111111101;
    assign weights1[38][202] = 16'b1111111111110001;
    assign weights1[38][203] = 16'b1111111111110110;
    assign weights1[38][204] = 16'b1111111111101101;
    assign weights1[38][205] = 16'b1111111111100011;
    assign weights1[38][206] = 16'b1111111111100000;
    assign weights1[38][207] = 16'b1111111111011011;
    assign weights1[38][208] = 16'b1111111111011101;
    assign weights1[38][209] = 16'b1111111111100110;
    assign weights1[38][210] = 16'b1111111111100111;
    assign weights1[38][211] = 16'b1111111111111111;
    assign weights1[38][212] = 16'b0000000000001101;
    assign weights1[38][213] = 16'b0000000000001111;
    assign weights1[38][214] = 16'b1111111111111100;
    assign weights1[38][215] = 16'b1111111111101111;
    assign weights1[38][216] = 16'b1111111111100111;
    assign weights1[38][217] = 16'b1111111111011010;
    assign weights1[38][218] = 16'b1111111111010111;
    assign weights1[38][219] = 16'b1111111111100111;
    assign weights1[38][220] = 16'b1111111111101100;
    assign weights1[38][221] = 16'b1111111111111000;
    assign weights1[38][222] = 16'b1111111111111110;
    assign weights1[38][223] = 16'b1111111111111111;
    assign weights1[38][224] = 16'b0000000000000000;
    assign weights1[38][225] = 16'b0000000000000000;
    assign weights1[38][226] = 16'b0000000000000000;
    assign weights1[38][227] = 16'b0000000000000000;
    assign weights1[38][228] = 16'b0000000000000011;
    assign weights1[38][229] = 16'b0000000000000010;
    assign weights1[38][230] = 16'b1111111111111010;
    assign weights1[38][231] = 16'b1111111111111100;
    assign weights1[38][232] = 16'b1111111111101101;
    assign weights1[38][233] = 16'b1111111111100001;
    assign weights1[38][234] = 16'b1111111111011100;
    assign weights1[38][235] = 16'b1111111111011000;
    assign weights1[38][236] = 16'b1111111111100101;
    assign weights1[38][237] = 16'b1111111111101011;
    assign weights1[38][238] = 16'b1111111111110011;
    assign weights1[38][239] = 16'b0000000000000100;
    assign weights1[38][240] = 16'b0000000000010011;
    assign weights1[38][241] = 16'b0000000000010011;
    assign weights1[38][242] = 16'b0000000000000110;
    assign weights1[38][243] = 16'b0000000000000001;
    assign weights1[38][244] = 16'b1111111111101011;
    assign weights1[38][245] = 16'b1111111111101101;
    assign weights1[38][246] = 16'b1111111111011100;
    assign weights1[38][247] = 16'b1111111111100101;
    assign weights1[38][248] = 16'b1111111111101100;
    assign weights1[38][249] = 16'b1111111111110010;
    assign weights1[38][250] = 16'b1111111111111000;
    assign weights1[38][251] = 16'b1111111111111100;
    assign weights1[38][252] = 16'b1111111111111110;
    assign weights1[38][253] = 16'b0000000000000010;
    assign weights1[38][254] = 16'b0000000000001001;
    assign weights1[38][255] = 16'b0000000000000010;
    assign weights1[38][256] = 16'b0000000000000100;
    assign weights1[38][257] = 16'b0000000000000111;
    assign weights1[38][258] = 16'b1111111111111111;
    assign weights1[38][259] = 16'b1111111111110101;
    assign weights1[38][260] = 16'b1111111111101100;
    assign weights1[38][261] = 16'b1111111111011011;
    assign weights1[38][262] = 16'b1111111111011011;
    assign weights1[38][263] = 16'b1111111111101010;
    assign weights1[38][264] = 16'b0000000000000000;
    assign weights1[38][265] = 16'b1111111111111010;
    assign weights1[38][266] = 16'b1111111111111001;
    assign weights1[38][267] = 16'b0000000000000100;
    assign weights1[38][268] = 16'b0000000000000111;
    assign weights1[38][269] = 16'b0000000000011000;
    assign weights1[38][270] = 16'b0000000000001000;
    assign weights1[38][271] = 16'b1111111111111101;
    assign weights1[38][272] = 16'b1111111111101011;
    assign weights1[38][273] = 16'b1111111111100101;
    assign weights1[38][274] = 16'b1111111111011011;
    assign weights1[38][275] = 16'b1111111111010101;
    assign weights1[38][276] = 16'b1111111111100101;
    assign weights1[38][277] = 16'b1111111111110101;
    assign weights1[38][278] = 16'b1111111111111000;
    assign weights1[38][279] = 16'b1111111111111100;
    assign weights1[38][280] = 16'b0000000000000010;
    assign weights1[38][281] = 16'b0000000000000011;
    assign weights1[38][282] = 16'b0000000000000110;
    assign weights1[38][283] = 16'b0000000000000011;
    assign weights1[38][284] = 16'b0000000000000110;
    assign weights1[38][285] = 16'b1111111111111000;
    assign weights1[38][286] = 16'b1111111111111000;
    assign weights1[38][287] = 16'b1111111111101111;
    assign weights1[38][288] = 16'b1111111111101101;
    assign weights1[38][289] = 16'b1111111111101100;
    assign weights1[38][290] = 16'b1111111111100000;
    assign weights1[38][291] = 16'b1111111111111011;
    assign weights1[38][292] = 16'b1111111111111001;
    assign weights1[38][293] = 16'b1111111111111000;
    assign weights1[38][294] = 16'b1111111111100111;
    assign weights1[38][295] = 16'b1111111111110010;
    assign weights1[38][296] = 16'b1111111111111111;
    assign weights1[38][297] = 16'b0000000000010100;
    assign weights1[38][298] = 16'b0000000000001001;
    assign weights1[38][299] = 16'b1111111111110100;
    assign weights1[38][300] = 16'b1111111111101010;
    assign weights1[38][301] = 16'b1111111111011001;
    assign weights1[38][302] = 16'b1111111111010001;
    assign weights1[38][303] = 16'b1111111111010010;
    assign weights1[38][304] = 16'b1111111111100010;
    assign weights1[38][305] = 16'b1111111111101001;
    assign weights1[38][306] = 16'b1111111111110010;
    assign weights1[38][307] = 16'b1111111111111100;
    assign weights1[38][308] = 16'b0000000000000001;
    assign weights1[38][309] = 16'b1111111111111111;
    assign weights1[38][310] = 16'b0000000000000100;
    assign weights1[38][311] = 16'b0000000000000101;
    assign weights1[38][312] = 16'b1111111111111111;
    assign weights1[38][313] = 16'b1111111111111101;
    assign weights1[38][314] = 16'b1111111111111010;
    assign weights1[38][315] = 16'b1111111111101100;
    assign weights1[38][316] = 16'b1111111111100000;
    assign weights1[38][317] = 16'b1111111111101010;
    assign weights1[38][318] = 16'b1111111111100010;
    assign weights1[38][319] = 16'b1111111111111100;
    assign weights1[38][320] = 16'b1111111111111010;
    assign weights1[38][321] = 16'b1111111111110011;
    assign weights1[38][322] = 16'b1111111111101011;
    assign weights1[38][323] = 16'b1111111111110110;
    assign weights1[38][324] = 16'b0000000000010101;
    assign weights1[38][325] = 16'b0000000000100001;
    assign weights1[38][326] = 16'b0000000000001011;
    assign weights1[38][327] = 16'b0000000000000010;
    assign weights1[38][328] = 16'b1111111111110110;
    assign weights1[38][329] = 16'b1111111111011011;
    assign weights1[38][330] = 16'b1111111111001000;
    assign weights1[38][331] = 16'b1111111111010100;
    assign weights1[38][332] = 16'b1111111111100001;
    assign weights1[38][333] = 16'b1111111111101101;
    assign weights1[38][334] = 16'b1111111111110101;
    assign weights1[38][335] = 16'b1111111111111000;
    assign weights1[38][336] = 16'b0000000000000001;
    assign weights1[38][337] = 16'b1111111111111011;
    assign weights1[38][338] = 16'b1111111111111111;
    assign weights1[38][339] = 16'b0000000000001000;
    assign weights1[38][340] = 16'b0000000000000010;
    assign weights1[38][341] = 16'b0000000000000101;
    assign weights1[38][342] = 16'b1111111111111000;
    assign weights1[38][343] = 16'b1111111111101101;
    assign weights1[38][344] = 16'b1111111111101000;
    assign weights1[38][345] = 16'b1111111111101110;
    assign weights1[38][346] = 16'b1111111111111001;
    assign weights1[38][347] = 16'b1111111111111110;
    assign weights1[38][348] = 16'b1111111111110010;
    assign weights1[38][349] = 16'b1111111111100011;
    assign weights1[38][350] = 16'b1111111111101010;
    assign weights1[38][351] = 16'b0000000000000100;
    assign weights1[38][352] = 16'b0000000000011100;
    assign weights1[38][353] = 16'b0000000000011000;
    assign weights1[38][354] = 16'b0000000000000110;
    assign weights1[38][355] = 16'b0000000000000000;
    assign weights1[38][356] = 16'b1111111111110011;
    assign weights1[38][357] = 16'b1111111111100010;
    assign weights1[38][358] = 16'b1111111111010001;
    assign weights1[38][359] = 16'b1111111111010100;
    assign weights1[38][360] = 16'b1111111111100110;
    assign weights1[38][361] = 16'b1111111111101110;
    assign weights1[38][362] = 16'b1111111111110100;
    assign weights1[38][363] = 16'b1111111111111010;
    assign weights1[38][364] = 16'b1111111111111111;
    assign weights1[38][365] = 16'b0000000000000000;
    assign weights1[38][366] = 16'b0000000000000011;
    assign weights1[38][367] = 16'b0000000000000001;
    assign weights1[38][368] = 16'b0000000000000001;
    assign weights1[38][369] = 16'b0000000000000111;
    assign weights1[38][370] = 16'b1111111111111111;
    assign weights1[38][371] = 16'b1111111111110010;
    assign weights1[38][372] = 16'b1111111111111011;
    assign weights1[38][373] = 16'b1111111111110101;
    assign weights1[38][374] = 16'b0000000000000000;
    assign weights1[38][375] = 16'b1111111111111010;
    assign weights1[38][376] = 16'b1111111111110000;
    assign weights1[38][377] = 16'b1111111111101000;
    assign weights1[38][378] = 16'b1111111111101011;
    assign weights1[38][379] = 16'b0000000000000111;
    assign weights1[38][380] = 16'b0000000000011001;
    assign weights1[38][381] = 16'b0000000000011000;
    assign weights1[38][382] = 16'b0000000000010000;
    assign weights1[38][383] = 16'b0000000000000100;
    assign weights1[38][384] = 16'b1111111111101110;
    assign weights1[38][385] = 16'b1111111111100000;
    assign weights1[38][386] = 16'b1111111111011110;
    assign weights1[38][387] = 16'b1111111111101010;
    assign weights1[38][388] = 16'b1111111111101100;
    assign weights1[38][389] = 16'b1111111111110111;
    assign weights1[38][390] = 16'b1111111111111001;
    assign weights1[38][391] = 16'b1111111111111111;
    assign weights1[38][392] = 16'b0000000000000001;
    assign weights1[38][393] = 16'b0000000000000010;
    assign weights1[38][394] = 16'b0000000000000000;
    assign weights1[38][395] = 16'b0000000000000011;
    assign weights1[38][396] = 16'b1111111111111101;
    assign weights1[38][397] = 16'b0000000000000101;
    assign weights1[38][398] = 16'b1111111111111011;
    assign weights1[38][399] = 16'b0000000000000000;
    assign weights1[38][400] = 16'b1111111111111110;
    assign weights1[38][401] = 16'b0000000000000110;
    assign weights1[38][402] = 16'b0000000000000000;
    assign weights1[38][403] = 16'b1111111111111010;
    assign weights1[38][404] = 16'b1111111111101010;
    assign weights1[38][405] = 16'b1111111111010111;
    assign weights1[38][406] = 16'b1111111111100100;
    assign weights1[38][407] = 16'b0000000000000000;
    assign weights1[38][408] = 16'b0000000000011010;
    assign weights1[38][409] = 16'b0000000000011011;
    assign weights1[38][410] = 16'b0000000000001100;
    assign weights1[38][411] = 16'b0000000000000111;
    assign weights1[38][412] = 16'b1111111111111011;
    assign weights1[38][413] = 16'b1111111111101100;
    assign weights1[38][414] = 16'b1111111111100001;
    assign weights1[38][415] = 16'b1111111111110110;
    assign weights1[38][416] = 16'b1111111111111000;
    assign weights1[38][417] = 16'b1111111111111100;
    assign weights1[38][418] = 16'b1111111111111110;
    assign weights1[38][419] = 16'b1111111111111100;
    assign weights1[38][420] = 16'b0000000000000011;
    assign weights1[38][421] = 16'b1111111111111110;
    assign weights1[38][422] = 16'b0000000000000010;
    assign weights1[38][423] = 16'b1111111111111100;
    assign weights1[38][424] = 16'b1111111111111100;
    assign weights1[38][425] = 16'b0000000000000011;
    assign weights1[38][426] = 16'b0000000000000100;
    assign weights1[38][427] = 16'b1111111111111110;
    assign weights1[38][428] = 16'b0000000000000101;
    assign weights1[38][429] = 16'b0000000000000001;
    assign weights1[38][430] = 16'b0000000000000011;
    assign weights1[38][431] = 16'b1111111111110101;
    assign weights1[38][432] = 16'b1111111111100100;
    assign weights1[38][433] = 16'b1111111111010001;
    assign weights1[38][434] = 16'b1111111111101011;
    assign weights1[38][435] = 16'b0000000000001011;
    assign weights1[38][436] = 16'b0000000000011111;
    assign weights1[38][437] = 16'b0000000000011110;
    assign weights1[38][438] = 16'b0000000000001110;
    assign weights1[38][439] = 16'b0000000000000001;
    assign weights1[38][440] = 16'b1111111111110010;
    assign weights1[38][441] = 16'b1111111111100101;
    assign weights1[38][442] = 16'b1111111111110001;
    assign weights1[38][443] = 16'b1111111111111011;
    assign weights1[38][444] = 16'b1111111111111000;
    assign weights1[38][445] = 16'b0000000000000001;
    assign weights1[38][446] = 16'b0000000000000001;
    assign weights1[38][447] = 16'b1111111111111011;
    assign weights1[38][448] = 16'b0000000000000101;
    assign weights1[38][449] = 16'b1111111111111011;
    assign weights1[38][450] = 16'b0000000000000011;
    assign weights1[38][451] = 16'b1111111111111001;
    assign weights1[38][452] = 16'b1111111111111111;
    assign weights1[38][453] = 16'b0000000000000000;
    assign weights1[38][454] = 16'b0000000000001011;
    assign weights1[38][455] = 16'b0000000000010000;
    assign weights1[38][456] = 16'b1111111111111100;
    assign weights1[38][457] = 16'b1111111111111001;
    assign weights1[38][458] = 16'b1111111111111001;
    assign weights1[38][459] = 16'b1111111111011100;
    assign weights1[38][460] = 16'b1111111111100100;
    assign weights1[38][461] = 16'b1111111111010100;
    assign weights1[38][462] = 16'b1111111111100010;
    assign weights1[38][463] = 16'b0000000000010011;
    assign weights1[38][464] = 16'b0000000000010010;
    assign weights1[38][465] = 16'b0000000000011001;
    assign weights1[38][466] = 16'b0000000000010110;
    assign weights1[38][467] = 16'b0000000000001000;
    assign weights1[38][468] = 16'b1111111111111110;
    assign weights1[38][469] = 16'b1111111111110010;
    assign weights1[38][470] = 16'b1111111111110100;
    assign weights1[38][471] = 16'b1111111111111111;
    assign weights1[38][472] = 16'b0000000000000011;
    assign weights1[38][473] = 16'b0000000000001000;
    assign weights1[38][474] = 16'b0000000000000000;
    assign weights1[38][475] = 16'b1111111111111101;
    assign weights1[38][476] = 16'b0000000000000001;
    assign weights1[38][477] = 16'b0000000000000000;
    assign weights1[38][478] = 16'b1111111111111111;
    assign weights1[38][479] = 16'b1111111111111101;
    assign weights1[38][480] = 16'b0000000000000110;
    assign weights1[38][481] = 16'b0000000000000010;
    assign weights1[38][482] = 16'b0000000000000001;
    assign weights1[38][483] = 16'b0000000000000011;
    assign weights1[38][484] = 16'b1111111111111011;
    assign weights1[38][485] = 16'b1111111111111000;
    assign weights1[38][486] = 16'b1111111111101111;
    assign weights1[38][487] = 16'b1111111111100100;
    assign weights1[38][488] = 16'b1111111111100000;
    assign weights1[38][489] = 16'b1111111111001001;
    assign weights1[38][490] = 16'b1111111111101001;
    assign weights1[38][491] = 16'b0000000000010110;
    assign weights1[38][492] = 16'b0000000000010010;
    assign weights1[38][493] = 16'b0000000000010110;
    assign weights1[38][494] = 16'b0000000000001110;
    assign weights1[38][495] = 16'b1111111111111010;
    assign weights1[38][496] = 16'b1111111111111001;
    assign weights1[38][497] = 16'b1111111111110001;
    assign weights1[38][498] = 16'b1111111111111110;
    assign weights1[38][499] = 16'b0000000000001010;
    assign weights1[38][500] = 16'b0000000000001011;
    assign weights1[38][501] = 16'b0000000000010000;
    assign weights1[38][502] = 16'b0000000000000011;
    assign weights1[38][503] = 16'b0000000000000000;
    assign weights1[38][504] = 16'b1111111111111111;
    assign weights1[38][505] = 16'b0000000000000001;
    assign weights1[38][506] = 16'b1111111111111111;
    assign weights1[38][507] = 16'b1111111111111101;
    assign weights1[38][508] = 16'b0000000000000011;
    assign weights1[38][509] = 16'b0000000000000010;
    assign weights1[38][510] = 16'b1111111111111100;
    assign weights1[38][511] = 16'b1111111111110101;
    assign weights1[38][512] = 16'b1111111111110010;
    assign weights1[38][513] = 16'b1111111111101010;
    assign weights1[38][514] = 16'b1111111111100010;
    assign weights1[38][515] = 16'b1111111111100000;
    assign weights1[38][516] = 16'b1111111111010100;
    assign weights1[38][517] = 16'b1111111111001011;
    assign weights1[38][518] = 16'b1111111111101010;
    assign weights1[38][519] = 16'b0000000000001010;
    assign weights1[38][520] = 16'b0000000000010010;
    assign weights1[38][521] = 16'b0000000000010011;
    assign weights1[38][522] = 16'b0000000000000110;
    assign weights1[38][523] = 16'b0000000000000010;
    assign weights1[38][524] = 16'b1111111111111011;
    assign weights1[38][525] = 16'b0000000000000100;
    assign weights1[38][526] = 16'b0000000000011000;
    assign weights1[38][527] = 16'b0000000000010001;
    assign weights1[38][528] = 16'b0000000000010110;
    assign weights1[38][529] = 16'b0000000000001101;
    assign weights1[38][530] = 16'b0000000000001000;
    assign weights1[38][531] = 16'b0000000000000000;
    assign weights1[38][532] = 16'b1111111111111110;
    assign weights1[38][533] = 16'b0000000000000001;
    assign weights1[38][534] = 16'b1111111111111011;
    assign weights1[38][535] = 16'b1111111111111100;
    assign weights1[38][536] = 16'b0000000000000001;
    assign weights1[38][537] = 16'b1111111111110100;
    assign weights1[38][538] = 16'b1111111111110110;
    assign weights1[38][539] = 16'b1111111111101110;
    assign weights1[38][540] = 16'b1111111111100111;
    assign weights1[38][541] = 16'b1111111111011111;
    assign weights1[38][542] = 16'b1111111111010011;
    assign weights1[38][543] = 16'b1111111111011000;
    assign weights1[38][544] = 16'b1111111111011011;
    assign weights1[38][545] = 16'b1111111111011111;
    assign weights1[38][546] = 16'b1111111111110001;
    assign weights1[38][547] = 16'b1111111111111111;
    assign weights1[38][548] = 16'b0000000000010100;
    assign weights1[38][549] = 16'b0000000000010010;
    assign weights1[38][550] = 16'b0000000000001010;
    assign weights1[38][551] = 16'b1111111111111101;
    assign weights1[38][552] = 16'b0000000000000011;
    assign weights1[38][553] = 16'b0000000000000101;
    assign weights1[38][554] = 16'b0000000000011001;
    assign weights1[38][555] = 16'b0000000000010010;
    assign weights1[38][556] = 16'b0000000000010101;
    assign weights1[38][557] = 16'b0000000000010000;
    assign weights1[38][558] = 16'b0000000000001100;
    assign weights1[38][559] = 16'b0000000000000011;
    assign weights1[38][560] = 16'b1111111111111100;
    assign weights1[38][561] = 16'b1111111111111110;
    assign weights1[38][562] = 16'b1111111111111011;
    assign weights1[38][563] = 16'b1111111111111000;
    assign weights1[38][564] = 16'b1111111111111101;
    assign weights1[38][565] = 16'b1111111111101111;
    assign weights1[38][566] = 16'b1111111111110001;
    assign weights1[38][567] = 16'b1111111111110100;
    assign weights1[38][568] = 16'b1111111111100110;
    assign weights1[38][569] = 16'b1111111111011010;
    assign weights1[38][570] = 16'b1111111111010101;
    assign weights1[38][571] = 16'b1111111111001111;
    assign weights1[38][572] = 16'b1111111111100111;
    assign weights1[38][573] = 16'b1111111111101001;
    assign weights1[38][574] = 16'b1111111111111100;
    assign weights1[38][575] = 16'b0000000000000011;
    assign weights1[38][576] = 16'b0000000000010011;
    assign weights1[38][577] = 16'b0000000000010001;
    assign weights1[38][578] = 16'b0000000000001101;
    assign weights1[38][579] = 16'b0000000000001000;
    assign weights1[38][580] = 16'b0000000000001110;
    assign weights1[38][581] = 16'b0000000000001000;
    assign weights1[38][582] = 16'b0000000000010010;
    assign weights1[38][583] = 16'b0000000000010110;
    assign weights1[38][584] = 16'b0000000000001101;
    assign weights1[38][585] = 16'b0000000000000100;
    assign weights1[38][586] = 16'b0000000000001001;
    assign weights1[38][587] = 16'b0000000000000110;
    assign weights1[38][588] = 16'b1111111111111111;
    assign weights1[38][589] = 16'b1111111111111110;
    assign weights1[38][590] = 16'b1111111111111001;
    assign weights1[38][591] = 16'b1111111111111010;
    assign weights1[38][592] = 16'b1111111111110110;
    assign weights1[38][593] = 16'b1111111111111001;
    assign weights1[38][594] = 16'b1111111111110110;
    assign weights1[38][595] = 16'b1111111111110100;
    assign weights1[38][596] = 16'b1111111111101101;
    assign weights1[38][597] = 16'b1111111111100110;
    assign weights1[38][598] = 16'b1111111111011001;
    assign weights1[38][599] = 16'b1111111111010110;
    assign weights1[38][600] = 16'b1111111111100000;
    assign weights1[38][601] = 16'b1111111111111001;
    assign weights1[38][602] = 16'b0000000000001000;
    assign weights1[38][603] = 16'b0000000000010000;
    assign weights1[38][604] = 16'b0000000000010011;
    assign weights1[38][605] = 16'b0000000000011001;
    assign weights1[38][606] = 16'b0000000000000111;
    assign weights1[38][607] = 16'b0000000000000111;
    assign weights1[38][608] = 16'b0000000000001110;
    assign weights1[38][609] = 16'b0000000000001011;
    assign weights1[38][610] = 16'b0000000000001110;
    assign weights1[38][611] = 16'b0000000000001000;
    assign weights1[38][612] = 16'b0000000000001101;
    assign weights1[38][613] = 16'b1111111111111100;
    assign weights1[38][614] = 16'b0000000000000010;
    assign weights1[38][615] = 16'b1111111111111111;
    assign weights1[38][616] = 16'b1111111111111110;
    assign weights1[38][617] = 16'b1111111111111101;
    assign weights1[38][618] = 16'b1111111111111000;
    assign weights1[38][619] = 16'b1111111111110101;
    assign weights1[38][620] = 16'b1111111111110011;
    assign weights1[38][621] = 16'b1111111111110011;
    assign weights1[38][622] = 16'b1111111111111001;
    assign weights1[38][623] = 16'b1111111111110110;
    assign weights1[38][624] = 16'b1111111111110010;
    assign weights1[38][625] = 16'b1111111111110000;
    assign weights1[38][626] = 16'b1111111111101110;
    assign weights1[38][627] = 16'b1111111111111011;
    assign weights1[38][628] = 16'b1111111111111011;
    assign weights1[38][629] = 16'b0000000000000001;
    assign weights1[38][630] = 16'b0000000000000101;
    assign weights1[38][631] = 16'b0000000000010001;
    assign weights1[38][632] = 16'b0000000000001110;
    assign weights1[38][633] = 16'b0000000000011011;
    assign weights1[38][634] = 16'b0000000000010001;
    assign weights1[38][635] = 16'b0000000000000110;
    assign weights1[38][636] = 16'b0000000000001010;
    assign weights1[38][637] = 16'b0000000000001011;
    assign weights1[38][638] = 16'b0000000000010000;
    assign weights1[38][639] = 16'b0000000000001100;
    assign weights1[38][640] = 16'b0000000000001101;
    assign weights1[38][641] = 16'b0000000000000111;
    assign weights1[38][642] = 16'b0000000000000011;
    assign weights1[38][643] = 16'b0000000000000001;
    assign weights1[38][644] = 16'b1111111111111110;
    assign weights1[38][645] = 16'b1111111111111110;
    assign weights1[38][646] = 16'b1111111111111001;
    assign weights1[38][647] = 16'b1111111111110110;
    assign weights1[38][648] = 16'b1111111111101110;
    assign weights1[38][649] = 16'b1111111111110011;
    assign weights1[38][650] = 16'b1111111111101110;
    assign weights1[38][651] = 16'b1111111111110001;
    assign weights1[38][652] = 16'b1111111111110000;
    assign weights1[38][653] = 16'b1111111111110000;
    assign weights1[38][654] = 16'b0000000000000001;
    assign weights1[38][655] = 16'b0000000000000101;
    assign weights1[38][656] = 16'b0000000000001010;
    assign weights1[38][657] = 16'b1111111111111110;
    assign weights1[38][658] = 16'b1111111111111000;
    assign weights1[38][659] = 16'b0000000000001100;
    assign weights1[38][660] = 16'b0000000000000000;
    assign weights1[38][661] = 16'b0000000000000111;
    assign weights1[38][662] = 16'b0000000000010100;
    assign weights1[38][663] = 16'b0000000000000010;
    assign weights1[38][664] = 16'b0000000000000111;
    assign weights1[38][665] = 16'b0000000000000111;
    assign weights1[38][666] = 16'b0000000000001010;
    assign weights1[38][667] = 16'b0000000000001001;
    assign weights1[38][668] = 16'b0000000000000001;
    assign weights1[38][669] = 16'b0000000000000011;
    assign weights1[38][670] = 16'b0000000000000011;
    assign weights1[38][671] = 16'b0000000000000010;
    assign weights1[38][672] = 16'b1111111111111111;
    assign weights1[38][673] = 16'b1111111111111110;
    assign weights1[38][674] = 16'b1111111111111001;
    assign weights1[38][675] = 16'b1111111111111000;
    assign weights1[38][676] = 16'b1111111111101111;
    assign weights1[38][677] = 16'b1111111111110001;
    assign weights1[38][678] = 16'b1111111111110001;
    assign weights1[38][679] = 16'b1111111111111000;
    assign weights1[38][680] = 16'b1111111111101110;
    assign weights1[38][681] = 16'b1111111111110110;
    assign weights1[38][682] = 16'b0000000000000000;
    assign weights1[38][683] = 16'b0000000000000011;
    assign weights1[38][684] = 16'b0000000000001011;
    assign weights1[38][685] = 16'b0000000000000111;
    assign weights1[38][686] = 16'b0000000000000001;
    assign weights1[38][687] = 16'b0000000000000011;
    assign weights1[38][688] = 16'b0000000000010010;
    assign weights1[38][689] = 16'b0000000000001100;
    assign weights1[38][690] = 16'b0000000000001011;
    assign weights1[38][691] = 16'b0000000000000001;
    assign weights1[38][692] = 16'b0000000000000111;
    assign weights1[38][693] = 16'b0000000000000100;
    assign weights1[38][694] = 16'b0000000000000110;
    assign weights1[38][695] = 16'b0000000000000110;
    assign weights1[38][696] = 16'b0000000000000011;
    assign weights1[38][697] = 16'b1111111111111111;
    assign weights1[38][698] = 16'b1111111111111101;
    assign weights1[38][699] = 16'b0000000000000001;
    assign weights1[38][700] = 16'b1111111111111111;
    assign weights1[38][701] = 16'b1111111111111110;
    assign weights1[38][702] = 16'b1111111111111100;
    assign weights1[38][703] = 16'b1111111111111110;
    assign weights1[38][704] = 16'b1111111111110100;
    assign weights1[38][705] = 16'b1111111111101101;
    assign weights1[38][706] = 16'b1111111111101111;
    assign weights1[38][707] = 16'b1111111111110101;
    assign weights1[38][708] = 16'b1111111111111001;
    assign weights1[38][709] = 16'b0000000000000100;
    assign weights1[38][710] = 16'b0000000000001010;
    assign weights1[38][711] = 16'b0000000000001101;
    assign weights1[38][712] = 16'b1111111111111010;
    assign weights1[38][713] = 16'b1111111111111110;
    assign weights1[38][714] = 16'b1111111111111101;
    assign weights1[38][715] = 16'b1111111111111110;
    assign weights1[38][716] = 16'b0000000000001011;
    assign weights1[38][717] = 16'b0000000000010010;
    assign weights1[38][718] = 16'b0000000000000110;
    assign weights1[38][719] = 16'b0000000000001000;
    assign weights1[38][720] = 16'b0000000000001101;
    assign weights1[38][721] = 16'b0000000000010000;
    assign weights1[38][722] = 16'b0000000000001010;
    assign weights1[38][723] = 16'b0000000000000100;
    assign weights1[38][724] = 16'b0000000000000010;
    assign weights1[38][725] = 16'b0000000000000000;
    assign weights1[38][726] = 16'b1111111111111111;
    assign weights1[38][727] = 16'b1111111111111111;
    assign weights1[38][728] = 16'b1111111111111101;
    assign weights1[38][729] = 16'b1111111111111101;
    assign weights1[38][730] = 16'b1111111111111111;
    assign weights1[38][731] = 16'b1111111111111110;
    assign weights1[38][732] = 16'b1111111111111001;
    assign weights1[38][733] = 16'b1111111111110101;
    assign weights1[38][734] = 16'b1111111111110101;
    assign weights1[38][735] = 16'b1111111111111001;
    assign weights1[38][736] = 16'b1111111111111100;
    assign weights1[38][737] = 16'b0000000000000111;
    assign weights1[38][738] = 16'b0000000000001011;
    assign weights1[38][739] = 16'b0000000000001001;
    assign weights1[38][740] = 16'b0000000000000001;
    assign weights1[38][741] = 16'b1111111111111110;
    assign weights1[38][742] = 16'b0000000000000110;
    assign weights1[38][743] = 16'b0000000000010001;
    assign weights1[38][744] = 16'b0000000000001101;
    assign weights1[38][745] = 16'b0000000000001000;
    assign weights1[38][746] = 16'b1111111111111010;
    assign weights1[38][747] = 16'b0000000000000000;
    assign weights1[38][748] = 16'b0000000000000110;
    assign weights1[38][749] = 16'b0000000000001101;
    assign weights1[38][750] = 16'b0000000000001001;
    assign weights1[38][751] = 16'b1111111111111111;
    assign weights1[38][752] = 16'b0000000000000000;
    assign weights1[38][753] = 16'b1111111111111111;
    assign weights1[38][754] = 16'b1111111111111111;
    assign weights1[38][755] = 16'b0000000000000000;
    assign weights1[38][756] = 16'b1111111111111110;
    assign weights1[38][757] = 16'b1111111111111110;
    assign weights1[38][758] = 16'b1111111111111110;
    assign weights1[38][759] = 16'b1111111111111111;
    assign weights1[38][760] = 16'b1111111111111101;
    assign weights1[38][761] = 16'b1111111111111101;
    assign weights1[38][762] = 16'b1111111111111110;
    assign weights1[38][763] = 16'b0000000000000101;
    assign weights1[38][764] = 16'b0000000000000100;
    assign weights1[38][765] = 16'b0000000000000110;
    assign weights1[38][766] = 16'b0000000000001000;
    assign weights1[38][767] = 16'b0000000000001111;
    assign weights1[38][768] = 16'b0000000000001100;
    assign weights1[38][769] = 16'b0000000000001010;
    assign weights1[38][770] = 16'b0000000000001011;
    assign weights1[38][771] = 16'b0000000000001010;
    assign weights1[38][772] = 16'b0000000000011010;
    assign weights1[38][773] = 16'b0000000000001111;
    assign weights1[38][774] = 16'b0000000000001001;
    assign weights1[38][775] = 16'b0000000000010010;
    assign weights1[38][776] = 16'b0000000000001000;
    assign weights1[38][777] = 16'b0000000000001001;
    assign weights1[38][778] = 16'b0000000000000100;
    assign weights1[38][779] = 16'b0000000000000011;
    assign weights1[38][780] = 16'b0000000000000010;
    assign weights1[38][781] = 16'b1111111111111111;
    assign weights1[38][782] = 16'b1111111111111111;
    assign weights1[38][783] = 16'b0000000000000000;
    assign weights1[39][0] = 16'b0000000000000001;
    assign weights1[39][1] = 16'b0000000000000001;
    assign weights1[39][2] = 16'b0000000000000001;
    assign weights1[39][3] = 16'b0000000000000000;
    assign weights1[39][4] = 16'b1111111111111101;
    assign weights1[39][5] = 16'b1111111111110111;
    assign weights1[39][6] = 16'b1111111111110110;
    assign weights1[39][7] = 16'b1111111111101110;
    assign weights1[39][8] = 16'b1111111111101011;
    assign weights1[39][9] = 16'b1111111111111101;
    assign weights1[39][10] = 16'b0000000000000001;
    assign weights1[39][11] = 16'b1111111111110101;
    assign weights1[39][12] = 16'b1111111111110101;
    assign weights1[39][13] = 16'b1111111111111111;
    assign weights1[39][14] = 16'b1111111111110110;
    assign weights1[39][15] = 16'b1111111111110000;
    assign weights1[39][16] = 16'b1111111111110000;
    assign weights1[39][17] = 16'b1111111111110011;
    assign weights1[39][18] = 16'b1111111111111101;
    assign weights1[39][19] = 16'b1111111111111111;
    assign weights1[39][20] = 16'b1111111111110110;
    assign weights1[39][21] = 16'b0000000000000101;
    assign weights1[39][22] = 16'b1111111111111111;
    assign weights1[39][23] = 16'b0000000000001101;
    assign weights1[39][24] = 16'b0000000000001000;
    assign weights1[39][25] = 16'b0000000000001000;
    assign weights1[39][26] = 16'b0000000000001000;
    assign weights1[39][27] = 16'b1111111111111110;
    assign weights1[39][28] = 16'b0000000000000001;
    assign weights1[39][29] = 16'b0000000000000000;
    assign weights1[39][30] = 16'b0000000000000000;
    assign weights1[39][31] = 16'b1111111111111111;
    assign weights1[39][32] = 16'b1111111111111101;
    assign weights1[39][33] = 16'b1111111111111111;
    assign weights1[39][34] = 16'b1111111111111100;
    assign weights1[39][35] = 16'b1111111111111110;
    assign weights1[39][36] = 16'b0000000000000011;
    assign weights1[39][37] = 16'b1111111111111001;
    assign weights1[39][38] = 16'b1111111111111100;
    assign weights1[39][39] = 16'b1111111111101110;
    assign weights1[39][40] = 16'b1111111111111011;
    assign weights1[39][41] = 16'b1111111111110100;
    assign weights1[39][42] = 16'b1111111111111001;
    assign weights1[39][43] = 16'b1111111111110111;
    assign weights1[39][44] = 16'b1111111111110001;
    assign weights1[39][45] = 16'b1111111111110001;
    assign weights1[39][46] = 16'b1111111111110001;
    assign weights1[39][47] = 16'b0000000000001001;
    assign weights1[39][48] = 16'b1111111111110001;
    assign weights1[39][49] = 16'b1111111111110100;
    assign weights1[39][50] = 16'b0000000000000110;
    assign weights1[39][51] = 16'b1111111111111101;
    assign weights1[39][52] = 16'b0000000000000101;
    assign weights1[39][53] = 16'b0000000000010000;
    assign weights1[39][54] = 16'b0000000000001101;
    assign weights1[39][55] = 16'b0000000000000110;
    assign weights1[39][56] = 16'b0000000000000011;
    assign weights1[39][57] = 16'b0000000000000011;
    assign weights1[39][58] = 16'b0000000000000111;
    assign weights1[39][59] = 16'b0000000000000001;
    assign weights1[39][60] = 16'b0000000000000011;
    assign weights1[39][61] = 16'b1111111111111111;
    assign weights1[39][62] = 16'b0000000000000010;
    assign weights1[39][63] = 16'b0000000000000011;
    assign weights1[39][64] = 16'b1111111111110010;
    assign weights1[39][65] = 16'b1111111111111110;
    assign weights1[39][66] = 16'b0000000000000111;
    assign weights1[39][67] = 16'b1111111111111111;
    assign weights1[39][68] = 16'b0000000000000001;
    assign weights1[39][69] = 16'b1111111111111011;
    assign weights1[39][70] = 16'b1111111111111000;
    assign weights1[39][71] = 16'b0000000000000100;
    assign weights1[39][72] = 16'b0000000000000010;
    assign weights1[39][73] = 16'b0000000000000100;
    assign weights1[39][74] = 16'b0000000000001011;
    assign weights1[39][75] = 16'b0000000000000111;
    assign weights1[39][76] = 16'b0000000000001100;
    assign weights1[39][77] = 16'b0000000000000111;
    assign weights1[39][78] = 16'b1111111111111010;
    assign weights1[39][79] = 16'b0000000000000111;
    assign weights1[39][80] = 16'b0000000000010010;
    assign weights1[39][81] = 16'b0000000000001111;
    assign weights1[39][82] = 16'b0000000000010010;
    assign weights1[39][83] = 16'b0000000000001100;
    assign weights1[39][84] = 16'b0000000000001001;
    assign weights1[39][85] = 16'b0000000000000101;
    assign weights1[39][86] = 16'b0000000000000110;
    assign weights1[39][87] = 16'b0000000000001010;
    assign weights1[39][88] = 16'b0000000000000011;
    assign weights1[39][89] = 16'b0000000000001010;
    assign weights1[39][90] = 16'b0000000000000000;
    assign weights1[39][91] = 16'b0000000000000010;
    assign weights1[39][92] = 16'b0000000000000101;
    assign weights1[39][93] = 16'b0000000000010001;
    assign weights1[39][94] = 16'b1111111111111000;
    assign weights1[39][95] = 16'b0000000000001011;
    assign weights1[39][96] = 16'b1111111111111001;
    assign weights1[39][97] = 16'b1111111111111101;
    assign weights1[39][98] = 16'b0000000000000001;
    assign weights1[39][99] = 16'b1111111111110101;
    assign weights1[39][100] = 16'b0000000000000001;
    assign weights1[39][101] = 16'b1111111111110000;
    assign weights1[39][102] = 16'b1111111111110110;
    assign weights1[39][103] = 16'b1111111111111010;
    assign weights1[39][104] = 16'b0000000000000000;
    assign weights1[39][105] = 16'b0000000000000101;
    assign weights1[39][106] = 16'b0000000000000111;
    assign weights1[39][107] = 16'b0000000000001101;
    assign weights1[39][108] = 16'b0000000000010111;
    assign weights1[39][109] = 16'b0000000000000010;
    assign weights1[39][110] = 16'b0000000000010000;
    assign weights1[39][111] = 16'b0000000000001001;
    assign weights1[39][112] = 16'b0000000000001100;
    assign weights1[39][113] = 16'b0000000000000101;
    assign weights1[39][114] = 16'b0000000000010000;
    assign weights1[39][115] = 16'b0000000000010100;
    assign weights1[39][116] = 16'b0000000000100000;
    assign weights1[39][117] = 16'b0000000000010101;
    assign weights1[39][118] = 16'b0000000000000010;
    assign weights1[39][119] = 16'b0000000000000001;
    assign weights1[39][120] = 16'b1111111111110001;
    assign weights1[39][121] = 16'b1111111111111010;
    assign weights1[39][122] = 16'b1111111111100111;
    assign weights1[39][123] = 16'b1111111111111001;
    assign weights1[39][124] = 16'b0000000000001100;
    assign weights1[39][125] = 16'b0000000000000011;
    assign weights1[39][126] = 16'b1111111111111110;
    assign weights1[39][127] = 16'b1111111111111110;
    assign weights1[39][128] = 16'b0000000000001001;
    assign weights1[39][129] = 16'b0000000000011001;
    assign weights1[39][130] = 16'b0000000000010001;
    assign weights1[39][131] = 16'b0000000000010100;
    assign weights1[39][132] = 16'b1111111111111011;
    assign weights1[39][133] = 16'b0000000000000101;
    assign weights1[39][134] = 16'b1111111111111110;
    assign weights1[39][135] = 16'b1111111111110110;
    assign weights1[39][136] = 16'b1111111111111111;
    assign weights1[39][137] = 16'b0000000000010011;
    assign weights1[39][138] = 16'b0000000000001010;
    assign weights1[39][139] = 16'b0000000000001101;
    assign weights1[39][140] = 16'b0000000000010100;
    assign weights1[39][141] = 16'b0000000000010100;
    assign weights1[39][142] = 16'b0000000000010010;
    assign weights1[39][143] = 16'b0000000000011011;
    assign weights1[39][144] = 16'b0000000000011011;
    assign weights1[39][145] = 16'b0000000000011001;
    assign weights1[39][146] = 16'b0000000000001001;
    assign weights1[39][147] = 16'b0000000000011001;
    assign weights1[39][148] = 16'b0000000000000011;
    assign weights1[39][149] = 16'b1111111111111101;
    assign weights1[39][150] = 16'b0000000000000000;
    assign weights1[39][151] = 16'b0000000000001010;
    assign weights1[39][152] = 16'b1111111111111111;
    assign weights1[39][153] = 16'b0000000000001001;
    assign weights1[39][154] = 16'b1111111111111101;
    assign weights1[39][155] = 16'b0000000000010111;
    assign weights1[39][156] = 16'b0000000000001001;
    assign weights1[39][157] = 16'b0000000000011011;
    assign weights1[39][158] = 16'b0000000000010101;
    assign weights1[39][159] = 16'b0000000000000100;
    assign weights1[39][160] = 16'b0000000000001110;
    assign weights1[39][161] = 16'b0000000000001011;
    assign weights1[39][162] = 16'b0000000000010000;
    assign weights1[39][163] = 16'b0000000000000011;
    assign weights1[39][164] = 16'b0000000000001010;
    assign weights1[39][165] = 16'b0000000000001101;
    assign weights1[39][166] = 16'b0000000000011101;
    assign weights1[39][167] = 16'b0000000000010101;
    assign weights1[39][168] = 16'b0000000000010010;
    assign weights1[39][169] = 16'b0000000000010001;
    assign weights1[39][170] = 16'b0000000000010101;
    assign weights1[39][171] = 16'b0000000000101010;
    assign weights1[39][172] = 16'b0000000000101010;
    assign weights1[39][173] = 16'b0000000000101100;
    assign weights1[39][174] = 16'b0000000000101001;
    assign weights1[39][175] = 16'b0000000000011011;
    assign weights1[39][176] = 16'b0000000000011010;
    assign weights1[39][177] = 16'b0000000000010101;
    assign weights1[39][178] = 16'b0000000000001000;
    assign weights1[39][179] = 16'b0000000000000111;
    assign weights1[39][180] = 16'b0000000000001000;
    assign weights1[39][181] = 16'b0000000000001100;
    assign weights1[39][182] = 16'b0000000000001111;
    assign weights1[39][183] = 16'b0000000000001011;
    assign weights1[39][184] = 16'b0000000000001110;
    assign weights1[39][185] = 16'b0000000000001000;
    assign weights1[39][186] = 16'b0000000000010101;
    assign weights1[39][187] = 16'b0000000000000101;
    assign weights1[39][188] = 16'b1111111111110010;
    assign weights1[39][189] = 16'b0000000000001111;
    assign weights1[39][190] = 16'b0000000000010101;
    assign weights1[39][191] = 16'b0000000000001111;
    assign weights1[39][192] = 16'b0000000000011000;
    assign weights1[39][193] = 16'b0000000000000100;
    assign weights1[39][194] = 16'b0000000000010101;
    assign weights1[39][195] = 16'b0000000000011100;
    assign weights1[39][196] = 16'b0000000000001100;
    assign weights1[39][197] = 16'b0000000000001100;
    assign weights1[39][198] = 16'b0000000000010011;
    assign weights1[39][199] = 16'b0000000000101111;
    assign weights1[39][200] = 16'b0000000000000000;
    assign weights1[39][201] = 16'b0000000000001111;
    assign weights1[39][202] = 16'b0000000000010101;
    assign weights1[39][203] = 16'b0000000001001001;
    assign weights1[39][204] = 16'b0000000000001110;
    assign weights1[39][205] = 16'b0000000000100010;
    assign weights1[39][206] = 16'b0000000000100011;
    assign weights1[39][207] = 16'b0000000000001111;
    assign weights1[39][208] = 16'b0000000000010111;
    assign weights1[39][209] = 16'b0000000000010111;
    assign weights1[39][210] = 16'b0000000000010110;
    assign weights1[39][211] = 16'b0000000000010011;
    assign weights1[39][212] = 16'b0000000000011001;
    assign weights1[39][213] = 16'b0000000000000010;
    assign weights1[39][214] = 16'b0000000000001101;
    assign weights1[39][215] = 16'b0000000000011001;
    assign weights1[39][216] = 16'b0000000000011001;
    assign weights1[39][217] = 16'b0000000000011001;
    assign weights1[39][218] = 16'b0000000000000001;
    assign weights1[39][219] = 16'b0000000000010000;
    assign weights1[39][220] = 16'b0000000000010011;
    assign weights1[39][221] = 16'b0000000000001100;
    assign weights1[39][222] = 16'b1111111111111010;
    assign weights1[39][223] = 16'b0000000000100000;
    assign weights1[39][224] = 16'b0000000000010010;
    assign weights1[39][225] = 16'b0000000000011011;
    assign weights1[39][226] = 16'b0000000000011011;
    assign weights1[39][227] = 16'b0000000000100100;
    assign weights1[39][228] = 16'b0000000000100111;
    assign weights1[39][229] = 16'b0000000000011100;
    assign weights1[39][230] = 16'b0000000000010110;
    assign weights1[39][231] = 16'b0000000000100111;
    assign weights1[39][232] = 16'b0000000000100101;
    assign weights1[39][233] = 16'b0000000000101000;
    assign weights1[39][234] = 16'b0000000000011010;
    assign weights1[39][235] = 16'b0000000000110101;
    assign weights1[39][236] = 16'b0000000000001010;
    assign weights1[39][237] = 16'b0000000000011110;
    assign weights1[39][238] = 16'b0000000000010100;
    assign weights1[39][239] = 16'b0000000000100110;
    assign weights1[39][240] = 16'b0000000000001011;
    assign weights1[39][241] = 16'b0000000000001011;
    assign weights1[39][242] = 16'b0000000000001001;
    assign weights1[39][243] = 16'b0000000000001011;
    assign weights1[39][244] = 16'b0000000000001011;
    assign weights1[39][245] = 16'b0000000000011100;
    assign weights1[39][246] = 16'b0000000000000110;
    assign weights1[39][247] = 16'b0000000000000001;
    assign weights1[39][248] = 16'b0000000000010101;
    assign weights1[39][249] = 16'b0000000000000011;
    assign weights1[39][250] = 16'b0000000000001010;
    assign weights1[39][251] = 16'b0000000000010000;
    assign weights1[39][252] = 16'b0000000000001100;
    assign weights1[39][253] = 16'b0000000000011000;
    assign weights1[39][254] = 16'b0000000000100101;
    assign weights1[39][255] = 16'b0000000000011111;
    assign weights1[39][256] = 16'b0000000000101100;
    assign weights1[39][257] = 16'b0000000000011111;
    assign weights1[39][258] = 16'b0000000000100110;
    assign weights1[39][259] = 16'b0000000000010111;
    assign weights1[39][260] = 16'b0000000000100100;
    assign weights1[39][261] = 16'b0000000000011000;
    assign weights1[39][262] = 16'b0000000000011100;
    assign weights1[39][263] = 16'b0000000000101001;
    assign weights1[39][264] = 16'b0000000000011101;
    assign weights1[39][265] = 16'b0000000000011001;
    assign weights1[39][266] = 16'b0000000000011001;
    assign weights1[39][267] = 16'b0000000000001101;
    assign weights1[39][268] = 16'b0000000000100100;
    assign weights1[39][269] = 16'b0000000000101101;
    assign weights1[39][270] = 16'b0000000000001111;
    assign weights1[39][271] = 16'b0000000000001110;
    assign weights1[39][272] = 16'b0000000000001011;
    assign weights1[39][273] = 16'b1111111111111110;
    assign weights1[39][274] = 16'b0000000000011001;
    assign weights1[39][275] = 16'b0000000000000100;
    assign weights1[39][276] = 16'b0000000000001101;
    assign weights1[39][277] = 16'b0000000000010001;
    assign weights1[39][278] = 16'b0000000000001111;
    assign weights1[39][279] = 16'b0000000000001101;
    assign weights1[39][280] = 16'b0000000000001110;
    assign weights1[39][281] = 16'b0000000000011000;
    assign weights1[39][282] = 16'b0000000000101010;
    assign weights1[39][283] = 16'b0000000000100101;
    assign weights1[39][284] = 16'b0000000000010100;
    assign weights1[39][285] = 16'b0000000000101100;
    assign weights1[39][286] = 16'b0000000000010011;
    assign weights1[39][287] = 16'b0000000000011011;
    assign weights1[39][288] = 16'b0000000000100111;
    assign weights1[39][289] = 16'b0000000000011110;
    assign weights1[39][290] = 16'b0000000000101001;
    assign weights1[39][291] = 16'b0000000000011000;
    assign weights1[39][292] = 16'b0000000000011010;
    assign weights1[39][293] = 16'b0000000000010001;
    assign weights1[39][294] = 16'b0000000000100011;
    assign weights1[39][295] = 16'b0000000000110111;
    assign weights1[39][296] = 16'b0000000000010000;
    assign weights1[39][297] = 16'b0000000000110001;
    assign weights1[39][298] = 16'b0000000000011000;
    assign weights1[39][299] = 16'b0000000000110100;
    assign weights1[39][300] = 16'b0000000000010101;
    assign weights1[39][301] = 16'b0000000000011000;
    assign weights1[39][302] = 16'b0000000000010011;
    assign weights1[39][303] = 16'b0000000000000110;
    assign weights1[39][304] = 16'b1111111111111110;
    assign weights1[39][305] = 16'b0000000000100110;
    assign weights1[39][306] = 16'b0000000000011010;
    assign weights1[39][307] = 16'b0000000000000101;
    assign weights1[39][308] = 16'b0000000000001010;
    assign weights1[39][309] = 16'b0000000000001110;
    assign weights1[39][310] = 16'b0000000000010101;
    assign weights1[39][311] = 16'b0000000000011111;
    assign weights1[39][312] = 16'b0000000000100001;
    assign weights1[39][313] = 16'b0000000000011100;
    assign weights1[39][314] = 16'b0000000000101001;
    assign weights1[39][315] = 16'b0000000000110010;
    assign weights1[39][316] = 16'b0000000000100001;
    assign weights1[39][317] = 16'b0000000000001001;
    assign weights1[39][318] = 16'b0000000000011011;
    assign weights1[39][319] = 16'b0000000000100100;
    assign weights1[39][320] = 16'b0000000000010101;
    assign weights1[39][321] = 16'b0000000000011001;
    assign weights1[39][322] = 16'b0000000000101001;
    assign weights1[39][323] = 16'b0000000000101001;
    assign weights1[39][324] = 16'b0000000000011010;
    assign weights1[39][325] = 16'b0000000000100010;
    assign weights1[39][326] = 16'b0000000000011111;
    assign weights1[39][327] = 16'b0000000000101100;
    assign weights1[39][328] = 16'b0000000000100001;
    assign weights1[39][329] = 16'b0000000000100110;
    assign weights1[39][330] = 16'b0000000000111011;
    assign weights1[39][331] = 16'b0000000000111001;
    assign weights1[39][332] = 16'b0000000000110111;
    assign weights1[39][333] = 16'b0000000000100011;
    assign weights1[39][334] = 16'b0000000000101100;
    assign weights1[39][335] = 16'b0000000000011010;
    assign weights1[39][336] = 16'b1111111111111101;
    assign weights1[39][337] = 16'b1111111111110000;
    assign weights1[39][338] = 16'b0000000000001110;
    assign weights1[39][339] = 16'b0000000000011010;
    assign weights1[39][340] = 16'b0000000000100111;
    assign weights1[39][341] = 16'b0000000000101000;
    assign weights1[39][342] = 16'b0000000000001000;
    assign weights1[39][343] = 16'b0000000000010010;
    assign weights1[39][344] = 16'b0000000000110000;
    assign weights1[39][345] = 16'b0000000000010001;
    assign weights1[39][346] = 16'b0000000000011101;
    assign weights1[39][347] = 16'b0000000000101110;
    assign weights1[39][348] = 16'b0000000000011111;
    assign weights1[39][349] = 16'b0000000000011010;
    assign weights1[39][350] = 16'b0000000000011000;
    assign weights1[39][351] = 16'b0000000000001100;
    assign weights1[39][352] = 16'b0000000000100100;
    assign weights1[39][353] = 16'b0000000000011110;
    assign weights1[39][354] = 16'b0000000000100110;
    assign weights1[39][355] = 16'b0000000000101011;
    assign weights1[39][356] = 16'b0000000000101011;
    assign weights1[39][357] = 16'b0000000000110011;
    assign weights1[39][358] = 16'b0000000000110010;
    assign weights1[39][359] = 16'b0000000000100010;
    assign weights1[39][360] = 16'b0000000000111000;
    assign weights1[39][361] = 16'b0000000000100011;
    assign weights1[39][362] = 16'b0000000000100001;
    assign weights1[39][363] = 16'b0000000000001111;
    assign weights1[39][364] = 16'b1111111111110110;
    assign weights1[39][365] = 16'b1111111111100100;
    assign weights1[39][366] = 16'b1111111111110010;
    assign weights1[39][367] = 16'b0000000000011100;
    assign weights1[39][368] = 16'b0000000000101001;
    assign weights1[39][369] = 16'b0000000000010111;
    assign weights1[39][370] = 16'b0000000000001001;
    assign weights1[39][371] = 16'b0000000000010111;
    assign weights1[39][372] = 16'b0000000000011101;
    assign weights1[39][373] = 16'b0000000000001110;
    assign weights1[39][374] = 16'b0000000000010110;
    assign weights1[39][375] = 16'b1111111111111100;
    assign weights1[39][376] = 16'b0000000000011001;
    assign weights1[39][377] = 16'b0000000000010011;
    assign weights1[39][378] = 16'b1111111111111101;
    assign weights1[39][379] = 16'b0000000000001010;
    assign weights1[39][380] = 16'b1111111111111101;
    assign weights1[39][381] = 16'b0000000000001011;
    assign weights1[39][382] = 16'b0000000000001101;
    assign weights1[39][383] = 16'b0000000000011001;
    assign weights1[39][384] = 16'b0000000000011110;
    assign weights1[39][385] = 16'b0000000000001010;
    assign weights1[39][386] = 16'b0000000000001101;
    assign weights1[39][387] = 16'b0000000000100111;
    assign weights1[39][388] = 16'b0000000000100000;
    assign weights1[39][389] = 16'b0000000000010100;
    assign weights1[39][390] = 16'b0000000000011010;
    assign weights1[39][391] = 16'b0000000000000110;
    assign weights1[39][392] = 16'b1111111111100010;
    assign weights1[39][393] = 16'b1111111111011000;
    assign weights1[39][394] = 16'b1111111111010000;
    assign weights1[39][395] = 16'b1111111111011000;
    assign weights1[39][396] = 16'b1111111111101111;
    assign weights1[39][397] = 16'b1111111111100101;
    assign weights1[39][398] = 16'b1111111111101111;
    assign weights1[39][399] = 16'b1111111111111001;
    assign weights1[39][400] = 16'b1111111111111111;
    assign weights1[39][401] = 16'b1111111111011100;
    assign weights1[39][402] = 16'b1111111110110101;
    assign weights1[39][403] = 16'b1111111110111100;
    assign weights1[39][404] = 16'b1111111111000000;
    assign weights1[39][405] = 16'b1111111111001100;
    assign weights1[39][406] = 16'b1111111111010110;
    assign weights1[39][407] = 16'b1111111111011000;
    assign weights1[39][408] = 16'b1111111111110100;
    assign weights1[39][409] = 16'b1111111111100011;
    assign weights1[39][410] = 16'b1111111111011001;
    assign weights1[39][411] = 16'b1111111111111000;
    assign weights1[39][412] = 16'b0000000000000010;
    assign weights1[39][413] = 16'b0000000000000100;
    assign weights1[39][414] = 16'b1111111111110111;
    assign weights1[39][415] = 16'b0000000000000101;
    assign weights1[39][416] = 16'b1111111111110111;
    assign weights1[39][417] = 16'b0000000000000010;
    assign weights1[39][418] = 16'b0000000000000111;
    assign weights1[39][419] = 16'b0000000000001001;
    assign weights1[39][420] = 16'b1111111111010111;
    assign weights1[39][421] = 16'b1111111111001010;
    assign weights1[39][422] = 16'b1111111110110001;
    assign weights1[39][423] = 16'b1111111110101100;
    assign weights1[39][424] = 16'b1111111110111101;
    assign weights1[39][425] = 16'b1111111110110100;
    assign weights1[39][426] = 16'b1111111110110000;
    assign weights1[39][427] = 16'b1111111110110110;
    assign weights1[39][428] = 16'b1111111110000100;
    assign weights1[39][429] = 16'b1111111101110010;
    assign weights1[39][430] = 16'b1111111110001000;
    assign weights1[39][431] = 16'b1111111110000110;
    assign weights1[39][432] = 16'b1111111110001101;
    assign weights1[39][433] = 16'b1111111110001111;
    assign weights1[39][434] = 16'b1111111110001111;
    assign weights1[39][435] = 16'b1111111110101100;
    assign weights1[39][436] = 16'b1111111110110011;
    assign weights1[39][437] = 16'b1111111110111111;
    assign weights1[39][438] = 16'b1111111111001001;
    assign weights1[39][439] = 16'b1111111111000110;
    assign weights1[39][440] = 16'b1111111110111100;
    assign weights1[39][441] = 16'b1111111111011100;
    assign weights1[39][442] = 16'b1111111111010011;
    assign weights1[39][443] = 16'b1111111111101001;
    assign weights1[39][444] = 16'b1111111111011011;
    assign weights1[39][445] = 16'b1111111111111011;
    assign weights1[39][446] = 16'b1111111111111001;
    assign weights1[39][447] = 16'b1111111111111010;
    assign weights1[39][448] = 16'b1111111111011010;
    assign weights1[39][449] = 16'b1111111111001000;
    assign weights1[39][450] = 16'b1111111110111001;
    assign weights1[39][451] = 16'b1111111110110000;
    assign weights1[39][452] = 16'b1111111110011001;
    assign weights1[39][453] = 16'b1111111110000111;
    assign weights1[39][454] = 16'b1111111101111110;
    assign weights1[39][455] = 16'b1111111101100111;
    assign weights1[39][456] = 16'b1111111101110100;
    assign weights1[39][457] = 16'b1111111101111011;
    assign weights1[39][458] = 16'b1111111110101100;
    assign weights1[39][459] = 16'b1111111110110100;
    assign weights1[39][460] = 16'b1111111110110010;
    assign weights1[39][461] = 16'b1111111110111000;
    assign weights1[39][462] = 16'b1111111110111000;
    assign weights1[39][463] = 16'b1111111110101111;
    assign weights1[39][464] = 16'b1111111110111000;
    assign weights1[39][465] = 16'b1111111110111001;
    assign weights1[39][466] = 16'b1111111110111010;
    assign weights1[39][467] = 16'b1111111111001001;
    assign weights1[39][468] = 16'b1111111110101111;
    assign weights1[39][469] = 16'b1111111111010110;
    assign weights1[39][470] = 16'b1111111111010001;
    assign weights1[39][471] = 16'b1111111111001001;
    assign weights1[39][472] = 16'b1111111111011010;
    assign weights1[39][473] = 16'b1111111111111011;
    assign weights1[39][474] = 16'b1111111111101100;
    assign weights1[39][475] = 16'b1111111111110010;
    assign weights1[39][476] = 16'b1111111111011110;
    assign weights1[39][477] = 16'b1111111111000101;
    assign weights1[39][478] = 16'b1111111111000111;
    assign weights1[39][479] = 16'b1111111110110011;
    assign weights1[39][480] = 16'b1111111110011001;
    assign weights1[39][481] = 16'b1111111110010100;
    assign weights1[39][482] = 16'b1111111101110101;
    assign weights1[39][483] = 16'b1111111110011000;
    assign weights1[39][484] = 16'b1111111111001001;
    assign weights1[39][485] = 16'b1111111111101011;
    assign weights1[39][486] = 16'b1111111111101001;
    assign weights1[39][487] = 16'b1111111111101001;
    assign weights1[39][488] = 16'b1111111111110001;
    assign weights1[39][489] = 16'b1111111111100110;
    assign weights1[39][490] = 16'b1111111111100100;
    assign weights1[39][491] = 16'b1111111111011100;
    assign weights1[39][492] = 16'b1111111111011110;
    assign weights1[39][493] = 16'b1111111111100011;
    assign weights1[39][494] = 16'b1111111111011100;
    assign weights1[39][495] = 16'b1111111111010011;
    assign weights1[39][496] = 16'b1111111111011101;
    assign weights1[39][497] = 16'b1111111110111000;
    assign weights1[39][498] = 16'b1111111111100110;
    assign weights1[39][499] = 16'b1111111111010101;
    assign weights1[39][500] = 16'b1111111111101000;
    assign weights1[39][501] = 16'b1111111111101100;
    assign weights1[39][502] = 16'b1111111111100101;
    assign weights1[39][503] = 16'b1111111111101101;
    assign weights1[39][504] = 16'b1111111111100001;
    assign weights1[39][505] = 16'b1111111111010101;
    assign weights1[39][506] = 16'b1111111111001001;
    assign weights1[39][507] = 16'b1111111110110000;
    assign weights1[39][508] = 16'b1111111111001010;
    assign weights1[39][509] = 16'b1111111110111001;
    assign weights1[39][510] = 16'b1111111111011001;
    assign weights1[39][511] = 16'b1111111111011111;
    assign weights1[39][512] = 16'b1111111111111010;
    assign weights1[39][513] = 16'b0000000000000010;
    assign weights1[39][514] = 16'b0000000000000010;
    assign weights1[39][515] = 16'b0000000000000000;
    assign weights1[39][516] = 16'b1111111111111111;
    assign weights1[39][517] = 16'b1111111111111000;
    assign weights1[39][518] = 16'b1111111111110011;
    assign weights1[39][519] = 16'b1111111111110010;
    assign weights1[39][520] = 16'b1111111111010111;
    assign weights1[39][521] = 16'b1111111111100100;
    assign weights1[39][522] = 16'b1111111111011101;
    assign weights1[39][523] = 16'b1111111111011100;
    assign weights1[39][524] = 16'b1111111111011011;
    assign weights1[39][525] = 16'b1111111111100101;
    assign weights1[39][526] = 16'b1111111111100111;
    assign weights1[39][527] = 16'b1111111111001011;
    assign weights1[39][528] = 16'b1111111111100101;
    assign weights1[39][529] = 16'b1111111111100011;
    assign weights1[39][530] = 16'b1111111111101011;
    assign weights1[39][531] = 16'b1111111111110001;
    assign weights1[39][532] = 16'b1111111111100110;
    assign weights1[39][533] = 16'b1111111111011110;
    assign weights1[39][534] = 16'b1111111111010111;
    assign weights1[39][535] = 16'b1111111111001110;
    assign weights1[39][536] = 16'b1111111111001111;
    assign weights1[39][537] = 16'b1111111111101011;
    assign weights1[39][538] = 16'b1111111111101001;
    assign weights1[39][539] = 16'b1111111111111000;
    assign weights1[39][540] = 16'b1111111111101111;
    assign weights1[39][541] = 16'b1111111111110100;
    assign weights1[39][542] = 16'b0000000000000001;
    assign weights1[39][543] = 16'b1111111111111100;
    assign weights1[39][544] = 16'b1111111111101100;
    assign weights1[39][545] = 16'b1111111111110001;
    assign weights1[39][546] = 16'b1111111111110100;
    assign weights1[39][547] = 16'b1111111111110110;
    assign weights1[39][548] = 16'b1111111111110001;
    assign weights1[39][549] = 16'b1111111111101101;
    assign weights1[39][550] = 16'b1111111111011101;
    assign weights1[39][551] = 16'b1111111111011011;
    assign weights1[39][552] = 16'b1111111111100010;
    assign weights1[39][553] = 16'b1111111111000011;
    assign weights1[39][554] = 16'b1111111111001110;
    assign weights1[39][555] = 16'b1111111111011111;
    assign weights1[39][556] = 16'b1111111111111001;
    assign weights1[39][557] = 16'b1111111111101001;
    assign weights1[39][558] = 16'b1111111111100111;
    assign weights1[39][559] = 16'b1111111111110000;
    assign weights1[39][560] = 16'b1111111111100101;
    assign weights1[39][561] = 16'b1111111111101010;
    assign weights1[39][562] = 16'b1111111111100011;
    assign weights1[39][563] = 16'b1111111111011001;
    assign weights1[39][564] = 16'b1111111111011111;
    assign weights1[39][565] = 16'b1111111111111111;
    assign weights1[39][566] = 16'b0000000000000111;
    assign weights1[39][567] = 16'b1111111111111101;
    assign weights1[39][568] = 16'b1111111111111001;
    assign weights1[39][569] = 16'b1111111111111100;
    assign weights1[39][570] = 16'b1111111111111000;
    assign weights1[39][571] = 16'b1111111111111000;
    assign weights1[39][572] = 16'b1111111111110101;
    assign weights1[39][573] = 16'b1111111111111011;
    assign weights1[39][574] = 16'b1111111111101100;
    assign weights1[39][575] = 16'b1111111111101010;
    assign weights1[39][576] = 16'b1111111111110100;
    assign weights1[39][577] = 16'b1111111111010111;
    assign weights1[39][578] = 16'b1111111111101011;
    assign weights1[39][579] = 16'b1111111111010111;
    assign weights1[39][580] = 16'b1111111111010101;
    assign weights1[39][581] = 16'b1111111111011010;
    assign weights1[39][582] = 16'b1111111111011011;
    assign weights1[39][583] = 16'b1111111111100100;
    assign weights1[39][584] = 16'b1111111111101101;
    assign weights1[39][585] = 16'b1111111111110001;
    assign weights1[39][586] = 16'b1111111111110001;
    assign weights1[39][587] = 16'b1111111111101111;
    assign weights1[39][588] = 16'b1111111111110101;
    assign weights1[39][589] = 16'b1111111111110011;
    assign weights1[39][590] = 16'b1111111111101111;
    assign weights1[39][591] = 16'b1111111111100100;
    assign weights1[39][592] = 16'b1111111111100010;
    assign weights1[39][593] = 16'b0000000000011010;
    assign weights1[39][594] = 16'b0000000000000101;
    assign weights1[39][595] = 16'b1111111111110011;
    assign weights1[39][596] = 16'b1111111111111101;
    assign weights1[39][597] = 16'b1111111111100101;
    assign weights1[39][598] = 16'b0000000000000010;
    assign weights1[39][599] = 16'b1111111111111111;
    assign weights1[39][600] = 16'b1111111111101001;
    assign weights1[39][601] = 16'b1111111111101110;
    assign weights1[39][602] = 16'b1111111111101100;
    assign weights1[39][603] = 16'b1111111111101100;
    assign weights1[39][604] = 16'b1111111111110101;
    assign weights1[39][605] = 16'b1111111111110001;
    assign weights1[39][606] = 16'b1111111111100101;
    assign weights1[39][607] = 16'b1111111111110001;
    assign weights1[39][608] = 16'b1111111111011110;
    assign weights1[39][609] = 16'b1111111111110100;
    assign weights1[39][610] = 16'b1111111111110111;
    assign weights1[39][611] = 16'b1111111111100100;
    assign weights1[39][612] = 16'b1111111111101000;
    assign weights1[39][613] = 16'b1111111111101100;
    assign weights1[39][614] = 16'b1111111111111001;
    assign weights1[39][615] = 16'b1111111111110100;
    assign weights1[39][616] = 16'b1111111111111100;
    assign weights1[39][617] = 16'b1111111111110100;
    assign weights1[39][618] = 16'b1111111111111101;
    assign weights1[39][619] = 16'b1111111111110100;
    assign weights1[39][620] = 16'b1111111111111111;
    assign weights1[39][621] = 16'b0000000000000001;
    assign weights1[39][622] = 16'b1111111111100101;
    assign weights1[39][623] = 16'b1111111111111011;
    assign weights1[39][624] = 16'b0000000000101000;
    assign weights1[39][625] = 16'b0000000000011100;
    assign weights1[39][626] = 16'b1111111111111100;
    assign weights1[39][627] = 16'b1111111111101011;
    assign weights1[39][628] = 16'b0000000000000010;
    assign weights1[39][629] = 16'b1111111111111101;
    assign weights1[39][630] = 16'b1111111111111111;
    assign weights1[39][631] = 16'b0000000000001000;
    assign weights1[39][632] = 16'b1111111111100111;
    assign weights1[39][633] = 16'b0000000000000101;
    assign weights1[39][634] = 16'b1111111111101010;
    assign weights1[39][635] = 16'b1111111111101011;
    assign weights1[39][636] = 16'b1111111111101000;
    assign weights1[39][637] = 16'b1111111111111001;
    assign weights1[39][638] = 16'b1111111111111010;
    assign weights1[39][639] = 16'b1111111111101000;
    assign weights1[39][640] = 16'b1111111111101000;
    assign weights1[39][641] = 16'b1111111111100110;
    assign weights1[39][642] = 16'b1111111111110100;
    assign weights1[39][643] = 16'b1111111111110100;
    assign weights1[39][644] = 16'b1111111111111000;
    assign weights1[39][645] = 16'b1111111111110011;
    assign weights1[39][646] = 16'b1111111111110101;
    assign weights1[39][647] = 16'b1111111111111110;
    assign weights1[39][648] = 16'b1111111111110111;
    assign weights1[39][649] = 16'b0000000000001110;
    assign weights1[39][650] = 16'b1111111111110101;
    assign weights1[39][651] = 16'b1111111111110101;
    assign weights1[39][652] = 16'b1111111111101001;
    assign weights1[39][653] = 16'b1111111111100100;
    assign weights1[39][654] = 16'b1111111111011111;
    assign weights1[39][655] = 16'b1111111111011101;
    assign weights1[39][656] = 16'b1111111111111111;
    assign weights1[39][657] = 16'b1111111111101110;
    assign weights1[39][658] = 16'b1111111111110100;
    assign weights1[39][659] = 16'b1111111111101010;
    assign weights1[39][660] = 16'b1111111111110100;
    assign weights1[39][661] = 16'b1111111111111111;
    assign weights1[39][662] = 16'b1111111111110000;
    assign weights1[39][663] = 16'b1111111111101001;
    assign weights1[39][664] = 16'b1111111111110101;
    assign weights1[39][665] = 16'b1111111111101101;
    assign weights1[39][666] = 16'b1111111111101011;
    assign weights1[39][667] = 16'b1111111111100010;
    assign weights1[39][668] = 16'b1111111111100101;
    assign weights1[39][669] = 16'b1111111111101001;
    assign weights1[39][670] = 16'b1111111111110110;
    assign weights1[39][671] = 16'b1111111111111001;
    assign weights1[39][672] = 16'b1111111111111111;
    assign weights1[39][673] = 16'b1111111111111110;
    assign weights1[39][674] = 16'b1111111111110111;
    assign weights1[39][675] = 16'b0000000000000000;
    assign weights1[39][676] = 16'b1111111111111001;
    assign weights1[39][677] = 16'b0000000000010010;
    assign weights1[39][678] = 16'b0000000000001000;
    assign weights1[39][679] = 16'b0000000000001100;
    assign weights1[39][680] = 16'b0000000000100000;
    assign weights1[39][681] = 16'b1111111111101100;
    assign weights1[39][682] = 16'b0000000000001001;
    assign weights1[39][683] = 16'b1111111111110110;
    assign weights1[39][684] = 16'b1111111111101001;
    assign weights1[39][685] = 16'b1111111111101001;
    assign weights1[39][686] = 16'b1111111111011010;
    assign weights1[39][687] = 16'b1111111111010100;
    assign weights1[39][688] = 16'b0000000000001100;
    assign weights1[39][689] = 16'b0000000000000101;
    assign weights1[39][690] = 16'b1111111111110001;
    assign weights1[39][691] = 16'b1111111111101111;
    assign weights1[39][692] = 16'b1111111111100011;
    assign weights1[39][693] = 16'b1111111111110010;
    assign weights1[39][694] = 16'b1111111111110010;
    assign weights1[39][695] = 16'b1111111111110000;
    assign weights1[39][696] = 16'b1111111111100110;
    assign weights1[39][697] = 16'b1111111111101100;
    assign weights1[39][698] = 16'b1111111111110111;
    assign weights1[39][699] = 16'b1111111111111110;
    assign weights1[39][700] = 16'b0000000000000011;
    assign weights1[39][701] = 16'b1111111111110110;
    assign weights1[39][702] = 16'b1111111111111111;
    assign weights1[39][703] = 16'b1111111111111010;
    assign weights1[39][704] = 16'b0000000000000010;
    assign weights1[39][705] = 16'b0000000000001100;
    assign weights1[39][706] = 16'b0000000000010000;
    assign weights1[39][707] = 16'b0000000000001000;
    assign weights1[39][708] = 16'b0000000000001001;
    assign weights1[39][709] = 16'b1111111111011110;
    assign weights1[39][710] = 16'b0000000000001100;
    assign weights1[39][711] = 16'b0000000000101100;
    assign weights1[39][712] = 16'b0000000000001110;
    assign weights1[39][713] = 16'b0000000000000101;
    assign weights1[39][714] = 16'b1111111111111110;
    assign weights1[39][715] = 16'b0000000000010001;
    assign weights1[39][716] = 16'b1111111111110010;
    assign weights1[39][717] = 16'b1111111111001011;
    assign weights1[39][718] = 16'b1111111111101001;
    assign weights1[39][719] = 16'b1111111111011001;
    assign weights1[39][720] = 16'b1111111111100110;
    assign weights1[39][721] = 16'b1111111111110100;
    assign weights1[39][722] = 16'b1111111111110001;
    assign weights1[39][723] = 16'b1111111111101101;
    assign weights1[39][724] = 16'b1111111111101111;
    assign weights1[39][725] = 16'b1111111111110110;
    assign weights1[39][726] = 16'b1111111111111011;
    assign weights1[39][727] = 16'b1111111111111111;
    assign weights1[39][728] = 16'b1111111111111101;
    assign weights1[39][729] = 16'b1111111111111010;
    assign weights1[39][730] = 16'b0000000000000110;
    assign weights1[39][731] = 16'b0000000000000100;
    assign weights1[39][732] = 16'b1111111111111001;
    assign weights1[39][733] = 16'b0000000000010100;
    assign weights1[39][734] = 16'b0000000000010111;
    assign weights1[39][735] = 16'b0000000000000111;
    assign weights1[39][736] = 16'b0000000000001000;
    assign weights1[39][737] = 16'b0000000000001010;
    assign weights1[39][738] = 16'b1111111111110101;
    assign weights1[39][739] = 16'b1111111111111011;
    assign weights1[39][740] = 16'b0000000000001000;
    assign weights1[39][741] = 16'b0000000000000110;
    assign weights1[39][742] = 16'b0000000000000110;
    assign weights1[39][743] = 16'b0000000000000010;
    assign weights1[39][744] = 16'b1111111111101110;
    assign weights1[39][745] = 16'b1111111111011100;
    assign weights1[39][746] = 16'b1111111111101000;
    assign weights1[39][747] = 16'b1111111111011010;
    assign weights1[39][748] = 16'b1111111111011010;
    assign weights1[39][749] = 16'b1111111111101000;
    assign weights1[39][750] = 16'b1111111111110101;
    assign weights1[39][751] = 16'b1111111111110101;
    assign weights1[39][752] = 16'b1111111111110111;
    assign weights1[39][753] = 16'b1111111111111010;
    assign weights1[39][754] = 16'b1111111111111101;
    assign weights1[39][755] = 16'b1111111111111111;
    assign weights1[39][756] = 16'b0000000000000011;
    assign weights1[39][757] = 16'b0000000000000011;
    assign weights1[39][758] = 16'b0000000000000000;
    assign weights1[39][759] = 16'b0000000000001001;
    assign weights1[39][760] = 16'b0000000000000110;
    assign weights1[39][761] = 16'b1111111111111101;
    assign weights1[39][762] = 16'b1111111111111101;
    assign weights1[39][763] = 16'b0000000000000100;
    assign weights1[39][764] = 16'b1111111111111100;
    assign weights1[39][765] = 16'b0000000000010000;
    assign weights1[39][766] = 16'b0000000000000011;
    assign weights1[39][767] = 16'b1111111111101000;
    assign weights1[39][768] = 16'b1111111111101101;
    assign weights1[39][769] = 16'b1111111111111100;
    assign weights1[39][770] = 16'b1111111111110100;
    assign weights1[39][771] = 16'b1111111111101111;
    assign weights1[39][772] = 16'b1111111111100011;
    assign weights1[39][773] = 16'b1111111111100011;
    assign weights1[39][774] = 16'b1111111111001101;
    assign weights1[39][775] = 16'b1111111111011111;
    assign weights1[39][776] = 16'b1111111111100010;
    assign weights1[39][777] = 16'b1111111111100101;
    assign weights1[39][778] = 16'b1111111111101101;
    assign weights1[39][779] = 16'b1111111111110101;
    assign weights1[39][780] = 16'b1111111111110111;
    assign weights1[39][781] = 16'b1111111111111111;
    assign weights1[39][782] = 16'b0000000000000000;
    assign weights1[39][783] = 16'b0000000000000000;
    assign weights1[40][0] = 16'b0000000000000000;
    assign weights1[40][1] = 16'b1111111111111111;
    assign weights1[40][2] = 16'b0000000000000010;
    assign weights1[40][3] = 16'b1111111111111110;
    assign weights1[40][4] = 16'b0000000000000001;
    assign weights1[40][5] = 16'b0000000000000101;
    assign weights1[40][6] = 16'b0000000000000100;
    assign weights1[40][7] = 16'b0000000000001011;
    assign weights1[40][8] = 16'b0000000000010000;
    assign weights1[40][9] = 16'b0000000000011000;
    assign weights1[40][10] = 16'b0000000000001010;
    assign weights1[40][11] = 16'b0000000000010101;
    assign weights1[40][12] = 16'b0000000000000101;
    assign weights1[40][13] = 16'b0000000000000011;
    assign weights1[40][14] = 16'b1111111111111011;
    assign weights1[40][15] = 16'b1111111111110110;
    assign weights1[40][16] = 16'b0000000000000011;
    assign weights1[40][17] = 16'b0000000000000011;
    assign weights1[40][18] = 16'b1111111111111110;
    assign weights1[40][19] = 16'b0000000000000001;
    assign weights1[40][20] = 16'b1111111111111100;
    assign weights1[40][21] = 16'b0000000000000011;
    assign weights1[40][22] = 16'b0000000000000110;
    assign weights1[40][23] = 16'b0000000000000001;
    assign weights1[40][24] = 16'b0000000000000101;
    assign weights1[40][25] = 16'b0000000000000010;
    assign weights1[40][26] = 16'b0000000000000100;
    assign weights1[40][27] = 16'b0000000000000000;
    assign weights1[40][28] = 16'b0000000000000000;
    assign weights1[40][29] = 16'b0000000000000001;
    assign weights1[40][30] = 16'b1111111111111111;
    assign weights1[40][31] = 16'b0000000000000010;
    assign weights1[40][32] = 16'b0000000000001011;
    assign weights1[40][33] = 16'b0000000000010111;
    assign weights1[40][34] = 16'b0000000000010011;
    assign weights1[40][35] = 16'b0000000000010000;
    assign weights1[40][36] = 16'b0000000000010101;
    assign weights1[40][37] = 16'b0000000000011110;
    assign weights1[40][38] = 16'b0000000000010110;
    assign weights1[40][39] = 16'b0000000000010111;
    assign weights1[40][40] = 16'b0000000000010001;
    assign weights1[40][41] = 16'b0000000000010010;
    assign weights1[40][42] = 16'b0000000000010111;
    assign weights1[40][43] = 16'b0000000000011011;
    assign weights1[40][44] = 16'b0000000000001101;
    assign weights1[40][45] = 16'b0000000000010101;
    assign weights1[40][46] = 16'b0000000000000111;
    assign weights1[40][47] = 16'b0000000000000101;
    assign weights1[40][48] = 16'b0000000000001110;
    assign weights1[40][49] = 16'b0000000000010000;
    assign weights1[40][50] = 16'b0000000000001010;
    assign weights1[40][51] = 16'b0000000000001101;
    assign weights1[40][52] = 16'b0000000000000000;
    assign weights1[40][53] = 16'b0000000000000100;
    assign weights1[40][54] = 16'b0000000000000100;
    assign weights1[40][55] = 16'b0000000000000010;
    assign weights1[40][56] = 16'b0000000000000010;
    assign weights1[40][57] = 16'b0000000000000010;
    assign weights1[40][58] = 16'b0000000000000111;
    assign weights1[40][59] = 16'b0000000000001110;
    assign weights1[40][60] = 16'b0000000000011001;
    assign weights1[40][61] = 16'b0000000000010101;
    assign weights1[40][62] = 16'b0000000000011110;
    assign weights1[40][63] = 16'b0000000000001101;
    assign weights1[40][64] = 16'b0000000000011000;
    assign weights1[40][65] = 16'b0000000000011100;
    assign weights1[40][66] = 16'b0000000000000110;
    assign weights1[40][67] = 16'b0000000000001110;
    assign weights1[40][68] = 16'b0000000000011001;
    assign weights1[40][69] = 16'b0000000000001011;
    assign weights1[40][70] = 16'b0000000000100100;
    assign weights1[40][71] = 16'b0000000000010111;
    assign weights1[40][72] = 16'b0000000000001010;
    assign weights1[40][73] = 16'b0000000000001110;
    assign weights1[40][74] = 16'b0000000000100001;
    assign weights1[40][75] = 16'b0000000000000101;
    assign weights1[40][76] = 16'b0000000000010111;
    assign weights1[40][77] = 16'b0000000000011110;
    assign weights1[40][78] = 16'b0000000000001111;
    assign weights1[40][79] = 16'b0000000000001011;
    assign weights1[40][80] = 16'b0000000000001001;
    assign weights1[40][81] = 16'b0000000000001100;
    assign weights1[40][82] = 16'b0000000000001011;
    assign weights1[40][83] = 16'b0000000000001000;
    assign weights1[40][84] = 16'b0000000000000011;
    assign weights1[40][85] = 16'b0000000000000100;
    assign weights1[40][86] = 16'b0000000000001010;
    assign weights1[40][87] = 16'b0000000000010110;
    assign weights1[40][88] = 16'b0000000000011011;
    assign weights1[40][89] = 16'b0000000000011110;
    assign weights1[40][90] = 16'b0000000000011111;
    assign weights1[40][91] = 16'b0000000000101011;
    assign weights1[40][92] = 16'b0000000000100101;
    assign weights1[40][93] = 16'b0000000000001001;
    assign weights1[40][94] = 16'b0000000000011101;
    assign weights1[40][95] = 16'b0000000000001111;
    assign weights1[40][96] = 16'b0000000000011011;
    assign weights1[40][97] = 16'b0000000000011010;
    assign weights1[40][98] = 16'b0000000000010011;
    assign weights1[40][99] = 16'b1111111111100101;
    assign weights1[40][100] = 16'b1111111111111001;
    assign weights1[40][101] = 16'b0000000000010101;
    assign weights1[40][102] = 16'b1111111111111110;
    assign weights1[40][103] = 16'b1111111111111101;
    assign weights1[40][104] = 16'b0000000000100000;
    assign weights1[40][105] = 16'b0000000000001101;
    assign weights1[40][106] = 16'b0000000000001011;
    assign weights1[40][107] = 16'b0000000000010110;
    assign weights1[40][108] = 16'b0000000000001101;
    assign weights1[40][109] = 16'b0000000000010010;
    assign weights1[40][110] = 16'b0000000000010010;
    assign weights1[40][111] = 16'b0000000000000110;
    assign weights1[40][112] = 16'b0000000000000000;
    assign weights1[40][113] = 16'b0000000000001011;
    assign weights1[40][114] = 16'b0000000000001110;
    assign weights1[40][115] = 16'b0000000000100000;
    assign weights1[40][116] = 16'b0000000000011011;
    assign weights1[40][117] = 16'b0000000000010001;
    assign weights1[40][118] = 16'b0000000000100001;
    assign weights1[40][119] = 16'b0000000000100000;
    assign weights1[40][120] = 16'b0000000000010111;
    assign weights1[40][121] = 16'b0000000000010101;
    assign weights1[40][122] = 16'b0000000000100000;
    assign weights1[40][123] = 16'b0000000000001011;
    assign weights1[40][124] = 16'b1111111111110100;
    assign weights1[40][125] = 16'b0000000000000011;
    assign weights1[40][126] = 16'b0000000000001011;
    assign weights1[40][127] = 16'b1111111111111001;
    assign weights1[40][128] = 16'b0000000000001000;
    assign weights1[40][129] = 16'b1111111111101110;
    assign weights1[40][130] = 16'b1111111111111111;
    assign weights1[40][131] = 16'b0000000000010010;
    assign weights1[40][132] = 16'b0000000000000110;
    assign weights1[40][133] = 16'b0000000000001000;
    assign weights1[40][134] = 16'b1111111111111100;
    assign weights1[40][135] = 16'b0000000000100000;
    assign weights1[40][136] = 16'b0000000000001111;
    assign weights1[40][137] = 16'b0000000000010010;
    assign weights1[40][138] = 16'b0000000000011001;
    assign weights1[40][139] = 16'b0000000000001100;
    assign weights1[40][140] = 16'b0000000000000010;
    assign weights1[40][141] = 16'b0000000000000111;
    assign weights1[40][142] = 16'b0000000000011010;
    assign weights1[40][143] = 16'b0000000000101100;
    assign weights1[40][144] = 16'b0000000000011111;
    assign weights1[40][145] = 16'b0000000000001110;
    assign weights1[40][146] = 16'b0000000000010010;
    assign weights1[40][147] = 16'b0000000000010110;
    assign weights1[40][148] = 16'b1111111111111010;
    assign weights1[40][149] = 16'b0000000000000101;
    assign weights1[40][150] = 16'b1111111111110110;
    assign weights1[40][151] = 16'b1111111111111101;
    assign weights1[40][152] = 16'b0000000000011010;
    assign weights1[40][153] = 16'b0000000000001100;
    assign weights1[40][154] = 16'b0000000000010111;
    assign weights1[40][155] = 16'b0000000000111011;
    assign weights1[40][156] = 16'b0000000000011000;
    assign weights1[40][157] = 16'b0000000000010010;
    assign weights1[40][158] = 16'b1111111111110000;
    assign weights1[40][159] = 16'b0000000000101000;
    assign weights1[40][160] = 16'b0000000000010010;
    assign weights1[40][161] = 16'b0000000000000110;
    assign weights1[40][162] = 16'b1111111111101111;
    assign weights1[40][163] = 16'b0000000000001110;
    assign weights1[40][164] = 16'b0000000000011000;
    assign weights1[40][165] = 16'b0000000000011100;
    assign weights1[40][166] = 16'b0000000000011100;
    assign weights1[40][167] = 16'b0000000000011010;
    assign weights1[40][168] = 16'b0000000000000101;
    assign weights1[40][169] = 16'b0000000000001011;
    assign weights1[40][170] = 16'b0000000000011000;
    assign weights1[40][171] = 16'b0000000000011111;
    assign weights1[40][172] = 16'b0000000000001111;
    assign weights1[40][173] = 16'b0000000000011000;
    assign weights1[40][174] = 16'b0000000000011100;
    assign weights1[40][175] = 16'b0000000000010110;
    assign weights1[40][176] = 16'b0000000000000110;
    assign weights1[40][177] = 16'b0000000000011101;
    assign weights1[40][178] = 16'b0000000000000011;
    assign weights1[40][179] = 16'b0000000000000001;
    assign weights1[40][180] = 16'b1111111111110111;
    assign weights1[40][181] = 16'b0000000000000010;
    assign weights1[40][182] = 16'b0000000000001010;
    assign weights1[40][183] = 16'b0000000000001100;
    assign weights1[40][184] = 16'b1111111111111001;
    assign weights1[40][185] = 16'b0000000000001101;
    assign weights1[40][186] = 16'b0000000000000010;
    assign weights1[40][187] = 16'b0000000000011001;
    assign weights1[40][188] = 16'b0000000000000101;
    assign weights1[40][189] = 16'b1111111111111000;
    assign weights1[40][190] = 16'b0000000000101010;
    assign weights1[40][191] = 16'b0000000000101010;
    assign weights1[40][192] = 16'b0000000000011011;
    assign weights1[40][193] = 16'b0000000000011011;
    assign weights1[40][194] = 16'b0000000000100100;
    assign weights1[40][195] = 16'b0000000000011010;
    assign weights1[40][196] = 16'b0000000000000100;
    assign weights1[40][197] = 16'b0000000000010010;
    assign weights1[40][198] = 16'b0000000000010011;
    assign weights1[40][199] = 16'b0000000000001100;
    assign weights1[40][200] = 16'b0000000000010110;
    assign weights1[40][201] = 16'b0000000000011111;
    assign weights1[40][202] = 16'b0000000000100000;
    assign weights1[40][203] = 16'b1111111111110110;
    assign weights1[40][204] = 16'b0000000000000101;
    assign weights1[40][205] = 16'b0000000000000101;
    assign weights1[40][206] = 16'b0000000000001100;
    assign weights1[40][207] = 16'b0000000000001001;
    assign weights1[40][208] = 16'b0000000000000101;
    assign weights1[40][209] = 16'b0000000000001000;
    assign weights1[40][210] = 16'b1111111111110101;
    assign weights1[40][211] = 16'b1111111111101000;
    assign weights1[40][212] = 16'b1111111111110111;
    assign weights1[40][213] = 16'b1111111111111101;
    assign weights1[40][214] = 16'b0000000000010101;
    assign weights1[40][215] = 16'b0000000000011010;
    assign weights1[40][216] = 16'b1111111111111001;
    assign weights1[40][217] = 16'b0000000000010001;
    assign weights1[40][218] = 16'b0000000000011101;
    assign weights1[40][219] = 16'b0000000000011110;
    assign weights1[40][220] = 16'b0000000000010111;
    assign weights1[40][221] = 16'b0000000000110011;
    assign weights1[40][222] = 16'b0000000000101010;
    assign weights1[40][223] = 16'b0000000000100110;
    assign weights1[40][224] = 16'b0000000000000010;
    assign weights1[40][225] = 16'b0000000000001110;
    assign weights1[40][226] = 16'b0000000000001111;
    assign weights1[40][227] = 16'b0000000000001001;
    assign weights1[40][228] = 16'b0000000000000100;
    assign weights1[40][229] = 16'b0000000000010101;
    assign weights1[40][230] = 16'b0000000000011011;
    assign weights1[40][231] = 16'b0000000000011010;
    assign weights1[40][232] = 16'b1111111111110110;
    assign weights1[40][233] = 16'b0000000000010011;
    assign weights1[40][234] = 16'b0000000000001100;
    assign weights1[40][235] = 16'b0000000000000000;
    assign weights1[40][236] = 16'b0000000000001001;
    assign weights1[40][237] = 16'b0000000000100001;
    assign weights1[40][238] = 16'b1111111111111000;
    assign weights1[40][239] = 16'b1111111111110001;
    assign weights1[40][240] = 16'b1111111111100111;
    assign weights1[40][241] = 16'b0000000000001000;
    assign weights1[40][242] = 16'b0000000000100010;
    assign weights1[40][243] = 16'b0000000000000001;
    assign weights1[40][244] = 16'b1111111111111110;
    assign weights1[40][245] = 16'b0000000000011100;
    assign weights1[40][246] = 16'b0000000000000001;
    assign weights1[40][247] = 16'b0000000000000011;
    assign weights1[40][248] = 16'b0000000000011000;
    assign weights1[40][249] = 16'b0000000000001000;
    assign weights1[40][250] = 16'b0000000000100100;
    assign weights1[40][251] = 16'b0000000000100111;
    assign weights1[40][252] = 16'b0000000000000111;
    assign weights1[40][253] = 16'b0000000000001110;
    assign weights1[40][254] = 16'b0000000000001001;
    assign weights1[40][255] = 16'b0000000000001101;
    assign weights1[40][256] = 16'b1111111111111110;
    assign weights1[40][257] = 16'b0000000000001110;
    assign weights1[40][258] = 16'b0000000000001101;
    assign weights1[40][259] = 16'b1111111111111011;
    assign weights1[40][260] = 16'b1111111111110011;
    assign weights1[40][261] = 16'b0000000000010000;
    assign weights1[40][262] = 16'b0000000000001100;
    assign weights1[40][263] = 16'b1111111111110100;
    assign weights1[40][264] = 16'b1111111111110000;
    assign weights1[40][265] = 16'b0000000000101010;
    assign weights1[40][266] = 16'b0000000000001111;
    assign weights1[40][267] = 16'b0000000000000001;
    assign weights1[40][268] = 16'b1111111111100100;
    assign weights1[40][269] = 16'b0000000000010110;
    assign weights1[40][270] = 16'b0000000000001111;
    assign weights1[40][271] = 16'b0000000000000011;
    assign weights1[40][272] = 16'b0000000000000110;
    assign weights1[40][273] = 16'b1111111111111111;
    assign weights1[40][274] = 16'b1111111111110000;
    assign weights1[40][275] = 16'b0000000000001011;
    assign weights1[40][276] = 16'b1111111111111011;
    assign weights1[40][277] = 16'b1111111111111111;
    assign weights1[40][278] = 16'b0000000000100011;
    assign weights1[40][279] = 16'b0000000000011011;
    assign weights1[40][280] = 16'b0000000000001000;
    assign weights1[40][281] = 16'b0000000000010001;
    assign weights1[40][282] = 16'b0000000000010010;
    assign weights1[40][283] = 16'b0000000000011010;
    assign weights1[40][284] = 16'b0000000000011011;
    assign weights1[40][285] = 16'b1111111111110101;
    assign weights1[40][286] = 16'b1111111111111111;
    assign weights1[40][287] = 16'b0000000000001000;
    assign weights1[40][288] = 16'b0000000000001001;
    assign weights1[40][289] = 16'b0000000000011011;
    assign weights1[40][290] = 16'b0000000000000111;
    assign weights1[40][291] = 16'b1111111111110001;
    assign weights1[40][292] = 16'b1111111111111010;
    assign weights1[40][293] = 16'b0000000000010110;
    assign weights1[40][294] = 16'b0000000000101011;
    assign weights1[40][295] = 16'b1111111111101110;
    assign weights1[40][296] = 16'b1111111111101001;
    assign weights1[40][297] = 16'b0000000000001011;
    assign weights1[40][298] = 16'b0000000000000011;
    assign weights1[40][299] = 16'b1111111111101001;
    assign weights1[40][300] = 16'b0000000000010010;
    assign weights1[40][301] = 16'b1111111111111100;
    assign weights1[40][302] = 16'b1111111111111100;
    assign weights1[40][303] = 16'b0000000000011001;
    assign weights1[40][304] = 16'b0000000000000010;
    assign weights1[40][305] = 16'b0000000000000100;
    assign weights1[40][306] = 16'b0000000000010010;
    assign weights1[40][307] = 16'b0000000000100001;
    assign weights1[40][308] = 16'b0000000000000010;
    assign weights1[40][309] = 16'b0000000000010001;
    assign weights1[40][310] = 16'b0000000000010010;
    assign weights1[40][311] = 16'b0000000000000100;
    assign weights1[40][312] = 16'b1111111111111101;
    assign weights1[40][313] = 16'b1111111111110111;
    assign weights1[40][314] = 16'b0000000000001010;
    assign weights1[40][315] = 16'b1111111111111110;
    assign weights1[40][316] = 16'b0000000000010001;
    assign weights1[40][317] = 16'b0000000000010000;
    assign weights1[40][318] = 16'b0000000000010101;
    assign weights1[40][319] = 16'b0000000000000010;
    assign weights1[40][320] = 16'b1111111111111011;
    assign weights1[40][321] = 16'b0000000000000010;
    assign weights1[40][322] = 16'b0000000000010001;
    assign weights1[40][323] = 16'b1111111111101010;
    assign weights1[40][324] = 16'b1111111111110111;
    assign weights1[40][325] = 16'b1111111111111111;
    assign weights1[40][326] = 16'b1111111111111111;
    assign weights1[40][327] = 16'b1111111111111000;
    assign weights1[40][328] = 16'b1111111111110010;
    assign weights1[40][329] = 16'b1111111111110010;
    assign weights1[40][330] = 16'b0000000000001110;
    assign weights1[40][331] = 16'b0000000000010000;
    assign weights1[40][332] = 16'b0000000000011001;
    assign weights1[40][333] = 16'b0000000000000010;
    assign weights1[40][334] = 16'b0000000000100001;
    assign weights1[40][335] = 16'b0000000000100100;
    assign weights1[40][336] = 16'b0000000000001010;
    assign weights1[40][337] = 16'b0000000000010110;
    assign weights1[40][338] = 16'b0000000000011111;
    assign weights1[40][339] = 16'b0000000000001011;
    assign weights1[40][340] = 16'b0000000000000110;
    assign weights1[40][341] = 16'b0000000000001100;
    assign weights1[40][342] = 16'b0000000000001000;
    assign weights1[40][343] = 16'b1111111111111011;
    assign weights1[40][344] = 16'b0000000000001011;
    assign weights1[40][345] = 16'b0000000000000011;
    assign weights1[40][346] = 16'b1111111111111001;
    assign weights1[40][347] = 16'b0000000000000101;
    assign weights1[40][348] = 16'b0000000000000010;
    assign weights1[40][349] = 16'b0000000000000110;
    assign weights1[40][350] = 16'b0000000000000010;
    assign weights1[40][351] = 16'b1111111111111010;
    assign weights1[40][352] = 16'b0000000000001000;
    assign weights1[40][353] = 16'b0000000000001010;
    assign weights1[40][354] = 16'b1111111111101111;
    assign weights1[40][355] = 16'b0000000000010010;
    assign weights1[40][356] = 16'b1111111111111000;
    assign weights1[40][357] = 16'b0000000000010000;
    assign weights1[40][358] = 16'b1111111111111010;
    assign weights1[40][359] = 16'b1111111111111100;
    assign weights1[40][360] = 16'b0000000000000110;
    assign weights1[40][361] = 16'b0000000000001010;
    assign weights1[40][362] = 16'b0000000000100100;
    assign weights1[40][363] = 16'b0000000000101111;
    assign weights1[40][364] = 16'b0000000000010000;
    assign weights1[40][365] = 16'b0000000000011110;
    assign weights1[40][366] = 16'b0000000000011011;
    assign weights1[40][367] = 16'b0000000000100001;
    assign weights1[40][368] = 16'b0000000000011010;
    assign weights1[40][369] = 16'b1111111111111111;
    assign weights1[40][370] = 16'b1111111111111111;
    assign weights1[40][371] = 16'b1111111111111001;
    assign weights1[40][372] = 16'b0000000000011011;
    assign weights1[40][373] = 16'b1111111111111000;
    assign weights1[40][374] = 16'b0000000000011111;
    assign weights1[40][375] = 16'b0000000000010010;
    assign weights1[40][376] = 16'b1111111111101110;
    assign weights1[40][377] = 16'b1111111111111010;
    assign weights1[40][378] = 16'b1111111111110001;
    assign weights1[40][379] = 16'b0000000000100000;
    assign weights1[40][380] = 16'b1111111111101111;
    assign weights1[40][381] = 16'b1111111111101010;
    assign weights1[40][382] = 16'b1111111111111111;
    assign weights1[40][383] = 16'b0000000000010101;
    assign weights1[40][384] = 16'b0000000000011110;
    assign weights1[40][385] = 16'b1111111111111110;
    assign weights1[40][386] = 16'b0000000000000100;
    assign weights1[40][387] = 16'b1111111111100101;
    assign weights1[40][388] = 16'b1111111111111001;
    assign weights1[40][389] = 16'b0000000000001011;
    assign weights1[40][390] = 16'b0000000000100111;
    assign weights1[40][391] = 16'b0000000000101111;
    assign weights1[40][392] = 16'b0000000000010001;
    assign weights1[40][393] = 16'b0000000000010101;
    assign weights1[40][394] = 16'b0000000000011001;
    assign weights1[40][395] = 16'b0000000000011011;
    assign weights1[40][396] = 16'b0000000000001000;
    assign weights1[40][397] = 16'b0000000000001001;
    assign weights1[40][398] = 16'b0000000000000110;
    assign weights1[40][399] = 16'b0000000000000111;
    assign weights1[40][400] = 16'b0000000000001101;
    assign weights1[40][401] = 16'b1111111111111000;
    assign weights1[40][402] = 16'b0000000000010000;
    assign weights1[40][403] = 16'b0000000000001101;
    assign weights1[40][404] = 16'b1111111111111100;
    assign weights1[40][405] = 16'b1111111111110011;
    assign weights1[40][406] = 16'b1111111111111101;
    assign weights1[40][407] = 16'b0000000000010010;
    assign weights1[40][408] = 16'b0000000000000110;
    assign weights1[40][409] = 16'b0000000000000110;
    assign weights1[40][410] = 16'b0000000000000000;
    assign weights1[40][411] = 16'b1111111111101110;
    assign weights1[40][412] = 16'b0000000000000011;
    assign weights1[40][413] = 16'b0000000000000100;
    assign weights1[40][414] = 16'b1111111111101001;
    assign weights1[40][415] = 16'b1111111111100111;
    assign weights1[40][416] = 16'b1111111111110111;
    assign weights1[40][417] = 16'b0000000000011001;
    assign weights1[40][418] = 16'b0000000000011100;
    assign weights1[40][419] = 16'b0000000000111100;
    assign weights1[40][420] = 16'b0000000000010100;
    assign weights1[40][421] = 16'b0000000000011011;
    assign weights1[40][422] = 16'b0000000000010100;
    assign weights1[40][423] = 16'b0000000000000100;
    assign weights1[40][424] = 16'b0000000000011000;
    assign weights1[40][425] = 16'b0000000000001001;
    assign weights1[40][426] = 16'b0000000000000010;
    assign weights1[40][427] = 16'b0000000000100001;
    assign weights1[40][428] = 16'b0000000000001011;
    assign weights1[40][429] = 16'b0000000000011010;
    assign weights1[40][430] = 16'b0000000000001110;
    assign weights1[40][431] = 16'b1111111111111111;
    assign weights1[40][432] = 16'b1111111111111011;
    assign weights1[40][433] = 16'b0000000000011010;
    assign weights1[40][434] = 16'b1111111111111010;
    assign weights1[40][435] = 16'b1111111111110100;
    assign weights1[40][436] = 16'b0000000000011000;
    assign weights1[40][437] = 16'b0000000000000101;
    assign weights1[40][438] = 16'b1111111111011101;
    assign weights1[40][439] = 16'b1111111111111101;
    assign weights1[40][440] = 16'b1111111111011110;
    assign weights1[40][441] = 16'b0000000000000010;
    assign weights1[40][442] = 16'b0000000000001100;
    assign weights1[40][443] = 16'b1111111111111010;
    assign weights1[40][444] = 16'b0000000000001000;
    assign weights1[40][445] = 16'b0000000000100101;
    assign weights1[40][446] = 16'b0000000000101101;
    assign weights1[40][447] = 16'b0000000000101001;
    assign weights1[40][448] = 16'b0000000000010000;
    assign weights1[40][449] = 16'b0000000000010110;
    assign weights1[40][450] = 16'b0000000000001011;
    assign weights1[40][451] = 16'b0000000000000010;
    assign weights1[40][452] = 16'b1111111111111101;
    assign weights1[40][453] = 16'b1111111111111111;
    assign weights1[40][454] = 16'b0000000000000101;
    assign weights1[40][455] = 16'b0000000000001000;
    assign weights1[40][456] = 16'b0000000000010100;
    assign weights1[40][457] = 16'b0000000000000101;
    assign weights1[40][458] = 16'b0000000000000000;
    assign weights1[40][459] = 16'b0000000000001101;
    assign weights1[40][460] = 16'b1111111111111100;
    assign weights1[40][461] = 16'b0000000000000100;
    assign weights1[40][462] = 16'b1111111111111100;
    assign weights1[40][463] = 16'b1111111111101010;
    assign weights1[40][464] = 16'b1111111111101110;
    assign weights1[40][465] = 16'b0000000000011010;
    assign weights1[40][466] = 16'b0000000000001101;
    assign weights1[40][467] = 16'b1111111111111001;
    assign weights1[40][468] = 16'b0000000000000000;
    assign weights1[40][469] = 16'b1111111111110000;
    assign weights1[40][470] = 16'b0000000000000011;
    assign weights1[40][471] = 16'b0000000000010010;
    assign weights1[40][472] = 16'b0000000000001110;
    assign weights1[40][473] = 16'b0000000000011111;
    assign weights1[40][474] = 16'b0000000000110100;
    assign weights1[40][475] = 16'b0000000000100110;
    assign weights1[40][476] = 16'b0000000000001101;
    assign weights1[40][477] = 16'b0000000000001001;
    assign weights1[40][478] = 16'b1111111111111010;
    assign weights1[40][479] = 16'b1111111111111001;
    assign weights1[40][480] = 16'b1111111111110111;
    assign weights1[40][481] = 16'b0000000000010111;
    assign weights1[40][482] = 16'b0000000000000011;
    assign weights1[40][483] = 16'b0000000000000010;
    assign weights1[40][484] = 16'b1111111111111001;
    assign weights1[40][485] = 16'b0000000000000101;
    assign weights1[40][486] = 16'b1111111111111110;
    assign weights1[40][487] = 16'b0000000000000101;
    assign weights1[40][488] = 16'b0000000000001111;
    assign weights1[40][489] = 16'b1111111111111100;
    assign weights1[40][490] = 16'b0000000000000101;
    assign weights1[40][491] = 16'b1111111111010111;
    assign weights1[40][492] = 16'b0000000000010101;
    assign weights1[40][493] = 16'b0000000000010100;
    assign weights1[40][494] = 16'b0000000000001001;
    assign weights1[40][495] = 16'b0000000000001011;
    assign weights1[40][496] = 16'b0000000000001101;
    assign weights1[40][497] = 16'b0000000000000110;
    assign weights1[40][498] = 16'b0000000000001101;
    assign weights1[40][499] = 16'b0000000000010000;
    assign weights1[40][500] = 16'b0000000000010110;
    assign weights1[40][501] = 16'b0000000000010110;
    assign weights1[40][502] = 16'b0000000000100010;
    assign weights1[40][503] = 16'b0000000000100001;
    assign weights1[40][504] = 16'b1111111111111110;
    assign weights1[40][505] = 16'b0000000000000111;
    assign weights1[40][506] = 16'b0000000000000101;
    assign weights1[40][507] = 16'b0000000000000101;
    assign weights1[40][508] = 16'b1111111111111100;
    assign weights1[40][509] = 16'b0000000000001110;
    assign weights1[40][510] = 16'b1111111111111110;
    assign weights1[40][511] = 16'b0000000000010101;
    assign weights1[40][512] = 16'b0000000000000011;
    assign weights1[40][513] = 16'b0000000000000010;
    assign weights1[40][514] = 16'b0000000000001110;
    assign weights1[40][515] = 16'b0000000000001010;
    assign weights1[40][516] = 16'b1111111111111000;
    assign weights1[40][517] = 16'b0000000000100011;
    assign weights1[40][518] = 16'b0000000000011100;
    assign weights1[40][519] = 16'b0000000000000110;
    assign weights1[40][520] = 16'b1111111111111000;
    assign weights1[40][521] = 16'b0000000000001001;
    assign weights1[40][522] = 16'b0000000000000110;
    assign weights1[40][523] = 16'b0000000000001101;
    assign weights1[40][524] = 16'b0000000000011111;
    assign weights1[40][525] = 16'b0000000000001001;
    assign weights1[40][526] = 16'b0000000000100011;
    assign weights1[40][527] = 16'b0000000000011111;
    assign weights1[40][528] = 16'b0000000000011111;
    assign weights1[40][529] = 16'b0000000000011111;
    assign weights1[40][530] = 16'b0000000000101001;
    assign weights1[40][531] = 16'b0000000000010110;
    assign weights1[40][532] = 16'b0000000000000111;
    assign weights1[40][533] = 16'b0000000000001001;
    assign weights1[40][534] = 16'b0000000000000110;
    assign weights1[40][535] = 16'b0000000000000000;
    assign weights1[40][536] = 16'b0000000000000001;
    assign weights1[40][537] = 16'b0000000000001110;
    assign weights1[40][538] = 16'b0000000000010011;
    assign weights1[40][539] = 16'b0000000000011110;
    assign weights1[40][540] = 16'b0000000000001001;
    assign weights1[40][541] = 16'b1111111111110000;
    assign weights1[40][542] = 16'b0000000000001110;
    assign weights1[40][543] = 16'b0000000000000011;
    assign weights1[40][544] = 16'b1111111111111100;
    assign weights1[40][545] = 16'b1111111111111010;
    assign weights1[40][546] = 16'b1111111111111011;
    assign weights1[40][547] = 16'b0000000000010000;
    assign weights1[40][548] = 16'b0000000000000111;
    assign weights1[40][549] = 16'b1111111111110100;
    assign weights1[40][550] = 16'b1111111111111111;
    assign weights1[40][551] = 16'b0000000000100011;
    assign weights1[40][552] = 16'b0000000000010100;
    assign weights1[40][553] = 16'b0000000000011010;
    assign weights1[40][554] = 16'b0000000000101101;
    assign weights1[40][555] = 16'b0000000000110001;
    assign weights1[40][556] = 16'b0000000000010001;
    assign weights1[40][557] = 16'b0000000000101000;
    assign weights1[40][558] = 16'b0000000000100101;
    assign weights1[40][559] = 16'b0000000000100000;
    assign weights1[40][560] = 16'b0000000000011001;
    assign weights1[40][561] = 16'b0000000000001111;
    assign weights1[40][562] = 16'b0000000000010100;
    assign weights1[40][563] = 16'b0000000000011001;
    assign weights1[40][564] = 16'b0000000000011110;
    assign weights1[40][565] = 16'b0000000000010110;
    assign weights1[40][566] = 16'b0000000000011010;
    assign weights1[40][567] = 16'b0000000000100000;
    assign weights1[40][568] = 16'b0000000000001001;
    assign weights1[40][569] = 16'b1111111111111000;
    assign weights1[40][570] = 16'b0000000000111100;
    assign weights1[40][571] = 16'b1111111111101011;
    assign weights1[40][572] = 16'b0000000000000110;
    assign weights1[40][573] = 16'b1111111111111000;
    assign weights1[40][574] = 16'b1111111111101011;
    assign weights1[40][575] = 16'b0000000000011011;
    assign weights1[40][576] = 16'b0000000000011010;
    assign weights1[40][577] = 16'b1111111111101100;
    assign weights1[40][578] = 16'b0000000000001010;
    assign weights1[40][579] = 16'b0000000000001111;
    assign weights1[40][580] = 16'b0000000000000000;
    assign weights1[40][581] = 16'b0000000000101000;
    assign weights1[40][582] = 16'b0000000000101001;
    assign weights1[40][583] = 16'b0000000000101010;
    assign weights1[40][584] = 16'b0000000000011011;
    assign weights1[40][585] = 16'b0000000000100100;
    assign weights1[40][586] = 16'b0000000000011111;
    assign weights1[40][587] = 16'b0000000000100000;
    assign weights1[40][588] = 16'b0000000000010010;
    assign weights1[40][589] = 16'b0000000000010001;
    assign weights1[40][590] = 16'b0000000000001010;
    assign weights1[40][591] = 16'b0000000000000111;
    assign weights1[40][592] = 16'b0000000000000011;
    assign weights1[40][593] = 16'b0000000000011000;
    assign weights1[40][594] = 16'b1111111111111100;
    assign weights1[40][595] = 16'b0000000000011000;
    assign weights1[40][596] = 16'b0000000000001000;
    assign weights1[40][597] = 16'b0000000000011111;
    assign weights1[40][598] = 16'b1111111111110111;
    assign weights1[40][599] = 16'b0000000000010011;
    assign weights1[40][600] = 16'b0000000000010101;
    assign weights1[40][601] = 16'b1111111111101001;
    assign weights1[40][602] = 16'b1111111111011111;
    assign weights1[40][603] = 16'b0000000000101001;
    assign weights1[40][604] = 16'b0000000000010110;
    assign weights1[40][605] = 16'b1111111111101001;
    assign weights1[40][606] = 16'b0000000000001010;
    assign weights1[40][607] = 16'b0000000000101010;
    assign weights1[40][608] = 16'b0000000000011011;
    assign weights1[40][609] = 16'b0000000000001110;
    assign weights1[40][610] = 16'b0000000000011010;
    assign weights1[40][611] = 16'b0000000000101010;
    assign weights1[40][612] = 16'b0000000000011010;
    assign weights1[40][613] = 16'b0000000000101001;
    assign weights1[40][614] = 16'b0000000000011101;
    assign weights1[40][615] = 16'b0000000000011110;
    assign weights1[40][616] = 16'b0000000000011001;
    assign weights1[40][617] = 16'b0000000000011111;
    assign weights1[40][618] = 16'b0000000000010100;
    assign weights1[40][619] = 16'b0000000000001111;
    assign weights1[40][620] = 16'b1111111111111101;
    assign weights1[40][621] = 16'b0000000000010101;
    assign weights1[40][622] = 16'b0000000000001010;
    assign weights1[40][623] = 16'b0000000000010000;
    assign weights1[40][624] = 16'b0000000000000101;
    assign weights1[40][625] = 16'b0000000000010111;
    assign weights1[40][626] = 16'b1111111111110100;
    assign weights1[40][627] = 16'b0000000000001111;
    assign weights1[40][628] = 16'b0000000001000111;
    assign weights1[40][629] = 16'b0000000000011100;
    assign weights1[40][630] = 16'b1111111111111000;
    assign weights1[40][631] = 16'b0000000000110100;
    assign weights1[40][632] = 16'b0000000000010000;
    assign weights1[40][633] = 16'b1111111111011110;
    assign weights1[40][634] = 16'b0000000000010110;
    assign weights1[40][635] = 16'b0000000000011111;
    assign weights1[40][636] = 16'b0000000000011011;
    assign weights1[40][637] = 16'b0000000000011011;
    assign weights1[40][638] = 16'b0000000000001001;
    assign weights1[40][639] = 16'b0000000000100101;
    assign weights1[40][640] = 16'b0000000000101100;
    assign weights1[40][641] = 16'b0000000000101100;
    assign weights1[40][642] = 16'b0000000000011010;
    assign weights1[40][643] = 16'b0000000000010001;
    assign weights1[40][644] = 16'b0000000000010100;
    assign weights1[40][645] = 16'b0000000000010110;
    assign weights1[40][646] = 16'b0000000000011010;
    assign weights1[40][647] = 16'b0000000000011100;
    assign weights1[40][648] = 16'b0000000000010100;
    assign weights1[40][649] = 16'b0000000000010010;
    assign weights1[40][650] = 16'b0000000000011111;
    assign weights1[40][651] = 16'b1111111111111100;
    assign weights1[40][652] = 16'b0000000000011011;
    assign weights1[40][653] = 16'b0000000000000010;
    assign weights1[40][654] = 16'b1111111111111111;
    assign weights1[40][655] = 16'b0000000000010111;
    assign weights1[40][656] = 16'b0000000000110001;
    assign weights1[40][657] = 16'b0000000000101100;
    assign weights1[40][658] = 16'b0000000000001100;
    assign weights1[40][659] = 16'b0000000000010001;
    assign weights1[40][660] = 16'b0000000000100111;
    assign weights1[40][661] = 16'b1111111111111110;
    assign weights1[40][662] = 16'b0000000000001110;
    assign weights1[40][663] = 16'b0000000000101010;
    assign weights1[40][664] = 16'b0000000000001010;
    assign weights1[40][665] = 16'b1111111111111100;
    assign weights1[40][666] = 16'b0000000000000101;
    assign weights1[40][667] = 16'b0000000000100011;
    assign weights1[40][668] = 16'b0000000000011001;
    assign weights1[40][669] = 16'b0000000000011111;
    assign weights1[40][670] = 16'b0000000000001100;
    assign weights1[40][671] = 16'b0000000000010000;
    assign weights1[40][672] = 16'b0000000000001100;
    assign weights1[40][673] = 16'b0000000000001101;
    assign weights1[40][674] = 16'b0000000000001110;
    assign weights1[40][675] = 16'b0000000000010011;
    assign weights1[40][676] = 16'b0000000000010000;
    assign weights1[40][677] = 16'b0000000000001110;
    assign weights1[40][678] = 16'b1111111111110101;
    assign weights1[40][679] = 16'b1111111111111111;
    assign weights1[40][680] = 16'b0000000000000111;
    assign weights1[40][681] = 16'b1111111111110011;
    assign weights1[40][682] = 16'b0000000000000011;
    assign weights1[40][683] = 16'b0000000000011001;
    assign weights1[40][684] = 16'b0000000000000000;
    assign weights1[40][685] = 16'b1111111111111110;
    assign weights1[40][686] = 16'b0000000000000100;
    assign weights1[40][687] = 16'b0000000000001000;
    assign weights1[40][688] = 16'b0000000000001101;
    assign weights1[40][689] = 16'b1111111111101000;
    assign weights1[40][690] = 16'b0000000000010000;
    assign weights1[40][691] = 16'b0000000000010010;
    assign weights1[40][692] = 16'b0000000000000010;
    assign weights1[40][693] = 16'b1111111111111011;
    assign weights1[40][694] = 16'b0000000000000001;
    assign weights1[40][695] = 16'b0000000000001101;
    assign weights1[40][696] = 16'b0000000000010101;
    assign weights1[40][697] = 16'b0000000000100000;
    assign weights1[40][698] = 16'b0000000000010010;
    assign weights1[40][699] = 16'b0000000000000101;
    assign weights1[40][700] = 16'b0000000000000101;
    assign weights1[40][701] = 16'b0000000000001101;
    assign weights1[40][702] = 16'b0000000000000100;
    assign weights1[40][703] = 16'b0000000000010001;
    assign weights1[40][704] = 16'b0000000000001100;
    assign weights1[40][705] = 16'b0000000000001111;
    assign weights1[40][706] = 16'b0000000000001001;
    assign weights1[40][707] = 16'b0000000000001011;
    assign weights1[40][708] = 16'b0000000000001101;
    assign weights1[40][709] = 16'b0000000000010001;
    assign weights1[40][710] = 16'b0000000000011011;
    assign weights1[40][711] = 16'b0000000000001010;
    assign weights1[40][712] = 16'b1111111111101001;
    assign weights1[40][713] = 16'b1111111111011011;
    assign weights1[40][714] = 16'b1111111111110111;
    assign weights1[40][715] = 16'b0000000000000100;
    assign weights1[40][716] = 16'b1111111111111010;
    assign weights1[40][717] = 16'b0000000000000001;
    assign weights1[40][718] = 16'b0000000000001110;
    assign weights1[40][719] = 16'b0000000000001011;
    assign weights1[40][720] = 16'b0000000000001111;
    assign weights1[40][721] = 16'b1111111111110100;
    assign weights1[40][722] = 16'b0000000000000010;
    assign weights1[40][723] = 16'b0000000000010010;
    assign weights1[40][724] = 16'b0000000000010011;
    assign weights1[40][725] = 16'b0000000000010111;
    assign weights1[40][726] = 16'b0000000000010001;
    assign weights1[40][727] = 16'b0000000000000110;
    assign weights1[40][728] = 16'b0000000000000010;
    assign weights1[40][729] = 16'b0000000000000110;
    assign weights1[40][730] = 16'b0000000000000100;
    assign weights1[40][731] = 16'b1111111111111110;
    assign weights1[40][732] = 16'b0000000000000111;
    assign weights1[40][733] = 16'b0000000000001010;
    assign weights1[40][734] = 16'b0000000000000111;
    assign weights1[40][735] = 16'b0000000000011000;
    assign weights1[40][736] = 16'b0000000000011100;
    assign weights1[40][737] = 16'b0000000000011011;
    assign weights1[40][738] = 16'b0000000000001011;
    assign weights1[40][739] = 16'b0000000000011100;
    assign weights1[40][740] = 16'b0000000000001111;
    assign weights1[40][741] = 16'b0000000000001001;
    assign weights1[40][742] = 16'b0000000000100000;
    assign weights1[40][743] = 16'b0000000000011101;
    assign weights1[40][744] = 16'b0000000000010101;
    assign weights1[40][745] = 16'b0000000000011111;
    assign weights1[40][746] = 16'b0000000000011010;
    assign weights1[40][747] = 16'b0000000000010111;
    assign weights1[40][748] = 16'b0000000000000101;
    assign weights1[40][749] = 16'b0000000000010001;
    assign weights1[40][750] = 16'b0000000000010010;
    assign weights1[40][751] = 16'b0000000000010000;
    assign weights1[40][752] = 16'b0000000000010101;
    assign weights1[40][753] = 16'b0000000000001111;
    assign weights1[40][754] = 16'b0000000000000100;
    assign weights1[40][755] = 16'b1111111111111111;
    assign weights1[40][756] = 16'b0000000000000010;
    assign weights1[40][757] = 16'b1111111111111111;
    assign weights1[40][758] = 16'b0000000000000011;
    assign weights1[40][759] = 16'b1111111111111110;
    assign weights1[40][760] = 16'b0000000000000001;
    assign weights1[40][761] = 16'b0000000000001011;
    assign weights1[40][762] = 16'b0000000000001010;
    assign weights1[40][763] = 16'b0000000000010011;
    assign weights1[40][764] = 16'b0000000000010100;
    assign weights1[40][765] = 16'b0000000000010001;
    assign weights1[40][766] = 16'b0000000000001001;
    assign weights1[40][767] = 16'b0000000000100111;
    assign weights1[40][768] = 16'b0000000000011110;
    assign weights1[40][769] = 16'b0000000000011111;
    assign weights1[40][770] = 16'b0000000000100110;
    assign weights1[40][771] = 16'b0000000000100010;
    assign weights1[40][772] = 16'b0000000000000111;
    assign weights1[40][773] = 16'b0000000000010110;
    assign weights1[40][774] = 16'b0000000000010000;
    assign weights1[40][775] = 16'b0000000000001110;
    assign weights1[40][776] = 16'b0000000000001001;
    assign weights1[40][777] = 16'b0000000000010000;
    assign weights1[40][778] = 16'b0000000000001100;
    assign weights1[40][779] = 16'b0000000000010001;
    assign weights1[40][780] = 16'b0000000000001100;
    assign weights1[40][781] = 16'b0000000000000110;
    assign weights1[40][782] = 16'b0000000000000000;
    assign weights1[40][783] = 16'b1111111111111100;
    assign weights1[41][0] = 16'b0000000000000000;
    assign weights1[41][1] = 16'b0000000000000000;
    assign weights1[41][2] = 16'b1111111111111111;
    assign weights1[41][3] = 16'b1111111111111110;
    assign weights1[41][4] = 16'b1111111111111111;
    assign weights1[41][5] = 16'b1111111111111110;
    assign weights1[41][6] = 16'b1111111111111010;
    assign weights1[41][7] = 16'b1111111111110100;
    assign weights1[41][8] = 16'b1111111111100011;
    assign weights1[41][9] = 16'b1111111111100110;
    assign weights1[41][10] = 16'b1111111111100100;
    assign weights1[41][11] = 16'b1111111111010001;
    assign weights1[41][12] = 16'b1111111111001010;
    assign weights1[41][13] = 16'b1111111111001011;
    assign weights1[41][14] = 16'b1111111111010101;
    assign weights1[41][15] = 16'b1111111111001010;
    assign weights1[41][16] = 16'b1111111111001010;
    assign weights1[41][17] = 16'b1111111111010100;
    assign weights1[41][18] = 16'b1111111111011011;
    assign weights1[41][19] = 16'b1111111111100101;
    assign weights1[41][20] = 16'b1111111111100100;
    assign weights1[41][21] = 16'b1111111111110110;
    assign weights1[41][22] = 16'b1111111111110110;
    assign weights1[41][23] = 16'b1111111111111011;
    assign weights1[41][24] = 16'b0000000000000010;
    assign weights1[41][25] = 16'b0000000000000110;
    assign weights1[41][26] = 16'b0000000000000000;
    assign weights1[41][27] = 16'b0000000000000000;
    assign weights1[41][28] = 16'b0000000000000000;
    assign weights1[41][29] = 16'b0000000000000000;
    assign weights1[41][30] = 16'b1111111111111100;
    assign weights1[41][31] = 16'b1111111111111110;
    assign weights1[41][32] = 16'b1111111111111100;
    assign weights1[41][33] = 16'b1111111111111000;
    assign weights1[41][34] = 16'b1111111111111010;
    assign weights1[41][35] = 16'b1111111111110000;
    assign weights1[41][36] = 16'b1111111111011011;
    assign weights1[41][37] = 16'b1111111111010111;
    assign weights1[41][38] = 16'b1111111111011011;
    assign weights1[41][39] = 16'b1111111111100100;
    assign weights1[41][40] = 16'b1111111111100100;
    assign weights1[41][41] = 16'b1111111111100100;
    assign weights1[41][42] = 16'b1111111111100100;
    assign weights1[41][43] = 16'b1111111111010101;
    assign weights1[41][44] = 16'b1111111111100010;
    assign weights1[41][45] = 16'b1111111111100000;
    assign weights1[41][46] = 16'b1111111111100111;
    assign weights1[41][47] = 16'b1111111111111000;
    assign weights1[41][48] = 16'b1111111111110100;
    assign weights1[41][49] = 16'b0000000000000010;
    assign weights1[41][50] = 16'b0000000000000011;
    assign weights1[41][51] = 16'b0000000000000110;
    assign weights1[41][52] = 16'b0000000000000001;
    assign weights1[41][53] = 16'b0000000000000101;
    assign weights1[41][54] = 16'b0000000000000010;
    assign weights1[41][55] = 16'b0000000000000000;
    assign weights1[41][56] = 16'b0000000000000010;
    assign weights1[41][57] = 16'b0000000000000001;
    assign weights1[41][58] = 16'b1111111111111001;
    assign weights1[41][59] = 16'b1111111111111011;
    assign weights1[41][60] = 16'b0000000000000011;
    assign weights1[41][61] = 16'b0000000000000010;
    assign weights1[41][62] = 16'b1111111111111001;
    assign weights1[41][63] = 16'b1111111111111000;
    assign weights1[41][64] = 16'b1111111111101001;
    assign weights1[41][65] = 16'b1111111111101011;
    assign weights1[41][66] = 16'b1111111111101111;
    assign weights1[41][67] = 16'b0000000000000010;
    assign weights1[41][68] = 16'b1111111111100101;
    assign weights1[41][69] = 16'b1111111111110010;
    assign weights1[41][70] = 16'b1111111111110010;
    assign weights1[41][71] = 16'b1111111111111111;
    assign weights1[41][72] = 16'b0000000000000011;
    assign weights1[41][73] = 16'b0000000000000000;
    assign weights1[41][74] = 16'b0000000000000110;
    assign weights1[41][75] = 16'b1111111111110110;
    assign weights1[41][76] = 16'b0000000000000111;
    assign weights1[41][77] = 16'b0000000000000011;
    assign weights1[41][78] = 16'b1111111111111101;
    assign weights1[41][79] = 16'b1111111111111010;
    assign weights1[41][80] = 16'b0000000000000110;
    assign weights1[41][81] = 16'b1111111111111101;
    assign weights1[41][82] = 16'b1111111111111001;
    assign weights1[41][83] = 16'b1111111111111010;
    assign weights1[41][84] = 16'b0000000000000010;
    assign weights1[41][85] = 16'b1111111111111101;
    assign weights1[41][86] = 16'b1111111111111000;
    assign weights1[41][87] = 16'b0000000000000000;
    assign weights1[41][88] = 16'b0000000000001010;
    assign weights1[41][89] = 16'b0000000000001101;
    assign weights1[41][90] = 16'b0000000000001011;
    assign weights1[41][91] = 16'b0000000000000110;
    assign weights1[41][92] = 16'b0000000000000001;
    assign weights1[41][93] = 16'b0000000000000111;
    assign weights1[41][94] = 16'b0000000000000111;
    assign weights1[41][95] = 16'b1111111111111110;
    assign weights1[41][96] = 16'b1111111111110110;
    assign weights1[41][97] = 16'b0000000000010010;
    assign weights1[41][98] = 16'b0000000000001111;
    assign weights1[41][99] = 16'b1111111111110100;
    assign weights1[41][100] = 16'b0000000000000000;
    assign weights1[41][101] = 16'b0000000000000000;
    assign weights1[41][102] = 16'b1111111111110011;
    assign weights1[41][103] = 16'b1111111111101001;
    assign weights1[41][104] = 16'b1111111111111001;
    assign weights1[41][105] = 16'b0000000000000111;
    assign weights1[41][106] = 16'b1111111111100010;
    assign weights1[41][107] = 16'b1111111111101101;
    assign weights1[41][108] = 16'b0000000000000011;
    assign weights1[41][109] = 16'b1111111111111011;
    assign weights1[41][110] = 16'b1111111111111010;
    assign weights1[41][111] = 16'b1111111111111100;
    assign weights1[41][112] = 16'b0000000000000001;
    assign weights1[41][113] = 16'b0000000000000000;
    assign weights1[41][114] = 16'b1111111111111101;
    assign weights1[41][115] = 16'b0000000000000011;
    assign weights1[41][116] = 16'b0000000000010000;
    assign weights1[41][117] = 16'b0000000000010100;
    assign weights1[41][118] = 16'b0000000000010101;
    assign weights1[41][119] = 16'b0000000000001110;
    assign weights1[41][120] = 16'b0000000000001011;
    assign weights1[41][121] = 16'b0000000000010011;
    assign weights1[41][122] = 16'b0000000000000111;
    assign weights1[41][123] = 16'b0000000000011000;
    assign weights1[41][124] = 16'b0000000000010100;
    assign weights1[41][125] = 16'b0000000000001101;
    assign weights1[41][126] = 16'b0000000000011011;
    assign weights1[41][127] = 16'b0000000000011011;
    assign weights1[41][128] = 16'b0000000000001011;
    assign weights1[41][129] = 16'b0000000000000100;
    assign weights1[41][130] = 16'b0000000000001100;
    assign weights1[41][131] = 16'b0000000000001111;
    assign weights1[41][132] = 16'b1111111111100100;
    assign weights1[41][133] = 16'b1111111111110110;
    assign weights1[41][134] = 16'b1111111111101011;
    assign weights1[41][135] = 16'b1111111111101010;
    assign weights1[41][136] = 16'b0000000000001011;
    assign weights1[41][137] = 16'b1111111111111000;
    assign weights1[41][138] = 16'b1111111111111001;
    assign weights1[41][139] = 16'b0000000000000000;
    assign weights1[41][140] = 16'b0000000000000010;
    assign weights1[41][141] = 16'b0000000000001000;
    assign weights1[41][142] = 16'b0000000000001011;
    assign weights1[41][143] = 16'b1111111111111111;
    assign weights1[41][144] = 16'b0000000000000101;
    assign weights1[41][145] = 16'b0000000000101101;
    assign weights1[41][146] = 16'b0000000000011010;
    assign weights1[41][147] = 16'b0000000000010011;
    assign weights1[41][148] = 16'b1111111111110000;
    assign weights1[41][149] = 16'b0000000000010011;
    assign weights1[41][150] = 16'b1111111111101111;
    assign weights1[41][151] = 16'b0000000000010111;
    assign weights1[41][152] = 16'b0000000000100011;
    assign weights1[41][153] = 16'b0000000000010011;
    assign weights1[41][154] = 16'b0000000000000001;
    assign weights1[41][155] = 16'b1111111111111011;
    assign weights1[41][156] = 16'b0000000000001100;
    assign weights1[41][157] = 16'b0000000000000100;
    assign weights1[41][158] = 16'b1111111111111000;
    assign weights1[41][159] = 16'b1111111111110110;
    assign weights1[41][160] = 16'b0000000000011010;
    assign weights1[41][161] = 16'b0000000000001001;
    assign weights1[41][162] = 16'b0000000000010000;
    assign weights1[41][163] = 16'b0000000000101100;
    assign weights1[41][164] = 16'b0000000000010111;
    assign weights1[41][165] = 16'b0000000000000010;
    assign weights1[41][166] = 16'b1111111111111110;
    assign weights1[41][167] = 16'b1111111111111010;
    assign weights1[41][168] = 16'b0000000000000000;
    assign weights1[41][169] = 16'b1111111111111001;
    assign weights1[41][170] = 16'b0000000000000011;
    assign weights1[41][171] = 16'b0000000000000010;
    assign weights1[41][172] = 16'b1111111111111010;
    assign weights1[41][173] = 16'b0000000000011101;
    assign weights1[41][174] = 16'b0000000000010001;
    assign weights1[41][175] = 16'b0000000000011110;
    assign weights1[41][176] = 16'b0000000000001111;
    assign weights1[41][177] = 16'b1111111111111000;
    assign weights1[41][178] = 16'b0000000000100011;
    assign weights1[41][179] = 16'b0000000000100001;
    assign weights1[41][180] = 16'b0000000000010110;
    assign weights1[41][181] = 16'b0000000000001100;
    assign weights1[41][182] = 16'b0000000000001000;
    assign weights1[41][183] = 16'b0000000000001011;
    assign weights1[41][184] = 16'b0000000000000111;
    assign weights1[41][185] = 16'b0000000000100011;
    assign weights1[41][186] = 16'b0000000000011100;
    assign weights1[41][187] = 16'b0000000000011100;
    assign weights1[41][188] = 16'b0000000000011000;
    assign weights1[41][189] = 16'b0000000000011100;
    assign weights1[41][190] = 16'b0000000000010110;
    assign weights1[41][191] = 16'b0000000000010001;
    assign weights1[41][192] = 16'b0000000000000001;
    assign weights1[41][193] = 16'b0000000000000101;
    assign weights1[41][194] = 16'b0000000000000111;
    assign weights1[41][195] = 16'b0000000000000100;
    assign weights1[41][196] = 16'b1111111111111111;
    assign weights1[41][197] = 16'b1111111111110011;
    assign weights1[41][198] = 16'b1111111111110000;
    assign weights1[41][199] = 16'b1111111111111110;
    assign weights1[41][200] = 16'b0000000000010100;
    assign weights1[41][201] = 16'b0000000000011111;
    assign weights1[41][202] = 16'b0000000000010100;
    assign weights1[41][203] = 16'b1111111111111100;
    assign weights1[41][204] = 16'b1111111111111111;
    assign weights1[41][205] = 16'b1111111111111010;
    assign weights1[41][206] = 16'b0000000000000010;
    assign weights1[41][207] = 16'b0000000000010100;
    assign weights1[41][208] = 16'b1111111111101011;
    assign weights1[41][209] = 16'b0000000000001110;
    assign weights1[41][210] = 16'b0000000000001010;
    assign weights1[41][211] = 16'b0000000000100110;
    assign weights1[41][212] = 16'b0000000000101101;
    assign weights1[41][213] = 16'b0000000000101000;
    assign weights1[41][214] = 16'b0000000000010110;
    assign weights1[41][215] = 16'b0000000000110011;
    assign weights1[41][216] = 16'b0000000000001100;
    assign weights1[41][217] = 16'b0000000000010000;
    assign weights1[41][218] = 16'b1111111111111000;
    assign weights1[41][219] = 16'b0000000000010111;
    assign weights1[41][220] = 16'b0000000000100011;
    assign weights1[41][221] = 16'b0000000000101000;
    assign weights1[41][222] = 16'b0000000000010111;
    assign weights1[41][223] = 16'b0000000000001011;
    assign weights1[41][224] = 16'b1111111111110110;
    assign weights1[41][225] = 16'b1111111111110000;
    assign weights1[41][226] = 16'b1111111111110010;
    assign weights1[41][227] = 16'b0000000000000001;
    assign weights1[41][228] = 16'b0000000000000100;
    assign weights1[41][229] = 16'b0000000000101001;
    assign weights1[41][230] = 16'b0000000000110100;
    assign weights1[41][231] = 16'b1111111111111000;
    assign weights1[41][232] = 16'b1111111111110001;
    assign weights1[41][233] = 16'b0000000000000010;
    assign weights1[41][234] = 16'b1111111111110000;
    assign weights1[41][235] = 16'b1111111111111101;
    assign weights1[41][236] = 16'b0000000000010101;
    assign weights1[41][237] = 16'b0000000000100010;
    assign weights1[41][238] = 16'b0000000000011010;
    assign weights1[41][239] = 16'b0000000000101100;
    assign weights1[41][240] = 16'b0000000000011001;
    assign weights1[41][241] = 16'b0000000000000001;
    assign weights1[41][242] = 16'b0000000000100110;
    assign weights1[41][243] = 16'b0000000000001110;
    assign weights1[41][244] = 16'b0000000000001011;
    assign weights1[41][245] = 16'b0000000000000000;
    assign weights1[41][246] = 16'b0000000000010011;
    assign weights1[41][247] = 16'b0000000000110001;
    assign weights1[41][248] = 16'b0000000000111101;
    assign weights1[41][249] = 16'b0000000000110001;
    assign weights1[41][250] = 16'b0000000000011000;
    assign weights1[41][251] = 16'b0000000000000101;
    assign weights1[41][252] = 16'b1111111111110101;
    assign weights1[41][253] = 16'b1111111111101011;
    assign weights1[41][254] = 16'b1111111111110000;
    assign weights1[41][255] = 16'b0000000000000101;
    assign weights1[41][256] = 16'b0000000000011100;
    assign weights1[41][257] = 16'b0000000000111001;
    assign weights1[41][258] = 16'b0000000000111011;
    assign weights1[41][259] = 16'b0000000000011101;
    assign weights1[41][260] = 16'b0000000000100011;
    assign weights1[41][261] = 16'b0000000000010011;
    assign weights1[41][262] = 16'b0000000000000011;
    assign weights1[41][263] = 16'b1111111111110011;
    assign weights1[41][264] = 16'b1111111111011010;
    assign weights1[41][265] = 16'b1111111111110000;
    assign weights1[41][266] = 16'b1111111111100101;
    assign weights1[41][267] = 16'b1111111111101011;
    assign weights1[41][268] = 16'b1111111111101000;
    assign weights1[41][269] = 16'b1111111111111010;
    assign weights1[41][270] = 16'b1111111111111001;
    assign weights1[41][271] = 16'b1111111111110100;
    assign weights1[41][272] = 16'b0000000000010100;
    assign weights1[41][273] = 16'b0000000000100001;
    assign weights1[41][274] = 16'b0000000000100101;
    assign weights1[41][275] = 16'b0000000000111110;
    assign weights1[41][276] = 16'b0000000000110111;
    assign weights1[41][277] = 16'b0000000000001100;
    assign weights1[41][278] = 16'b0000000000001010;
    assign weights1[41][279] = 16'b1111111111111010;
    assign weights1[41][280] = 16'b1111111111110110;
    assign weights1[41][281] = 16'b1111111111110011;
    assign weights1[41][282] = 16'b1111111111100011;
    assign weights1[41][283] = 16'b0000000000000010;
    assign weights1[41][284] = 16'b0000000000011000;
    assign weights1[41][285] = 16'b0000000000101000;
    assign weights1[41][286] = 16'b0000000000101011;
    assign weights1[41][287] = 16'b0000000000100010;
    assign weights1[41][288] = 16'b0000000000100100;
    assign weights1[41][289] = 16'b0000000000101101;
    assign weights1[41][290] = 16'b0000000000010011;
    assign weights1[41][291] = 16'b1111111111100010;
    assign weights1[41][292] = 16'b1111111111110010;
    assign weights1[41][293] = 16'b1111111111001101;
    assign weights1[41][294] = 16'b1111111111011011;
    assign weights1[41][295] = 16'b1111111111001001;
    assign weights1[41][296] = 16'b1111111111011110;
    assign weights1[41][297] = 16'b1111111111011100;
    assign weights1[41][298] = 16'b1111111111101000;
    assign weights1[41][299] = 16'b1111111111110110;
    assign weights1[41][300] = 16'b0000000000001000;
    assign weights1[41][301] = 16'b1111111111111101;
    assign weights1[41][302] = 16'b0000000000100101;
    assign weights1[41][303] = 16'b0000000000001110;
    assign weights1[41][304] = 16'b0000000000010010;
    assign weights1[41][305] = 16'b1111111111101010;
    assign weights1[41][306] = 16'b1111111111100000;
    assign weights1[41][307] = 16'b1111111111100001;
    assign weights1[41][308] = 16'b1111111111110111;
    assign weights1[41][309] = 16'b1111111111100000;
    assign weights1[41][310] = 16'b1111111111010011;
    assign weights1[41][311] = 16'b1111111111110101;
    assign weights1[41][312] = 16'b0000000000000100;
    assign weights1[41][313] = 16'b0000000000010010;
    assign weights1[41][314] = 16'b0000000000100010;
    assign weights1[41][315] = 16'b0000000000110000;
    assign weights1[41][316] = 16'b0000000000010111;
    assign weights1[41][317] = 16'b0000000000100100;
    assign weights1[41][318] = 16'b0000000000101111;
    assign weights1[41][319] = 16'b0000000000010100;
    assign weights1[41][320] = 16'b0000000000011100;
    assign weights1[41][321] = 16'b0000000000000101;
    assign weights1[41][322] = 16'b0000000000101000;
    assign weights1[41][323] = 16'b1111111111110100;
    assign weights1[41][324] = 16'b0000000000001101;
    assign weights1[41][325] = 16'b0000000000011111;
    assign weights1[41][326] = 16'b0000000000010101;
    assign weights1[41][327] = 16'b0000000000010000;
    assign weights1[41][328] = 16'b1111111111110100;
    assign weights1[41][329] = 16'b0000000000001101;
    assign weights1[41][330] = 16'b1111111111011111;
    assign weights1[41][331] = 16'b1111111111011101;
    assign weights1[41][332] = 16'b1111111111010101;
    assign weights1[41][333] = 16'b1111111110111101;
    assign weights1[41][334] = 16'b1111111111000111;
    assign weights1[41][335] = 16'b1111111111011100;
    assign weights1[41][336] = 16'b1111111111101101;
    assign weights1[41][337] = 16'b1111111111011111;
    assign weights1[41][338] = 16'b1111111111001100;
    assign weights1[41][339] = 16'b1111111111010000;
    assign weights1[41][340] = 16'b1111111111111011;
    assign weights1[41][341] = 16'b0000000000011010;
    assign weights1[41][342] = 16'b0000000000010111;
    assign weights1[41][343] = 16'b0000000000110001;
    assign weights1[41][344] = 16'b0000000000110011;
    assign weights1[41][345] = 16'b0000000000110010;
    assign weights1[41][346] = 16'b0000000000001001;
    assign weights1[41][347] = 16'b0000000000100011;
    assign weights1[41][348] = 16'b0000000000011111;
    assign weights1[41][349] = 16'b0000000000010101;
    assign weights1[41][350] = 16'b0000000000110100;
    assign weights1[41][351] = 16'b0000000000010010;
    assign weights1[41][352] = 16'b0000000000001011;
    assign weights1[41][353] = 16'b0000000000011011;
    assign weights1[41][354] = 16'b0000000000010101;
    assign weights1[41][355] = 16'b0000000000100001;
    assign weights1[41][356] = 16'b0000000000101110;
    assign weights1[41][357] = 16'b0000000000001000;
    assign weights1[41][358] = 16'b1111111111110000;
    assign weights1[41][359] = 16'b1111111111010000;
    assign weights1[41][360] = 16'b1111111110101011;
    assign weights1[41][361] = 16'b1111111110110010;
    assign weights1[41][362] = 16'b1111111111000011;
    assign weights1[41][363] = 16'b1111111111010011;
    assign weights1[41][364] = 16'b1111111111101001;
    assign weights1[41][365] = 16'b1111111111011011;
    assign weights1[41][366] = 16'b1111111111000010;
    assign weights1[41][367] = 16'b1111111110111101;
    assign weights1[41][368] = 16'b1111111111011101;
    assign weights1[41][369] = 16'b1111111111100111;
    assign weights1[41][370] = 16'b0000000000010100;
    assign weights1[41][371] = 16'b0000000000110100;
    assign weights1[41][372] = 16'b0000000000110010;
    assign weights1[41][373] = 16'b0000000000011110;
    assign weights1[41][374] = 16'b0000000000100101;
    assign weights1[41][375] = 16'b0000000001001100;
    assign weights1[41][376] = 16'b0000000000101000;
    assign weights1[41][377] = 16'b0000000000100011;
    assign weights1[41][378] = 16'b0000000000001001;
    assign weights1[41][379] = 16'b0000000000010110;
    assign weights1[41][380] = 16'b0000000000011110;
    assign weights1[41][381] = 16'b0000000000010100;
    assign weights1[41][382] = 16'b0000000000011100;
    assign weights1[41][383] = 16'b0000000000001100;
    assign weights1[41][384] = 16'b0000000000011000;
    assign weights1[41][385] = 16'b0000000000000111;
    assign weights1[41][386] = 16'b1111111111010111;
    assign weights1[41][387] = 16'b1111111111010101;
    assign weights1[41][388] = 16'b1111111111000011;
    assign weights1[41][389] = 16'b1111111111001110;
    assign weights1[41][390] = 16'b1111111111010100;
    assign weights1[41][391] = 16'b1111111111011000;
    assign weights1[41][392] = 16'b1111111111100101;
    assign weights1[41][393] = 16'b1111111111010110;
    assign weights1[41][394] = 16'b1111111110111001;
    assign weights1[41][395] = 16'b1111111110100100;
    assign weights1[41][396] = 16'b1111111110100011;
    assign weights1[41][397] = 16'b1111111110111001;
    assign weights1[41][398] = 16'b1111111111110001;
    assign weights1[41][399] = 16'b1111111111111110;
    assign weights1[41][400] = 16'b0000000000101110;
    assign weights1[41][401] = 16'b0000000000100101;
    assign weights1[41][402] = 16'b0000000001001101;
    assign weights1[41][403] = 16'b0000000000010100;
    assign weights1[41][404] = 16'b0000000000100100;
    assign weights1[41][405] = 16'b0000000000101101;
    assign weights1[41][406] = 16'b0000000000011100;
    assign weights1[41][407] = 16'b0000000000100001;
    assign weights1[41][408] = 16'b0000000000011101;
    assign weights1[41][409] = 16'b0000000000010110;
    assign weights1[41][410] = 16'b0000000000010011;
    assign weights1[41][411] = 16'b1111111111011111;
    assign weights1[41][412] = 16'b1111111111100101;
    assign weights1[41][413] = 16'b1111111111100111;
    assign weights1[41][414] = 16'b1111111111001101;
    assign weights1[41][415] = 16'b1111111111100100;
    assign weights1[41][416] = 16'b1111111111101000;
    assign weights1[41][417] = 16'b1111111111101000;
    assign weights1[41][418] = 16'b1111111111011110;
    assign weights1[41][419] = 16'b1111111111011111;
    assign weights1[41][420] = 16'b1111111111101111;
    assign weights1[41][421] = 16'b1111111111100001;
    assign weights1[41][422] = 16'b1111111110111101;
    assign weights1[41][423] = 16'b1111111110110110;
    assign weights1[41][424] = 16'b1111111110001001;
    assign weights1[41][425] = 16'b1111111101100111;
    assign weights1[41][426] = 16'b1111111110000101;
    assign weights1[41][427] = 16'b1111111110101001;
    assign weights1[41][428] = 16'b1111111111010010;
    assign weights1[41][429] = 16'b1111111111111100;
    assign weights1[41][430] = 16'b0000000000101111;
    assign weights1[41][431] = 16'b0000000000100111;
    assign weights1[41][432] = 16'b0000000000010101;
    assign weights1[41][433] = 16'b0000000001000100;
    assign weights1[41][434] = 16'b0000000000100110;
    assign weights1[41][435] = 16'b0000000000100100;
    assign weights1[41][436] = 16'b0000000000010010;
    assign weights1[41][437] = 16'b0000000000001100;
    assign weights1[41][438] = 16'b1111111111101011;
    assign weights1[41][439] = 16'b1111111111110100;
    assign weights1[41][440] = 16'b1111111111101010;
    assign weights1[41][441] = 16'b1111111111011011;
    assign weights1[41][442] = 16'b1111111111110110;
    assign weights1[41][443] = 16'b1111111111111001;
    assign weights1[41][444] = 16'b1111111111111000;
    assign weights1[41][445] = 16'b1111111111101110;
    assign weights1[41][446] = 16'b1111111111011101;
    assign weights1[41][447] = 16'b1111111111100011;
    assign weights1[41][448] = 16'b1111111111110011;
    assign weights1[41][449] = 16'b1111111111101100;
    assign weights1[41][450] = 16'b1111111111010110;
    assign weights1[41][451] = 16'b1111111111000010;
    assign weights1[41][452] = 16'b1111111110001101;
    assign weights1[41][453] = 16'b1111111110001000;
    assign weights1[41][454] = 16'b1111111101010011;
    assign weights1[41][455] = 16'b1111111101010101;
    assign weights1[41][456] = 16'b1111111101111001;
    assign weights1[41][457] = 16'b1111111110010111;
    assign weights1[41][458] = 16'b1111111110111100;
    assign weights1[41][459] = 16'b1111111111110001;
    assign weights1[41][460] = 16'b0000000000010111;
    assign weights1[41][461] = 16'b0000000000010011;
    assign weights1[41][462] = 16'b0000000000001110;
    assign weights1[41][463] = 16'b0000000000010010;
    assign weights1[41][464] = 16'b0000000000001000;
    assign weights1[41][465] = 16'b1111111111101010;
    assign weights1[41][466] = 16'b1111111111101010;
    assign weights1[41][467] = 16'b1111111111101101;
    assign weights1[41][468] = 16'b1111111111010101;
    assign weights1[41][469] = 16'b1111111111110111;
    assign weights1[41][470] = 16'b1111111111111001;
    assign weights1[41][471] = 16'b0000000000010000;
    assign weights1[41][472] = 16'b0000000000010000;
    assign weights1[41][473] = 16'b1111111111111011;
    assign weights1[41][474] = 16'b1111111111101010;
    assign weights1[41][475] = 16'b1111111111100110;
    assign weights1[41][476] = 16'b1111111111111100;
    assign weights1[41][477] = 16'b1111111111111011;
    assign weights1[41][478] = 16'b1111111111110111;
    assign weights1[41][479] = 16'b1111111111110010;
    assign weights1[41][480] = 16'b1111111111100100;
    assign weights1[41][481] = 16'b1111111111010111;
    assign weights1[41][482] = 16'b1111111110100111;
    assign weights1[41][483] = 16'b1111111110001111;
    assign weights1[41][484] = 16'b1111111101111010;
    assign weights1[41][485] = 16'b1111111101101010;
    assign weights1[41][486] = 16'b1111111110000010;
    assign weights1[41][487] = 16'b1111111110011001;
    assign weights1[41][488] = 16'b1111111110100010;
    assign weights1[41][489] = 16'b1111111110100011;
    assign weights1[41][490] = 16'b1111111110111010;
    assign weights1[41][491] = 16'b1111111111001111;
    assign weights1[41][492] = 16'b1111111111110000;
    assign weights1[41][493] = 16'b1111111111101010;
    assign weights1[41][494] = 16'b1111111111110010;
    assign weights1[41][495] = 16'b1111111111011111;
    assign weights1[41][496] = 16'b0000000000000101;
    assign weights1[41][497] = 16'b0000000000011100;
    assign weights1[41][498] = 16'b1111111111111101;
    assign weights1[41][499] = 16'b0000000000100111;
    assign weights1[41][500] = 16'b0000000000000100;
    assign weights1[41][501] = 16'b1111111111111011;
    assign weights1[41][502] = 16'b0000000000000000;
    assign weights1[41][503] = 16'b1111111111100110;
    assign weights1[41][504] = 16'b1111111111111100;
    assign weights1[41][505] = 16'b1111111111111100;
    assign weights1[41][506] = 16'b0000000000000010;
    assign weights1[41][507] = 16'b0000000000001101;
    assign weights1[41][508] = 16'b0000000000001001;
    assign weights1[41][509] = 16'b0000000000010111;
    assign weights1[41][510] = 16'b0000000000011001;
    assign weights1[41][511] = 16'b1111111111101110;
    assign weights1[41][512] = 16'b1111111111001100;
    assign weights1[41][513] = 16'b1111111110110100;
    assign weights1[41][514] = 16'b1111111110111110;
    assign weights1[41][515] = 16'b1111111110111101;
    assign weights1[41][516] = 16'b1111111110100101;
    assign weights1[41][517] = 16'b1111111110111001;
    assign weights1[41][518] = 16'b1111111110101110;
    assign weights1[41][519] = 16'b1111111111011000;
    assign weights1[41][520] = 16'b1111111111100000;
    assign weights1[41][521] = 16'b1111111111100001;
    assign weights1[41][522] = 16'b1111111111100101;
    assign weights1[41][523] = 16'b1111111111111111;
    assign weights1[41][524] = 16'b0000000000001001;
    assign weights1[41][525] = 16'b0000000000000010;
    assign weights1[41][526] = 16'b0000000000001001;
    assign weights1[41][527] = 16'b0000000000010110;
    assign weights1[41][528] = 16'b0000000000000110;
    assign weights1[41][529] = 16'b0000000000000111;
    assign weights1[41][530] = 16'b1111111111110010;
    assign weights1[41][531] = 16'b1111111111101011;
    assign weights1[41][532] = 16'b0000000000000011;
    assign weights1[41][533] = 16'b0000000000001110;
    assign weights1[41][534] = 16'b0000000000001001;
    assign weights1[41][535] = 16'b0000000000001111;
    assign weights1[41][536] = 16'b0000000000100000;
    assign weights1[41][537] = 16'b0000000001000000;
    assign weights1[41][538] = 16'b0000000000111010;
    assign weights1[41][539] = 16'b0000000000101101;
    assign weights1[41][540] = 16'b0000000000100011;
    assign weights1[41][541] = 16'b0000000000001101;
    assign weights1[41][542] = 16'b0000000000000101;
    assign weights1[41][543] = 16'b1111111111100101;
    assign weights1[41][544] = 16'b1111111111110111;
    assign weights1[41][545] = 16'b1111111111110110;
    assign weights1[41][546] = 16'b1111111111101100;
    assign weights1[41][547] = 16'b1111111111100010;
    assign weights1[41][548] = 16'b1111111111101011;
    assign weights1[41][549] = 16'b0000000000001001;
    assign weights1[41][550] = 16'b1111111111110010;
    assign weights1[41][551] = 16'b1111111111101011;
    assign weights1[41][552] = 16'b1111111111101100;
    assign weights1[41][553] = 16'b1111111111101111;
    assign weights1[41][554] = 16'b1111111111110100;
    assign weights1[41][555] = 16'b1111111111110100;
    assign weights1[41][556] = 16'b0000000000001100;
    assign weights1[41][557] = 16'b0000000000010001;
    assign weights1[41][558] = 16'b1111111111111011;
    assign weights1[41][559] = 16'b1111111111110011;
    assign weights1[41][560] = 16'b0000000000000101;
    assign weights1[41][561] = 16'b0000000000001000;
    assign weights1[41][562] = 16'b0000000000001101;
    assign weights1[41][563] = 16'b0000000000010001;
    assign weights1[41][564] = 16'b0000000000001011;
    assign weights1[41][565] = 16'b0000000000001101;
    assign weights1[41][566] = 16'b0000000000010011;
    assign weights1[41][567] = 16'b0000000000010100;
    assign weights1[41][568] = 16'b0000000000011010;
    assign weights1[41][569] = 16'b0000000000000101;
    assign weights1[41][570] = 16'b0000000000001001;
    assign weights1[41][571] = 16'b0000000000010101;
    assign weights1[41][572] = 16'b1111111111111001;
    assign weights1[41][573] = 16'b1111111111111111;
    assign weights1[41][574] = 16'b0000000000001010;
    assign weights1[41][575] = 16'b0000000000000001;
    assign weights1[41][576] = 16'b1111111111110010;
    assign weights1[41][577] = 16'b0000000000000111;
    assign weights1[41][578] = 16'b1111111111101011;
    assign weights1[41][579] = 16'b1111111111110011;
    assign weights1[41][580] = 16'b1111111111110000;
    assign weights1[41][581] = 16'b0000000000001101;
    assign weights1[41][582] = 16'b1111111111110100;
    assign weights1[41][583] = 16'b1111111111111111;
    assign weights1[41][584] = 16'b0000000000000101;
    assign weights1[41][585] = 16'b0000000000001110;
    assign weights1[41][586] = 16'b1111111111111101;
    assign weights1[41][587] = 16'b1111111111101101;
    assign weights1[41][588] = 16'b1111111111111110;
    assign weights1[41][589] = 16'b0000000000000111;
    assign weights1[41][590] = 16'b1111111111111110;
    assign weights1[41][591] = 16'b1111111111111010;
    assign weights1[41][592] = 16'b1111111111110110;
    assign weights1[41][593] = 16'b0000000000100011;
    assign weights1[41][594] = 16'b0000000000010101;
    assign weights1[41][595] = 16'b1111111111110011;
    assign weights1[41][596] = 16'b0000000000000000;
    assign weights1[41][597] = 16'b0000000000011000;
    assign weights1[41][598] = 16'b0000000000001101;
    assign weights1[41][599] = 16'b1111111111110010;
    assign weights1[41][600] = 16'b0000000000010001;
    assign weights1[41][601] = 16'b1111111111101010;
    assign weights1[41][602] = 16'b1111111111110001;
    assign weights1[41][603] = 16'b1111111111101001;
    assign weights1[41][604] = 16'b1111111111101011;
    assign weights1[41][605] = 16'b1111111111111110;
    assign weights1[41][606] = 16'b1111111111110101;
    assign weights1[41][607] = 16'b1111111111111011;
    assign weights1[41][608] = 16'b0000000000010000;
    assign weights1[41][609] = 16'b0000000000010000;
    assign weights1[41][610] = 16'b0000000000001010;
    assign weights1[41][611] = 16'b1111111111011011;
    assign weights1[41][612] = 16'b0000000000001011;
    assign weights1[41][613] = 16'b0000000000010000;
    assign weights1[41][614] = 16'b1111111111111011;
    assign weights1[41][615] = 16'b1111111111111001;
    assign weights1[41][616] = 16'b1111111111110100;
    assign weights1[41][617] = 16'b1111111111111000;
    assign weights1[41][618] = 16'b1111111111101011;
    assign weights1[41][619] = 16'b1111111111110111;
    assign weights1[41][620] = 16'b0000000000001001;
    assign weights1[41][621] = 16'b0000000000010000;
    assign weights1[41][622] = 16'b1111111111101100;
    assign weights1[41][623] = 16'b0000000000001110;
    assign weights1[41][624] = 16'b1111111111110001;
    assign weights1[41][625] = 16'b0000000000001111;
    assign weights1[41][626] = 16'b1111111111101100;
    assign weights1[41][627] = 16'b1111111111101011;
    assign weights1[41][628] = 16'b1111111111111101;
    assign weights1[41][629] = 16'b0000000000000010;
    assign weights1[41][630] = 16'b0000000000001010;
    assign weights1[41][631] = 16'b0000000000000110;
    assign weights1[41][632] = 16'b0000000000001101;
    assign weights1[41][633] = 16'b0000000000000101;
    assign weights1[41][634] = 16'b1111111111101001;
    assign weights1[41][635] = 16'b1111111111110001;
    assign weights1[41][636] = 16'b1111111111110100;
    assign weights1[41][637] = 16'b0000000000011010;
    assign weights1[41][638] = 16'b1111111111101110;
    assign weights1[41][639] = 16'b1111111111111111;
    assign weights1[41][640] = 16'b1111111111111000;
    assign weights1[41][641] = 16'b1111111111111001;
    assign weights1[41][642] = 16'b1111111111110001;
    assign weights1[41][643] = 16'b1111111111111011;
    assign weights1[41][644] = 16'b1111111111111000;
    assign weights1[41][645] = 16'b1111111111110011;
    assign weights1[41][646] = 16'b1111111111101101;
    assign weights1[41][647] = 16'b1111111111110100;
    assign weights1[41][648] = 16'b1111111111101110;
    assign weights1[41][649] = 16'b1111111111101111;
    assign weights1[41][650] = 16'b0000000000001000;
    assign weights1[41][651] = 16'b1111111111110000;
    assign weights1[41][652] = 16'b0000000000010000;
    assign weights1[41][653] = 16'b0000000000000100;
    assign weights1[41][654] = 16'b1111111111111101;
    assign weights1[41][655] = 16'b0000000000100111;
    assign weights1[41][656] = 16'b0000000000001110;
    assign weights1[41][657] = 16'b0000000000000000;
    assign weights1[41][658] = 16'b0000000000010010;
    assign weights1[41][659] = 16'b1111111111110001;
    assign weights1[41][660] = 16'b1111111111111000;
    assign weights1[41][661] = 16'b1111111111110111;
    assign weights1[41][662] = 16'b1111111111110011;
    assign weights1[41][663] = 16'b1111111111111101;
    assign weights1[41][664] = 16'b1111111111101110;
    assign weights1[41][665] = 16'b0000000000010011;
    assign weights1[41][666] = 16'b1111111111101100;
    assign weights1[41][667] = 16'b1111111111111100;
    assign weights1[41][668] = 16'b1111111111101110;
    assign weights1[41][669] = 16'b1111111111111001;
    assign weights1[41][670] = 16'b1111111111111101;
    assign weights1[41][671] = 16'b1111111111111110;
    assign weights1[41][672] = 16'b1111111111110111;
    assign weights1[41][673] = 16'b1111111111111011;
    assign weights1[41][674] = 16'b1111111111110001;
    assign weights1[41][675] = 16'b1111111111101110;
    assign weights1[41][676] = 16'b1111111111111001;
    assign weights1[41][677] = 16'b1111111111110000;
    assign weights1[41][678] = 16'b1111111111110011;
    assign weights1[41][679] = 16'b0000000000000111;
    assign weights1[41][680] = 16'b0000000000000110;
    assign weights1[41][681] = 16'b1111111111100011;
    assign weights1[41][682] = 16'b0000000000000110;
    assign weights1[41][683] = 16'b0000000000010100;
    assign weights1[41][684] = 16'b1111111111101010;
    assign weights1[41][685] = 16'b0000000000001101;
    assign weights1[41][686] = 16'b0000000000000010;
    assign weights1[41][687] = 16'b1111111111110100;
    assign weights1[41][688] = 16'b1111111111101010;
    assign weights1[41][689] = 16'b1111111111101010;
    assign weights1[41][690] = 16'b1111111111100101;
    assign weights1[41][691] = 16'b1111111111111100;
    assign weights1[41][692] = 16'b0000000000001010;
    assign weights1[41][693] = 16'b0000000000000110;
    assign weights1[41][694] = 16'b1111111111101110;
    assign weights1[41][695] = 16'b1111111111110010;
    assign weights1[41][696] = 16'b1111111111110011;
    assign weights1[41][697] = 16'b1111111111110000;
    assign weights1[41][698] = 16'b0000000000000001;
    assign weights1[41][699] = 16'b1111111111111110;
    assign weights1[41][700] = 16'b1111111111111011;
    assign weights1[41][701] = 16'b1111111111110111;
    assign weights1[41][702] = 16'b1111111111110110;
    assign weights1[41][703] = 16'b1111111111110100;
    assign weights1[41][704] = 16'b1111111111100111;
    assign weights1[41][705] = 16'b1111111111100111;
    assign weights1[41][706] = 16'b1111111111011010;
    assign weights1[41][707] = 16'b1111111111110101;
    assign weights1[41][708] = 16'b1111111111110001;
    assign weights1[41][709] = 16'b1111111111101011;
    assign weights1[41][710] = 16'b1111111111110111;
    assign weights1[41][711] = 16'b0000000000000010;
    assign weights1[41][712] = 16'b1111111111100110;
    assign weights1[41][713] = 16'b0000000000010000;
    assign weights1[41][714] = 16'b1111111111100110;
    assign weights1[41][715] = 16'b1111111111110000;
    assign weights1[41][716] = 16'b0000000000000001;
    assign weights1[41][717] = 16'b0000000000000100;
    assign weights1[41][718] = 16'b1111111111110110;
    assign weights1[41][719] = 16'b0000000000010000;
    assign weights1[41][720] = 16'b0000000000010000;
    assign weights1[41][721] = 16'b0000000000000000;
    assign weights1[41][722] = 16'b0000000000000110;
    assign weights1[41][723] = 16'b1111111111111101;
    assign weights1[41][724] = 16'b1111111111111001;
    assign weights1[41][725] = 16'b1111111111111000;
    assign weights1[41][726] = 16'b1111111111111011;
    assign weights1[41][727] = 16'b1111111111111110;
    assign weights1[41][728] = 16'b1111111111111110;
    assign weights1[41][729] = 16'b1111111111110111;
    assign weights1[41][730] = 16'b1111111111110101;
    assign weights1[41][731] = 16'b1111111111111010;
    assign weights1[41][732] = 16'b1111111111110111;
    assign weights1[41][733] = 16'b1111111111111010;
    assign weights1[41][734] = 16'b1111111111101001;
    assign weights1[41][735] = 16'b1111111111101001;
    assign weights1[41][736] = 16'b1111111111101001;
    assign weights1[41][737] = 16'b1111111111100010;
    assign weights1[41][738] = 16'b1111111111110110;
    assign weights1[41][739] = 16'b1111111111101110;
    assign weights1[41][740] = 16'b1111111111110010;
    assign weights1[41][741] = 16'b1111111111111101;
    assign weights1[41][742] = 16'b0000000000001001;
    assign weights1[41][743] = 16'b1111111111101110;
    assign weights1[41][744] = 16'b0000000000010110;
    assign weights1[41][745] = 16'b0000000000001001;
    assign weights1[41][746] = 16'b1111111111101110;
    assign weights1[41][747] = 16'b1111111111110111;
    assign weights1[41][748] = 16'b1111111111111010;
    assign weights1[41][749] = 16'b1111111111111010;
    assign weights1[41][750] = 16'b0000000000000111;
    assign weights1[41][751] = 16'b0000000000000010;
    assign weights1[41][752] = 16'b1111111111111011;
    assign weights1[41][753] = 16'b1111111111111011;
    assign weights1[41][754] = 16'b1111111111111101;
    assign weights1[41][755] = 16'b0000000000000000;
    assign weights1[41][756] = 16'b0000000000000000;
    assign weights1[41][757] = 16'b1111111111111100;
    assign weights1[41][758] = 16'b1111111111111100;
    assign weights1[41][759] = 16'b1111111111110110;
    assign weights1[41][760] = 16'b1111111111110110;
    assign weights1[41][761] = 16'b1111111111110101;
    assign weights1[41][762] = 16'b1111111111110110;
    assign weights1[41][763] = 16'b1111111111101011;
    assign weights1[41][764] = 16'b1111111111011110;
    assign weights1[41][765] = 16'b1111111111011111;
    assign weights1[41][766] = 16'b1111111111100100;
    assign weights1[41][767] = 16'b1111111111100000;
    assign weights1[41][768] = 16'b1111111111011110;
    assign weights1[41][769] = 16'b1111111111110000;
    assign weights1[41][770] = 16'b1111111111111110;
    assign weights1[41][771] = 16'b1111111111110001;
    assign weights1[41][772] = 16'b1111111111110000;
    assign weights1[41][773] = 16'b1111111111110100;
    assign weights1[41][774] = 16'b1111111111111011;
    assign weights1[41][775] = 16'b1111111111111100;
    assign weights1[41][776] = 16'b1111111111111101;
    assign weights1[41][777] = 16'b1111111111111001;
    assign weights1[41][778] = 16'b1111111111111010;
    assign weights1[41][779] = 16'b1111111111111010;
    assign weights1[41][780] = 16'b1111111111111011;
    assign weights1[41][781] = 16'b1111111111111101;
    assign weights1[41][782] = 16'b1111111111111110;
    assign weights1[41][783] = 16'b0000000000000000;
    assign weights1[42][0] = 16'b0000000000000000;
    assign weights1[42][1] = 16'b0000000000000000;
    assign weights1[42][2] = 16'b1111111111111111;
    assign weights1[42][3] = 16'b1111111111111111;
    assign weights1[42][4] = 16'b1111111111111111;
    assign weights1[42][5] = 16'b1111111111111110;
    assign weights1[42][6] = 16'b1111111111111110;
    assign weights1[42][7] = 16'b1111111111111010;
    assign weights1[42][8] = 16'b1111111111110110;
    assign weights1[42][9] = 16'b1111111111101110;
    assign weights1[42][10] = 16'b1111111111110000;
    assign weights1[42][11] = 16'b1111111111110111;
    assign weights1[42][12] = 16'b1111111111110110;
    assign weights1[42][13] = 16'b1111111111110000;
    assign weights1[42][14] = 16'b1111111111101111;
    assign weights1[42][15] = 16'b1111111111101111;
    assign weights1[42][16] = 16'b1111111111111011;
    assign weights1[42][17] = 16'b1111111111111000;
    assign weights1[42][18] = 16'b1111111111110110;
    assign weights1[42][19] = 16'b1111111111110110;
    assign weights1[42][20] = 16'b1111111111111000;
    assign weights1[42][21] = 16'b1111111111110111;
    assign weights1[42][22] = 16'b1111111111111101;
    assign weights1[42][23] = 16'b1111111111111110;
    assign weights1[42][24] = 16'b1111111111111110;
    assign weights1[42][25] = 16'b1111111111111111;
    assign weights1[42][26] = 16'b0000000000000000;
    assign weights1[42][27] = 16'b0000000000000000;
    assign weights1[42][28] = 16'b0000000000000000;
    assign weights1[42][29] = 16'b0000000000000000;
    assign weights1[42][30] = 16'b0000000000000000;
    assign weights1[42][31] = 16'b1111111111111111;
    assign weights1[42][32] = 16'b0000000000000000;
    assign weights1[42][33] = 16'b1111111111111111;
    assign weights1[42][34] = 16'b1111111111111001;
    assign weights1[42][35] = 16'b1111111111110100;
    assign weights1[42][36] = 16'b1111111111101100;
    assign weights1[42][37] = 16'b1111111111100011;
    assign weights1[42][38] = 16'b1111111111011111;
    assign weights1[42][39] = 16'b1111111111110001;
    assign weights1[42][40] = 16'b1111111111110010;
    assign weights1[42][41] = 16'b1111111111100111;
    assign weights1[42][42] = 16'b1111111111011100;
    assign weights1[42][43] = 16'b1111111111100011;
    assign weights1[42][44] = 16'b1111111111101010;
    assign weights1[42][45] = 16'b1111111111101110;
    assign weights1[42][46] = 16'b1111111111101100;
    assign weights1[42][47] = 16'b1111111111110010;
    assign weights1[42][48] = 16'b1111111111110101;
    assign weights1[42][49] = 16'b1111111111110111;
    assign weights1[42][50] = 16'b1111111111111100;
    assign weights1[42][51] = 16'b1111111111111100;
    assign weights1[42][52] = 16'b1111111111111011;
    assign weights1[42][53] = 16'b1111111111111111;
    assign weights1[42][54] = 16'b1111111111111110;
    assign weights1[42][55] = 16'b1111111111111110;
    assign weights1[42][56] = 16'b0000000000000000;
    assign weights1[42][57] = 16'b0000000000000000;
    assign weights1[42][58] = 16'b0000000000000000;
    assign weights1[42][59] = 16'b1111111111111111;
    assign weights1[42][60] = 16'b1111111111111111;
    assign weights1[42][61] = 16'b1111111111111011;
    assign weights1[42][62] = 16'b1111111111110100;
    assign weights1[42][63] = 16'b1111111111101111;
    assign weights1[42][64] = 16'b1111111111101000;
    assign weights1[42][65] = 16'b1111111111100010;
    assign weights1[42][66] = 16'b1111111111011011;
    assign weights1[42][67] = 16'b1111111111010100;
    assign weights1[42][68] = 16'b1111111111101100;
    assign weights1[42][69] = 16'b1111111111011111;
    assign weights1[42][70] = 16'b1111111111001110;
    assign weights1[42][71] = 16'b1111111111010111;
    assign weights1[42][72] = 16'b1111111111100001;
    assign weights1[42][73] = 16'b1111111111101111;
    assign weights1[42][74] = 16'b1111111111101101;
    assign weights1[42][75] = 16'b1111111111101010;
    assign weights1[42][76] = 16'b1111111111101011;
    assign weights1[42][77] = 16'b1111111111101000;
    assign weights1[42][78] = 16'b1111111111101100;
    assign weights1[42][79] = 16'b1111111111110101;
    assign weights1[42][80] = 16'b1111111111111010;
    assign weights1[42][81] = 16'b1111111111111110;
    assign weights1[42][82] = 16'b0000000000000010;
    assign weights1[42][83] = 16'b1111111111111101;
    assign weights1[42][84] = 16'b0000000000000000;
    assign weights1[42][85] = 16'b1111111111111111;
    assign weights1[42][86] = 16'b1111111111111101;
    assign weights1[42][87] = 16'b1111111111111111;
    assign weights1[42][88] = 16'b1111111111111011;
    assign weights1[42][89] = 16'b1111111111111100;
    assign weights1[42][90] = 16'b1111111111101110;
    assign weights1[42][91] = 16'b1111111111100111;
    assign weights1[42][92] = 16'b1111111111101011;
    assign weights1[42][93] = 16'b1111111111001111;
    assign weights1[42][94] = 16'b1111111111001011;
    assign weights1[42][95] = 16'b1111111111001111;
    assign weights1[42][96] = 16'b1111111111101101;
    assign weights1[42][97] = 16'b1111111111001100;
    assign weights1[42][98] = 16'b1111111111001001;
    assign weights1[42][99] = 16'b1111111110110011;
    assign weights1[42][100] = 16'b1111111111010101;
    assign weights1[42][101] = 16'b1111111111001011;
    assign weights1[42][102] = 16'b1111111111001001;
    assign weights1[42][103] = 16'b1111111111010001;
    assign weights1[42][104] = 16'b1111111111011111;
    assign weights1[42][105] = 16'b1111111111100000;
    assign weights1[42][106] = 16'b1111111111101001;
    assign weights1[42][107] = 16'b1111111111101111;
    assign weights1[42][108] = 16'b1111111111110110;
    assign weights1[42][109] = 16'b0000000000000000;
    assign weights1[42][110] = 16'b0000000000000011;
    assign weights1[42][111] = 16'b1111111111111110;
    assign weights1[42][112] = 16'b1111111111111111;
    assign weights1[42][113] = 16'b1111111111111011;
    assign weights1[42][114] = 16'b1111111111111100;
    assign weights1[42][115] = 16'b1111111111111011;
    assign weights1[42][116] = 16'b1111111111111110;
    assign weights1[42][117] = 16'b1111111111110101;
    assign weights1[42][118] = 16'b1111111111101110;
    assign weights1[42][119] = 16'b1111111111010010;
    assign weights1[42][120] = 16'b1111111111010110;
    assign weights1[42][121] = 16'b1111111110110111;
    assign weights1[42][122] = 16'b1111111110111110;
    assign weights1[42][123] = 16'b1111111111000001;
    assign weights1[42][124] = 16'b1111111111010001;
    assign weights1[42][125] = 16'b1111111111010111;
    assign weights1[42][126] = 16'b1111111111010100;
    assign weights1[42][127] = 16'b1111111111001101;
    assign weights1[42][128] = 16'b1111111111111101;
    assign weights1[42][129] = 16'b1111111111101101;
    assign weights1[42][130] = 16'b1111111111011110;
    assign weights1[42][131] = 16'b1111111111011000;
    assign weights1[42][132] = 16'b1111111111011000;
    assign weights1[42][133] = 16'b1111111111101100;
    assign weights1[42][134] = 16'b1111111111111001;
    assign weights1[42][135] = 16'b1111111111111100;
    assign weights1[42][136] = 16'b0000000000000001;
    assign weights1[42][137] = 16'b0000000000000101;
    assign weights1[42][138] = 16'b0000000000000011;
    assign weights1[42][139] = 16'b1111111111111101;
    assign weights1[42][140] = 16'b1111111111111101;
    assign weights1[42][141] = 16'b1111111111111010;
    assign weights1[42][142] = 16'b1111111111111011;
    assign weights1[42][143] = 16'b1111111111111001;
    assign weights1[42][144] = 16'b1111111111110111;
    assign weights1[42][145] = 16'b1111111111101111;
    assign weights1[42][146] = 16'b1111111111111010;
    assign weights1[42][147] = 16'b1111111111101010;
    assign weights1[42][148] = 16'b1111111111101000;
    assign weights1[42][149] = 16'b1111111111011001;
    assign weights1[42][150] = 16'b1111111111101110;
    assign weights1[42][151] = 16'b1111111111000101;
    assign weights1[42][152] = 16'b1111111111011010;
    assign weights1[42][153] = 16'b1111111111011011;
    assign weights1[42][154] = 16'b1111111111110001;
    assign weights1[42][155] = 16'b1111111111101001;
    assign weights1[42][156] = 16'b1111111111101000;
    assign weights1[42][157] = 16'b1111111111101011;
    assign weights1[42][158] = 16'b1111111111110100;
    assign weights1[42][159] = 16'b1111111111100110;
    assign weights1[42][160] = 16'b1111111111110001;
    assign weights1[42][161] = 16'b1111111111101100;
    assign weights1[42][162] = 16'b1111111111111000;
    assign weights1[42][163] = 16'b1111111111111100;
    assign weights1[42][164] = 16'b0000000000001100;
    assign weights1[42][165] = 16'b0000000000000110;
    assign weights1[42][166] = 16'b1111111111111010;
    assign weights1[42][167] = 16'b1111111111111011;
    assign weights1[42][168] = 16'b1111111111111100;
    assign weights1[42][169] = 16'b1111111111110111;
    assign weights1[42][170] = 16'b1111111111110000;
    assign weights1[42][171] = 16'b1111111111101110;
    assign weights1[42][172] = 16'b1111111111110110;
    assign weights1[42][173] = 16'b1111111111111101;
    assign weights1[42][174] = 16'b1111111111111000;
    assign weights1[42][175] = 16'b0000000000000010;
    assign weights1[42][176] = 16'b0000000000010100;
    assign weights1[42][177] = 16'b1111111111011110;
    assign weights1[42][178] = 16'b0000000000010100;
    assign weights1[42][179] = 16'b1111111111110001;
    assign weights1[42][180] = 16'b0000000000010010;
    assign weights1[42][181] = 16'b0000000000010001;
    assign weights1[42][182] = 16'b1111111111100110;
    assign weights1[42][183] = 16'b1111111111111001;
    assign weights1[42][184] = 16'b1111111111101110;
    assign weights1[42][185] = 16'b1111111111110000;
    assign weights1[42][186] = 16'b0000000000010100;
    assign weights1[42][187] = 16'b0000000000001000;
    assign weights1[42][188] = 16'b1111111111111010;
    assign weights1[42][189] = 16'b0000000000001010;
    assign weights1[42][190] = 16'b0000000000001001;
    assign weights1[42][191] = 16'b0000000000010011;
    assign weights1[42][192] = 16'b0000000000010110;
    assign weights1[42][193] = 16'b1111111111111100;
    assign weights1[42][194] = 16'b1111111111111011;
    assign weights1[42][195] = 16'b1111111111111101;
    assign weights1[42][196] = 16'b1111111111111011;
    assign weights1[42][197] = 16'b1111111111110111;
    assign weights1[42][198] = 16'b1111111111101101;
    assign weights1[42][199] = 16'b1111111111101100;
    assign weights1[42][200] = 16'b1111111111101011;
    assign weights1[42][201] = 16'b1111111111101000;
    assign weights1[42][202] = 16'b1111111111111000;
    assign weights1[42][203] = 16'b0000000000010000;
    assign weights1[42][204] = 16'b0000000000001111;
    assign weights1[42][205] = 16'b0000000000010000;
    assign weights1[42][206] = 16'b0000000000010110;
    assign weights1[42][207] = 16'b0000000000011101;
    assign weights1[42][208] = 16'b0000000000100000;
    assign weights1[42][209] = 16'b1111111111111000;
    assign weights1[42][210] = 16'b1111111111111000;
    assign weights1[42][211] = 16'b1111111111111000;
    assign weights1[42][212] = 16'b0000000000000110;
    assign weights1[42][213] = 16'b1111111111111000;
    assign weights1[42][214] = 16'b0000000000010010;
    assign weights1[42][215] = 16'b0000000000010100;
    assign weights1[42][216] = 16'b0000000000000000;
    assign weights1[42][217] = 16'b0000000000010001;
    assign weights1[42][218] = 16'b0000000000010001;
    assign weights1[42][219] = 16'b0000000000010101;
    assign weights1[42][220] = 16'b0000000000001101;
    assign weights1[42][221] = 16'b0000000000001001;
    assign weights1[42][222] = 16'b1111111111111110;
    assign weights1[42][223] = 16'b0000000000000001;
    assign weights1[42][224] = 16'b1111111111111010;
    assign weights1[42][225] = 16'b1111111111110010;
    assign weights1[42][226] = 16'b1111111111101101;
    assign weights1[42][227] = 16'b1111111111011110;
    assign weights1[42][228] = 16'b1111111111001001;
    assign weights1[42][229] = 16'b1111111111110011;
    assign weights1[42][230] = 16'b1111111111010100;
    assign weights1[42][231] = 16'b0000000000000010;
    assign weights1[42][232] = 16'b0000000000011101;
    assign weights1[42][233] = 16'b1111111111111101;
    assign weights1[42][234] = 16'b0000000000011010;
    assign weights1[42][235] = 16'b0000000000110001;
    assign weights1[42][236] = 16'b0000000000110000;
    assign weights1[42][237] = 16'b0000000000010000;
    assign weights1[42][238] = 16'b0000000000010011;
    assign weights1[42][239] = 16'b0000000000001101;
    assign weights1[42][240] = 16'b0000000000010010;
    assign weights1[42][241] = 16'b0000000000010010;
    assign weights1[42][242] = 16'b0000000000010000;
    assign weights1[42][243] = 16'b0000000000000010;
    assign weights1[42][244] = 16'b0000000000100000;
    assign weights1[42][245] = 16'b0000000000000011;
    assign weights1[42][246] = 16'b1111111111110111;
    assign weights1[42][247] = 16'b0000000000001110;
    assign weights1[42][248] = 16'b0000000000000110;
    assign weights1[42][249] = 16'b0000000000000110;
    assign weights1[42][250] = 16'b0000000000000011;
    assign weights1[42][251] = 16'b1111111111111010;
    assign weights1[42][252] = 16'b1111111111111000;
    assign weights1[42][253] = 16'b1111111111110110;
    assign weights1[42][254] = 16'b1111111111101011;
    assign weights1[42][255] = 16'b1111111111101011;
    assign weights1[42][256] = 16'b1111111111101111;
    assign weights1[42][257] = 16'b0000000000000000;
    assign weights1[42][258] = 16'b0000000000001101;
    assign weights1[42][259] = 16'b1111111111110100;
    assign weights1[42][260] = 16'b0000000000100011;
    assign weights1[42][261] = 16'b0000000000011111;
    assign weights1[42][262] = 16'b0000000000111110;
    assign weights1[42][263] = 16'b0000000000101010;
    assign weights1[42][264] = 16'b0000000000011001;
    assign weights1[42][265] = 16'b0000000000110001;
    assign weights1[42][266] = 16'b0000000000101100;
    assign weights1[42][267] = 16'b0000000000011010;
    assign weights1[42][268] = 16'b1111111111110010;
    assign weights1[42][269] = 16'b0000000000010110;
    assign weights1[42][270] = 16'b0000000000011100;
    assign weights1[42][271] = 16'b0000000000010100;
    assign weights1[42][272] = 16'b0000000000101110;
    assign weights1[42][273] = 16'b0000000000011001;
    assign weights1[42][274] = 16'b0000000000010011;
    assign weights1[42][275] = 16'b0000000000000000;
    assign weights1[42][276] = 16'b0000000000000100;
    assign weights1[42][277] = 16'b0000000000000000;
    assign weights1[42][278] = 16'b1111111111101110;
    assign weights1[42][279] = 16'b0000000000010001;
    assign weights1[42][280] = 16'b1111111111111010;
    assign weights1[42][281] = 16'b1111111111101111;
    assign weights1[42][282] = 16'b1111111111110010;
    assign weights1[42][283] = 16'b1111111111110001;
    assign weights1[42][284] = 16'b0000000000000001;
    assign weights1[42][285] = 16'b1111111111111011;
    assign weights1[42][286] = 16'b0000000000000011;
    assign weights1[42][287] = 16'b0000000000000110;
    assign weights1[42][288] = 16'b0000000000001101;
    assign weights1[42][289] = 16'b0000000000010111;
    assign weights1[42][290] = 16'b0000000000000001;
    assign weights1[42][291] = 16'b0000000000110100;
    assign weights1[42][292] = 16'b0000000000101010;
    assign weights1[42][293] = 16'b0000000000111100;
    assign weights1[42][294] = 16'b0000000000110000;
    assign weights1[42][295] = 16'b0000000000101110;
    assign weights1[42][296] = 16'b0000000000001011;
    assign weights1[42][297] = 16'b0000000000101110;
    assign weights1[42][298] = 16'b0000000000000001;
    assign weights1[42][299] = 16'b0000000000001101;
    assign weights1[42][300] = 16'b0000000000001001;
    assign weights1[42][301] = 16'b0000000000011011;
    assign weights1[42][302] = 16'b0000000000011101;
    assign weights1[42][303] = 16'b0000000000000001;
    assign weights1[42][304] = 16'b0000000000000100;
    assign weights1[42][305] = 16'b0000000000000001;
    assign weights1[42][306] = 16'b0000000000000110;
    assign weights1[42][307] = 16'b0000000000010001;
    assign weights1[42][308] = 16'b1111111111111001;
    assign weights1[42][309] = 16'b1111111111110111;
    assign weights1[42][310] = 16'b1111111111110111;
    assign weights1[42][311] = 16'b1111111111111000;
    assign weights1[42][312] = 16'b1111111111101101;
    assign weights1[42][313] = 16'b1111111111101111;
    assign weights1[42][314] = 16'b1111111111111101;
    assign weights1[42][315] = 16'b1111111111111000;
    assign weights1[42][316] = 16'b1111111111101000;
    assign weights1[42][317] = 16'b0000000000001100;
    assign weights1[42][318] = 16'b0000000000100010;
    assign weights1[42][319] = 16'b0000000000011100;
    assign weights1[42][320] = 16'b0000000000010100;
    assign weights1[42][321] = 16'b1111111111110001;
    assign weights1[42][322] = 16'b1111111111101010;
    assign weights1[42][323] = 16'b0000000000001110;
    assign weights1[42][324] = 16'b1111111111111000;
    assign weights1[42][325] = 16'b0000000000010001;
    assign weights1[42][326] = 16'b0000000000100010;
    assign weights1[42][327] = 16'b0000000000001111;
    assign weights1[42][328] = 16'b0000000000100101;
    assign weights1[42][329] = 16'b0000000000000010;
    assign weights1[42][330] = 16'b0000000000011111;
    assign weights1[42][331] = 16'b0000000000000111;
    assign weights1[42][332] = 16'b1111111111111011;
    assign weights1[42][333] = 16'b1111111111101000;
    assign weights1[42][334] = 16'b0000000000000101;
    assign weights1[42][335] = 16'b0000000000010111;
    assign weights1[42][336] = 16'b1111111111111100;
    assign weights1[42][337] = 16'b0000000000000010;
    assign weights1[42][338] = 16'b0000000000000011;
    assign weights1[42][339] = 16'b1111111111101111;
    assign weights1[42][340] = 16'b1111111111110111;
    assign weights1[42][341] = 16'b1111111111101001;
    assign weights1[42][342] = 16'b0000000000001001;
    assign weights1[42][343] = 16'b1111111111110100;
    assign weights1[42][344] = 16'b1111111111111011;
    assign weights1[42][345] = 16'b0000000000000101;
    assign weights1[42][346] = 16'b0000000000001001;
    assign weights1[42][347] = 16'b0000000000001111;
    assign weights1[42][348] = 16'b0000000000000010;
    assign weights1[42][349] = 16'b1111111110110111;
    assign weights1[42][350] = 16'b1111111110111100;
    assign weights1[42][351] = 16'b1111111111010110;
    assign weights1[42][352] = 16'b1111111111110010;
    assign weights1[42][353] = 16'b1111111111111111;
    assign weights1[42][354] = 16'b1111111111110100;
    assign weights1[42][355] = 16'b1111111111110000;
    assign weights1[42][356] = 16'b0000000000001011;
    assign weights1[42][357] = 16'b1111111111110101;
    assign weights1[42][358] = 16'b0000000000001110;
    assign weights1[42][359] = 16'b0000000000000101;
    assign weights1[42][360] = 16'b0000000000000010;
    assign weights1[42][361] = 16'b1111111111101010;
    assign weights1[42][362] = 16'b1111111111111100;
    assign weights1[42][363] = 16'b0000000000001111;
    assign weights1[42][364] = 16'b1111111111111101;
    assign weights1[42][365] = 16'b0000000000001000;
    assign weights1[42][366] = 16'b1111111111111001;
    assign weights1[42][367] = 16'b1111111111110010;
    assign weights1[42][368] = 16'b1111111111111101;
    assign weights1[42][369] = 16'b1111111111111100;
    assign weights1[42][370] = 16'b1111111111111001;
    assign weights1[42][371] = 16'b0000000000000011;
    assign weights1[42][372] = 16'b0000000000010011;
    assign weights1[42][373] = 16'b0000000000001000;
    assign weights1[42][374] = 16'b0000000000001110;
    assign weights1[42][375] = 16'b0000000000000100;
    assign weights1[42][376] = 16'b1111111111001111;
    assign weights1[42][377] = 16'b1111111110000001;
    assign weights1[42][378] = 16'b1111111110001010;
    assign weights1[42][379] = 16'b1111111111010011;
    assign weights1[42][380] = 16'b1111111111101101;
    assign weights1[42][381] = 16'b0000000000000100;
    assign weights1[42][382] = 16'b1111111111010110;
    assign weights1[42][383] = 16'b0000000000000111;
    assign weights1[42][384] = 16'b1111111111111001;
    assign weights1[42][385] = 16'b1111111111111100;
    assign weights1[42][386] = 16'b0000000000000001;
    assign weights1[42][387] = 16'b1111111111111010;
    assign weights1[42][388] = 16'b1111111111111100;
    assign weights1[42][389] = 16'b1111111111101111;
    assign weights1[42][390] = 16'b0000000000000000;
    assign weights1[42][391] = 16'b0000000000000111;
    assign weights1[42][392] = 16'b0000000000000110;
    assign weights1[42][393] = 16'b0000000000001011;
    assign weights1[42][394] = 16'b1111111111110101;
    assign weights1[42][395] = 16'b1111111111111011;
    assign weights1[42][396] = 16'b1111111111110010;
    assign weights1[42][397] = 16'b0000000000100110;
    assign weights1[42][398] = 16'b0000000000000100;
    assign weights1[42][399] = 16'b0000000000010101;
    assign weights1[42][400] = 16'b0000000000000001;
    assign weights1[42][401] = 16'b1111111111111100;
    assign weights1[42][402] = 16'b0000000000011100;
    assign weights1[42][403] = 16'b0000000000000110;
    assign weights1[42][404] = 16'b1111111110100011;
    assign weights1[42][405] = 16'b1111111101011011;
    assign weights1[42][406] = 16'b1111111111010010;
    assign weights1[42][407] = 16'b1111111111101111;
    assign weights1[42][408] = 16'b1111111111110000;
    assign weights1[42][409] = 16'b1111111111010110;
    assign weights1[42][410] = 16'b1111111111011101;
    assign weights1[42][411] = 16'b1111111111011111;
    assign weights1[42][412] = 16'b1111111111110110;
    assign weights1[42][413] = 16'b1111111111101101;
    assign weights1[42][414] = 16'b1111111111111111;
    assign weights1[42][415] = 16'b0000000000000111;
    assign weights1[42][416] = 16'b0000000000001000;
    assign weights1[42][417] = 16'b1111111111100001;
    assign weights1[42][418] = 16'b1111111111111011;
    assign weights1[42][419] = 16'b0000000000000000;
    assign weights1[42][420] = 16'b0000000000001000;
    assign weights1[42][421] = 16'b0000000000001100;
    assign weights1[42][422] = 16'b1111111111111000;
    assign weights1[42][423] = 16'b0000000000000011;
    assign weights1[42][424] = 16'b0000000000000000;
    assign weights1[42][425] = 16'b0000000000010010;
    assign weights1[42][426] = 16'b0000000000100001;
    assign weights1[42][427] = 16'b0000000000011101;
    assign weights1[42][428] = 16'b0000000000000100;
    assign weights1[42][429] = 16'b0000000000010000;
    assign weights1[42][430] = 16'b0000000000101100;
    assign weights1[42][431] = 16'b1111111111011100;
    assign weights1[42][432] = 16'b1111111101101111;
    assign weights1[42][433] = 16'b1111111100111110;
    assign weights1[42][434] = 16'b1111111111011011;
    assign weights1[42][435] = 16'b1111111111111011;
    assign weights1[42][436] = 16'b1111111111101010;
    assign weights1[42][437] = 16'b1111111111010101;
    assign weights1[42][438] = 16'b1111111111101001;
    assign weights1[42][439] = 16'b1111111111011101;
    assign weights1[42][440] = 16'b1111111111100011;
    assign weights1[42][441] = 16'b1111111111111110;
    assign weights1[42][442] = 16'b1111111111101010;
    assign weights1[42][443] = 16'b1111111111110011;
    assign weights1[42][444] = 16'b1111111111111100;
    assign weights1[42][445] = 16'b1111111111110000;
    assign weights1[42][446] = 16'b1111111111110000;
    assign weights1[42][447] = 16'b1111111111111111;
    assign weights1[42][448] = 16'b0000000000001100;
    assign weights1[42][449] = 16'b0000000000001100;
    assign weights1[42][450] = 16'b0000000000000111;
    assign weights1[42][451] = 16'b0000000000010001;
    assign weights1[42][452] = 16'b1111111111110101;
    assign weights1[42][453] = 16'b0000000000001110;
    assign weights1[42][454] = 16'b0000000000010010;
    assign weights1[42][455] = 16'b1111111111111100;
    assign weights1[42][456] = 16'b0000000000100000;
    assign weights1[42][457] = 16'b0000000000000111;
    assign weights1[42][458] = 16'b0000000000010100;
    assign weights1[42][459] = 16'b1111111110101000;
    assign weights1[42][460] = 16'b1111111101001100;
    assign weights1[42][461] = 16'b1111111110011101;
    assign weights1[42][462] = 16'b1111111111101010;
    assign weights1[42][463] = 16'b1111111111101101;
    assign weights1[42][464] = 16'b1111111111010101;
    assign weights1[42][465] = 16'b1111111111011111;
    assign weights1[42][466] = 16'b1111111111101100;
    assign weights1[42][467] = 16'b1111111111111101;
    assign weights1[42][468] = 16'b1111111111101111;
    assign weights1[42][469] = 16'b0000000000001001;
    assign weights1[42][470] = 16'b1111111111101101;
    assign weights1[42][471] = 16'b1111111111101011;
    assign weights1[42][472] = 16'b0000000000000001;
    assign weights1[42][473] = 16'b1111111111101101;
    assign weights1[42][474] = 16'b1111111111110111;
    assign weights1[42][475] = 16'b1111111111111101;
    assign weights1[42][476] = 16'b0000000000001010;
    assign weights1[42][477] = 16'b0000000000001100;
    assign weights1[42][478] = 16'b0000000000001110;
    assign weights1[42][479] = 16'b1111111111111101;
    assign weights1[42][480] = 16'b0000000000001000;
    assign weights1[42][481] = 16'b0000000000000111;
    assign weights1[42][482] = 16'b0000000000001010;
    assign weights1[42][483] = 16'b0000000000001100;
    assign weights1[42][484] = 16'b0000000000000000;
    assign weights1[42][485] = 16'b1111111111111111;
    assign weights1[42][486] = 16'b1111111111001010;
    assign weights1[42][487] = 16'b1111111101110000;
    assign weights1[42][488] = 16'b1111111101000101;
    assign weights1[42][489] = 16'b1111111111101111;
    assign weights1[42][490] = 16'b0000000000000011;
    assign weights1[42][491] = 16'b1111111111011100;
    assign weights1[42][492] = 16'b1111111111011101;
    assign weights1[42][493] = 16'b0000000000000010;
    assign weights1[42][494] = 16'b1111111111110110;
    assign weights1[42][495] = 16'b1111111111101100;
    assign weights1[42][496] = 16'b0000000000000000;
    assign weights1[42][497] = 16'b1111111111110000;
    assign weights1[42][498] = 16'b0000000000000011;
    assign weights1[42][499] = 16'b1111111111111011;
    assign weights1[42][500] = 16'b1111111111111000;
    assign weights1[42][501] = 16'b1111111111101010;
    assign weights1[42][502] = 16'b1111111111110110;
    assign weights1[42][503] = 16'b1111111111111011;
    assign weights1[42][504] = 16'b0000000000001110;
    assign weights1[42][505] = 16'b0000000000011100;
    assign weights1[42][506] = 16'b0000000000010100;
    assign weights1[42][507] = 16'b0000000000001110;
    assign weights1[42][508] = 16'b0000000000000111;
    assign weights1[42][509] = 16'b0000000000001110;
    assign weights1[42][510] = 16'b0000000000000111;
    assign weights1[42][511] = 16'b0000000000000010;
    assign weights1[42][512] = 16'b1111111111110011;
    assign weights1[42][513] = 16'b0000000000000010;
    assign weights1[42][514] = 16'b1111111111010100;
    assign weights1[42][515] = 16'b1111111101101101;
    assign weights1[42][516] = 16'b1111111110110000;
    assign weights1[42][517] = 16'b1111111111101111;
    assign weights1[42][518] = 16'b0000000000000111;
    assign weights1[42][519] = 16'b1111111111101111;
    assign weights1[42][520] = 16'b0000000000001011;
    assign weights1[42][521] = 16'b0000000000010000;
    assign weights1[42][522] = 16'b0000000000000011;
    assign weights1[42][523] = 16'b1111111111111111;
    assign weights1[42][524] = 16'b1111111111111001;
    assign weights1[42][525] = 16'b0000000000011110;
    assign weights1[42][526] = 16'b1111111111111110;
    assign weights1[42][527] = 16'b1111111111101111;
    assign weights1[42][528] = 16'b1111111111101110;
    assign weights1[42][529] = 16'b1111111111100011;
    assign weights1[42][530] = 16'b1111111111111000;
    assign weights1[42][531] = 16'b1111111111111111;
    assign weights1[42][532] = 16'b0000000000010011;
    assign weights1[42][533] = 16'b0000000000001010;
    assign weights1[42][534] = 16'b0000000000010000;
    assign weights1[42][535] = 16'b0000000000000001;
    assign weights1[42][536] = 16'b1111111111110100;
    assign weights1[42][537] = 16'b0000000000000100;
    assign weights1[42][538] = 16'b0000000000000100;
    assign weights1[42][539] = 16'b1111111111111001;
    assign weights1[42][540] = 16'b1111111111110110;
    assign weights1[42][541] = 16'b1111111111110011;
    assign weights1[42][542] = 16'b1111111111011110;
    assign weights1[42][543] = 16'b1111111110101100;
    assign weights1[42][544] = 16'b1111111111001111;
    assign weights1[42][545] = 16'b1111111111100111;
    assign weights1[42][546] = 16'b0000000000001101;
    assign weights1[42][547] = 16'b0000000000001010;
    assign weights1[42][548] = 16'b0000000000000011;
    assign weights1[42][549] = 16'b1111111111111101;
    assign weights1[42][550] = 16'b0000000000010010;
    assign weights1[42][551] = 16'b1111111111101101;
    assign weights1[42][552] = 16'b0000000000000010;
    assign weights1[42][553] = 16'b0000000000001111;
    assign weights1[42][554] = 16'b1111111111101101;
    assign weights1[42][555] = 16'b1111111111100110;
    assign weights1[42][556] = 16'b1111111111100010;
    assign weights1[42][557] = 16'b1111111111101001;
    assign weights1[42][558] = 16'b1111111111111001;
    assign weights1[42][559] = 16'b0000000000000100;
    assign weights1[42][560] = 16'b0000000000010100;
    assign weights1[42][561] = 16'b0000000000001111;
    assign weights1[42][562] = 16'b0000000000000111;
    assign weights1[42][563] = 16'b0000000000000011;
    assign weights1[42][564] = 16'b0000000000010100;
    assign weights1[42][565] = 16'b0000000000000111;
    assign weights1[42][566] = 16'b0000000000011010;
    assign weights1[42][567] = 16'b0000000000000000;
    assign weights1[42][568] = 16'b1111111111111010;
    assign weights1[42][569] = 16'b1111111111101111;
    assign weights1[42][570] = 16'b1111111111110011;
    assign weights1[42][571] = 16'b0000000000000001;
    assign weights1[42][572] = 16'b1111111111110111;
    assign weights1[42][573] = 16'b1111111111101010;
    assign weights1[42][574] = 16'b0000000000000010;
    assign weights1[42][575] = 16'b1111111111111100;
    assign weights1[42][576] = 16'b1111111111101101;
    assign weights1[42][577] = 16'b1111111111111000;
    assign weights1[42][578] = 16'b1111111111100011;
    assign weights1[42][579] = 16'b0000000000001111;
    assign weights1[42][580] = 16'b1111111111101001;
    assign weights1[42][581] = 16'b1111111111101111;
    assign weights1[42][582] = 16'b1111111111110001;
    assign weights1[42][583] = 16'b1111111111101101;
    assign weights1[42][584] = 16'b1111111111101101;
    assign weights1[42][585] = 16'b1111111111101100;
    assign weights1[42][586] = 16'b1111111111110011;
    assign weights1[42][587] = 16'b1111111111111101;
    assign weights1[42][588] = 16'b0000000000001101;
    assign weights1[42][589] = 16'b0000000000000111;
    assign weights1[42][590] = 16'b0000000000000011;
    assign weights1[42][591] = 16'b0000000000001011;
    assign weights1[42][592] = 16'b0000000000010001;
    assign weights1[42][593] = 16'b0000000000010100;
    assign weights1[42][594] = 16'b1111111111111110;
    assign weights1[42][595] = 16'b0000000000000110;
    assign weights1[42][596] = 16'b1111111111101101;
    assign weights1[42][597] = 16'b0000000000001011;
    assign weights1[42][598] = 16'b0000000000010101;
    assign weights1[42][599] = 16'b0000000000010100;
    assign weights1[42][600] = 16'b0000000000000010;
    assign weights1[42][601] = 16'b0000000000000100;
    assign weights1[42][602] = 16'b1111111111101101;
    assign weights1[42][603] = 16'b0000000000001101;
    assign weights1[42][604] = 16'b0000000000000001;
    assign weights1[42][605] = 16'b1111111111111001;
    assign weights1[42][606] = 16'b1111111111101100;
    assign weights1[42][607] = 16'b1111111111010010;
    assign weights1[42][608] = 16'b1111111111110010;
    assign weights1[42][609] = 16'b1111111111110100;
    assign weights1[42][610] = 16'b1111111111010101;
    assign weights1[42][611] = 16'b1111111111100010;
    assign weights1[42][612] = 16'b1111111111101010;
    assign weights1[42][613] = 16'b1111111111101110;
    assign weights1[42][614] = 16'b1111111111110110;
    assign weights1[42][615] = 16'b1111111111111100;
    assign weights1[42][616] = 16'b0000000000000111;
    assign weights1[42][617] = 16'b0000000000001001;
    assign weights1[42][618] = 16'b0000000000000010;
    assign weights1[42][619] = 16'b0000000000000111;
    assign weights1[42][620] = 16'b1111111111101101;
    assign weights1[42][621] = 16'b0000000000000010;
    assign weights1[42][622] = 16'b0000000000011101;
    assign weights1[42][623] = 16'b1111111111110100;
    assign weights1[42][624] = 16'b0000000000100100;
    assign weights1[42][625] = 16'b0000000000110001;
    assign weights1[42][626] = 16'b0000000000001011;
    assign weights1[42][627] = 16'b1111111111111111;
    assign weights1[42][628] = 16'b0000000000001010;
    assign weights1[42][629] = 16'b0000000000011101;
    assign weights1[42][630] = 16'b0000000000010111;
    assign weights1[42][631] = 16'b0000000000000101;
    assign weights1[42][632] = 16'b1111111111111010;
    assign weights1[42][633] = 16'b0000000000000101;
    assign weights1[42][634] = 16'b0000000000010011;
    assign weights1[42][635] = 16'b1111111111111000;
    assign weights1[42][636] = 16'b1111111111101000;
    assign weights1[42][637] = 16'b1111111111101100;
    assign weights1[42][638] = 16'b1111111111101011;
    assign weights1[42][639] = 16'b1111111111101101;
    assign weights1[42][640] = 16'b1111111111100101;
    assign weights1[42][641] = 16'b1111111111101100;
    assign weights1[42][642] = 16'b1111111111111010;
    assign weights1[42][643] = 16'b1111111111111100;
    assign weights1[42][644] = 16'b0000000000000101;
    assign weights1[42][645] = 16'b0000000000000010;
    assign weights1[42][646] = 16'b1111111111111100;
    assign weights1[42][647] = 16'b0000000000000100;
    assign weights1[42][648] = 16'b0000000000001111;
    assign weights1[42][649] = 16'b0000000000000100;
    assign weights1[42][650] = 16'b0000000000100010;
    assign weights1[42][651] = 16'b0000000000100111;
    assign weights1[42][652] = 16'b0000000000000001;
    assign weights1[42][653] = 16'b1111111111111111;
    assign weights1[42][654] = 16'b0000000000100001;
    assign weights1[42][655] = 16'b0000000000000000;
    assign weights1[42][656] = 16'b0000000000000101;
    assign weights1[42][657] = 16'b0000000000010000;
    assign weights1[42][658] = 16'b0000000000001101;
    assign weights1[42][659] = 16'b0000000000011001;
    assign weights1[42][660] = 16'b0000000000000001;
    assign weights1[42][661] = 16'b0000000000101010;
    assign weights1[42][662] = 16'b0000000000000001;
    assign weights1[42][663] = 16'b0000000000000001;
    assign weights1[42][664] = 16'b1111111111101110;
    assign weights1[42][665] = 16'b0000000000000101;
    assign weights1[42][666] = 16'b1111111111110010;
    assign weights1[42][667] = 16'b1111111111110111;
    assign weights1[42][668] = 16'b1111111111110010;
    assign weights1[42][669] = 16'b1111111111111000;
    assign weights1[42][670] = 16'b1111111111111111;
    assign weights1[42][671] = 16'b1111111111111111;
    assign weights1[42][672] = 16'b1111111111111011;
    assign weights1[42][673] = 16'b0000000000000111;
    assign weights1[42][674] = 16'b1111111111110011;
    assign weights1[42][675] = 16'b0000000000000011;
    assign weights1[42][676] = 16'b0000000000001111;
    assign weights1[42][677] = 16'b0000000000011101;
    assign weights1[42][678] = 16'b0000000000100011;
    assign weights1[42][679] = 16'b0000000000001101;
    assign weights1[42][680] = 16'b0000000000011011;
    assign weights1[42][681] = 16'b0000000000100010;
    assign weights1[42][682] = 16'b0000000000011111;
    assign weights1[42][683] = 16'b0000000000010010;
    assign weights1[42][684] = 16'b0000000000000100;
    assign weights1[42][685] = 16'b1111111111101010;
    assign weights1[42][686] = 16'b0000000000001010;
    assign weights1[42][687] = 16'b1111111111100010;
    assign weights1[42][688] = 16'b1111111111100001;
    assign weights1[42][689] = 16'b0000000000001000;
    assign weights1[42][690] = 16'b1111111111100000;
    assign weights1[42][691] = 16'b1111111111101000;
    assign weights1[42][692] = 16'b1111111111110001;
    assign weights1[42][693] = 16'b0000000000000100;
    assign weights1[42][694] = 16'b1111111111110101;
    assign weights1[42][695] = 16'b1111111111110111;
    assign weights1[42][696] = 16'b1111111111111000;
    assign weights1[42][697] = 16'b1111111111111001;
    assign weights1[42][698] = 16'b1111111111111101;
    assign weights1[42][699] = 16'b0000000000000001;
    assign weights1[42][700] = 16'b1111111111111111;
    assign weights1[42][701] = 16'b0000000000000000;
    assign weights1[42][702] = 16'b0000000000000011;
    assign weights1[42][703] = 16'b0000000000001010;
    assign weights1[42][704] = 16'b0000000000001101;
    assign weights1[42][705] = 16'b0000000000000111;
    assign weights1[42][706] = 16'b0000000000100011;
    assign weights1[42][707] = 16'b0000000000011000;
    assign weights1[42][708] = 16'b0000000000001101;
    assign weights1[42][709] = 16'b0000000000000010;
    assign weights1[42][710] = 16'b0000000000001010;
    assign weights1[42][711] = 16'b0000000000000101;
    assign weights1[42][712] = 16'b0000000000001011;
    assign weights1[42][713] = 16'b1111111111111101;
    assign weights1[42][714] = 16'b0000000000001011;
    assign weights1[42][715] = 16'b1111111111110010;
    assign weights1[42][716] = 16'b1111111111110000;
    assign weights1[42][717] = 16'b1111111111010110;
    assign weights1[42][718] = 16'b1111111111110100;
    assign weights1[42][719] = 16'b1111111111110010;
    assign weights1[42][720] = 16'b1111111111101011;
    assign weights1[42][721] = 16'b0000000000000110;
    assign weights1[42][722] = 16'b1111111111110000;
    assign weights1[42][723] = 16'b1111111111111000;
    assign weights1[42][724] = 16'b1111111111110011;
    assign weights1[42][725] = 16'b1111111111110110;
    assign weights1[42][726] = 16'b1111111111111000;
    assign weights1[42][727] = 16'b1111111111111011;
    assign weights1[42][728] = 16'b0000000000000000;
    assign weights1[42][729] = 16'b1111111111111001;
    assign weights1[42][730] = 16'b1111111111111111;
    assign weights1[42][731] = 16'b0000000000000000;
    assign weights1[42][732] = 16'b0000000000000001;
    assign weights1[42][733] = 16'b0000000000001011;
    assign weights1[42][734] = 16'b1111111111111111;
    assign weights1[42][735] = 16'b0000000000001101;
    assign weights1[42][736] = 16'b0000000000011011;
    assign weights1[42][737] = 16'b0000000000001000;
    assign weights1[42][738] = 16'b0000000000000100;
    assign weights1[42][739] = 16'b0000000000011101;
    assign weights1[42][740] = 16'b1111111111110110;
    assign weights1[42][741] = 16'b0000000000000010;
    assign weights1[42][742] = 16'b0000000000000111;
    assign weights1[42][743] = 16'b0000000000001001;
    assign weights1[42][744] = 16'b0000000000000011;
    assign weights1[42][745] = 16'b0000000000000001;
    assign weights1[42][746] = 16'b1111111111101111;
    assign weights1[42][747] = 16'b0000000000010000;
    assign weights1[42][748] = 16'b1111111111101010;
    assign weights1[42][749] = 16'b1111111111110001;
    assign weights1[42][750] = 16'b1111111111100110;
    assign weights1[42][751] = 16'b1111111111101011;
    assign weights1[42][752] = 16'b1111111111110001;
    assign weights1[42][753] = 16'b1111111111110111;
    assign weights1[42][754] = 16'b1111111111111101;
    assign weights1[42][755] = 16'b1111111111111101;
    assign weights1[42][756] = 16'b1111111111111110;
    assign weights1[42][757] = 16'b1111111111111110;
    assign weights1[42][758] = 16'b1111111111111110;
    assign weights1[42][759] = 16'b1111111111111101;
    assign weights1[42][760] = 16'b1111111111110011;
    assign weights1[42][761] = 16'b1111111111110011;
    assign weights1[42][762] = 16'b1111111111110000;
    assign weights1[42][763] = 16'b1111111111110100;
    assign weights1[42][764] = 16'b0000000000000111;
    assign weights1[42][765] = 16'b1111111111111010;
    assign weights1[42][766] = 16'b1111111111111100;
    assign weights1[42][767] = 16'b0000000000000010;
    assign weights1[42][768] = 16'b0000000000011000;
    assign weights1[42][769] = 16'b1111111111111111;
    assign weights1[42][770] = 16'b1111111111101001;
    assign weights1[42][771] = 16'b1111111111010101;
    assign weights1[42][772] = 16'b1111111111011100;
    assign weights1[42][773] = 16'b1111111111011001;
    assign weights1[42][774] = 16'b1111111111011010;
    assign weights1[42][775] = 16'b1111111111001101;
    assign weights1[42][776] = 16'b1111111111100010;
    assign weights1[42][777] = 16'b1111111111011011;
    assign weights1[42][778] = 16'b1111111111011111;
    assign weights1[42][779] = 16'b1111111111101101;
    assign weights1[42][780] = 16'b1111111111110000;
    assign weights1[42][781] = 16'b1111111111110110;
    assign weights1[42][782] = 16'b0000000000000110;
    assign weights1[42][783] = 16'b0000000000000010;
    assign weights1[43][0] = 16'b0000000000000001;
    assign weights1[43][1] = 16'b0000000000000001;
    assign weights1[43][2] = 16'b0000000000000001;
    assign weights1[43][3] = 16'b0000000000001000;
    assign weights1[43][4] = 16'b0000000000000000;
    assign weights1[43][5] = 16'b1111111111110001;
    assign weights1[43][6] = 16'b1111111111100100;
    assign weights1[43][7] = 16'b1111111111010110;
    assign weights1[43][8] = 16'b1111111111001101;
    assign weights1[43][9] = 16'b1111111111001101;
    assign weights1[43][10] = 16'b1111111111011110;
    assign weights1[43][11] = 16'b0000000000001000;
    assign weights1[43][12] = 16'b0000000000101100;
    assign weights1[43][13] = 16'b0000000000101100;
    assign weights1[43][14] = 16'b0000000000011100;
    assign weights1[43][15] = 16'b0000000000001011;
    assign weights1[43][16] = 16'b1111111111100010;
    assign weights1[43][17] = 16'b1111111110110001;
    assign weights1[43][18] = 16'b1111111110010101;
    assign weights1[43][19] = 16'b1111111110110111;
    assign weights1[43][20] = 16'b1111111111011011;
    assign weights1[43][21] = 16'b1111111111101101;
    assign weights1[43][22] = 16'b0000000000000001;
    assign weights1[43][23] = 16'b0000000000001000;
    assign weights1[43][24] = 16'b0000000000000101;
    assign weights1[43][25] = 16'b0000000000000100;
    assign weights1[43][26] = 16'b0000000000000101;
    assign weights1[43][27] = 16'b0000000000000101;
    assign weights1[43][28] = 16'b0000000000000001;
    assign weights1[43][29] = 16'b0000000000000001;
    assign weights1[43][30] = 16'b0000000000000011;
    assign weights1[43][31] = 16'b0000000000001110;
    assign weights1[43][32] = 16'b0000000000000010;
    assign weights1[43][33] = 16'b1111111111101000;
    assign weights1[43][34] = 16'b1111111111011000;
    assign weights1[43][35] = 16'b1111111111000111;
    assign weights1[43][36] = 16'b1111111110111000;
    assign weights1[43][37] = 16'b1111111111001101;
    assign weights1[43][38] = 16'b1111111111101101;
    assign weights1[43][39] = 16'b0000000000101101;
    assign weights1[43][40] = 16'b0000000000110001;
    assign weights1[43][41] = 16'b0000000000101111;
    assign weights1[43][42] = 16'b0000000000010000;
    assign weights1[43][43] = 16'b1111111111110101;
    assign weights1[43][44] = 16'b1111111110100110;
    assign weights1[43][45] = 16'b1111111110000011;
    assign weights1[43][46] = 16'b1111111110000000;
    assign weights1[43][47] = 16'b1111111110111001;
    assign weights1[43][48] = 16'b1111111111100010;
    assign weights1[43][49] = 16'b0000000000000111;
    assign weights1[43][50] = 16'b0000000000001000;
    assign weights1[43][51] = 16'b0000000000001101;
    assign weights1[43][52] = 16'b0000000000011001;
    assign weights1[43][53] = 16'b0000000000001001;
    assign weights1[43][54] = 16'b0000000000000011;
    assign weights1[43][55] = 16'b0000000000000001;
    assign weights1[43][56] = 16'b0000000000000010;
    assign weights1[43][57] = 16'b0000000000000100;
    assign weights1[43][58] = 16'b0000000000001001;
    assign weights1[43][59] = 16'b0000000000001100;
    assign weights1[43][60] = 16'b0000000000000011;
    assign weights1[43][61] = 16'b1111111111101010;
    assign weights1[43][62] = 16'b1111111111001010;
    assign weights1[43][63] = 16'b1111111110110000;
    assign weights1[43][64] = 16'b1111111110100101;
    assign weights1[43][65] = 16'b1111111111001011;
    assign weights1[43][66] = 16'b1111111111111011;
    assign weights1[43][67] = 16'b0000000000110100;
    assign weights1[43][68] = 16'b0000000000100110;
    assign weights1[43][69] = 16'b0000000000110100;
    assign weights1[43][70] = 16'b0000000000011010;
    assign weights1[43][71] = 16'b1111111111011011;
    assign weights1[43][72] = 16'b1111111101100101;
    assign weights1[43][73] = 16'b1111111101001100;
    assign weights1[43][74] = 16'b1111111110010001;
    assign weights1[43][75] = 16'b1111111111011011;
    assign weights1[43][76] = 16'b1111111111101111;
    assign weights1[43][77] = 16'b0000000000000110;
    assign weights1[43][78] = 16'b0000000000010110;
    assign weights1[43][79] = 16'b0000000000100000;
    assign weights1[43][80] = 16'b0000000000001111;
    assign weights1[43][81] = 16'b0000000000000111;
    assign weights1[43][82] = 16'b0000000000000000;
    assign weights1[43][83] = 16'b1111111111111100;
    assign weights1[43][84] = 16'b0000000000000000;
    assign weights1[43][85] = 16'b0000000000000011;
    assign weights1[43][86] = 16'b0000000000010000;
    assign weights1[43][87] = 16'b0000000000010100;
    assign weights1[43][88] = 16'b0000000000000100;
    assign weights1[43][89] = 16'b1111111111101100;
    assign weights1[43][90] = 16'b1111111111001010;
    assign weights1[43][91] = 16'b1111111110011000;
    assign weights1[43][92] = 16'b1111111110011000;
    assign weights1[43][93] = 16'b1111111111010111;
    assign weights1[43][94] = 16'b0000000000000111;
    assign weights1[43][95] = 16'b0000000000110110;
    assign weights1[43][96] = 16'b0000000000101011;
    assign weights1[43][97] = 16'b0000000000111000;
    assign weights1[43][98] = 16'b0000000000010011;
    assign weights1[43][99] = 16'b1111111110111001;
    assign weights1[43][100] = 16'b1111111100011101;
    assign weights1[43][101] = 16'b1111111101011001;
    assign weights1[43][102] = 16'b1111111111000000;
    assign weights1[43][103] = 16'b0000000000000000;
    assign weights1[43][104] = 16'b0000000000100100;
    assign weights1[43][105] = 16'b0000000000011100;
    assign weights1[43][106] = 16'b0000000000110110;
    assign weights1[43][107] = 16'b0000000000011111;
    assign weights1[43][108] = 16'b0000000000001101;
    assign weights1[43][109] = 16'b1111111111111101;
    assign weights1[43][110] = 16'b1111111111101101;
    assign weights1[43][111] = 16'b1111111111110001;
    assign weights1[43][112] = 16'b0000000000000010;
    assign weights1[43][113] = 16'b0000000000001010;
    assign weights1[43][114] = 16'b0000000000010100;
    assign weights1[43][115] = 16'b0000000000011010;
    assign weights1[43][116] = 16'b0000000000000101;
    assign weights1[43][117] = 16'b1111111111101010;
    assign weights1[43][118] = 16'b1111111110111011;
    assign weights1[43][119] = 16'b1111111110001111;
    assign weights1[43][120] = 16'b1111111110001100;
    assign weights1[43][121] = 16'b1111111111000111;
    assign weights1[43][122] = 16'b0000000000010101;
    assign weights1[43][123] = 16'b0000000000111101;
    assign weights1[43][124] = 16'b0000000000111011;
    assign weights1[43][125] = 16'b0000000000111100;
    assign weights1[43][126] = 16'b1111111111101011;
    assign weights1[43][127] = 16'b1111111101111010;
    assign weights1[43][128] = 16'b1111111100011001;
    assign weights1[43][129] = 16'b1111111101101111;
    assign weights1[43][130] = 16'b1111111111100000;
    assign weights1[43][131] = 16'b0000000000101111;
    assign weights1[43][132] = 16'b0000000000101011;
    assign weights1[43][133] = 16'b0000000000010110;
    assign weights1[43][134] = 16'b0000000000011100;
    assign weights1[43][135] = 16'b0000000000000110;
    assign weights1[43][136] = 16'b0000000000001110;
    assign weights1[43][137] = 16'b1111111111110010;
    assign weights1[43][138] = 16'b1111111111101000;
    assign weights1[43][139] = 16'b1111111111101110;
    assign weights1[43][140] = 16'b0000000000000110;
    assign weights1[43][141] = 16'b0000000000001000;
    assign weights1[43][142] = 16'b0000000000011111;
    assign weights1[43][143] = 16'b0000000000010111;
    assign weights1[43][144] = 16'b0000000000010100;
    assign weights1[43][145] = 16'b1111111111110110;
    assign weights1[43][146] = 16'b1111111111001000;
    assign weights1[43][147] = 16'b1111111110001100;
    assign weights1[43][148] = 16'b1111111101110101;
    assign weights1[43][149] = 16'b0000000000000000;
    assign weights1[43][150] = 16'b0000000000111100;
    assign weights1[43][151] = 16'b0000000000100010;
    assign weights1[43][152] = 16'b0000000001000011;
    assign weights1[43][153] = 16'b0000000000110101;
    assign weights1[43][154] = 16'b1111111111100101;
    assign weights1[43][155] = 16'b1111111101011110;
    assign weights1[43][156] = 16'b1111111100001110;
    assign weights1[43][157] = 16'b1111111111011010;
    assign weights1[43][158] = 16'b0000000001000011;
    assign weights1[43][159] = 16'b0000000000101000;
    assign weights1[43][160] = 16'b0000000000111011;
    assign weights1[43][161] = 16'b0000000000010110;
    assign weights1[43][162] = 16'b0000000000001010;
    assign weights1[43][163] = 16'b0000000000100111;
    assign weights1[43][164] = 16'b0000000000000110;
    assign weights1[43][165] = 16'b1111111111011101;
    assign weights1[43][166] = 16'b1111111111100100;
    assign weights1[43][167] = 16'b1111111111100011;
    assign weights1[43][168] = 16'b0000000000000001;
    assign weights1[43][169] = 16'b0000000000001101;
    assign weights1[43][170] = 16'b0000000000011110;
    assign weights1[43][171] = 16'b0000000000011000;
    assign weights1[43][172] = 16'b0000000000010000;
    assign weights1[43][173] = 16'b0000000000000110;
    assign weights1[43][174] = 16'b1111111111000011;
    assign weights1[43][175] = 16'b1111111101111110;
    assign weights1[43][176] = 16'b1111111101110000;
    assign weights1[43][177] = 16'b0000000000000000;
    assign weights1[43][178] = 16'b0000000000010100;
    assign weights1[43][179] = 16'b0000000000100101;
    assign weights1[43][180] = 16'b0000000000100111;
    assign weights1[43][181] = 16'b0000000000011100;
    assign weights1[43][182] = 16'b1111111111111101;
    assign weights1[43][183] = 16'b1111111100111111;
    assign weights1[43][184] = 16'b1111111101100011;
    assign weights1[43][185] = 16'b0000000000100011;
    assign weights1[43][186] = 16'b0000000000111000;
    assign weights1[43][187] = 16'b0000000000010001;
    assign weights1[43][188] = 16'b0000000000010010;
    assign weights1[43][189] = 16'b0000000000011011;
    assign weights1[43][190] = 16'b0000000000011000;
    assign weights1[43][191] = 16'b1111111111111100;
    assign weights1[43][192] = 16'b1111111111010000;
    assign weights1[43][193] = 16'b1111111111010011;
    assign weights1[43][194] = 16'b1111111111010100;
    assign weights1[43][195] = 16'b1111111111011001;
    assign weights1[43][196] = 16'b0000000000000101;
    assign weights1[43][197] = 16'b0000000000001011;
    assign weights1[43][198] = 16'b0000000000011111;
    assign weights1[43][199] = 16'b0000000000011000;
    assign weights1[43][200] = 16'b0000000000001110;
    assign weights1[43][201] = 16'b0000000000010011;
    assign weights1[43][202] = 16'b1111111111011110;
    assign weights1[43][203] = 16'b1111111110101001;
    assign weights1[43][204] = 16'b1111111110110010;
    assign weights1[43][205] = 16'b1111111111100010;
    assign weights1[43][206] = 16'b0000000000011011;
    assign weights1[43][207] = 16'b0000000000011000;
    assign weights1[43][208] = 16'b0000000000101010;
    assign weights1[43][209] = 16'b0000000000000001;
    assign weights1[43][210] = 16'b1111111111100001;
    assign weights1[43][211] = 16'b1111111101001000;
    assign weights1[43][212] = 16'b1111111111000101;
    assign weights1[43][213] = 16'b0000000000010100;
    assign weights1[43][214] = 16'b0000000000101100;
    assign weights1[43][215] = 16'b0000000000001111;
    assign weights1[43][216] = 16'b0000000000010001;
    assign weights1[43][217] = 16'b0000000000010110;
    assign weights1[43][218] = 16'b0000000000000100;
    assign weights1[43][219] = 16'b1111111111101010;
    assign weights1[43][220] = 16'b1111111110111101;
    assign weights1[43][221] = 16'b1111111111000110;
    assign weights1[43][222] = 16'b1111111111001001;
    assign weights1[43][223] = 16'b1111111111100010;
    assign weights1[43][224] = 16'b0000000000000100;
    assign weights1[43][225] = 16'b0000000000001011;
    assign weights1[43][226] = 16'b0000000000010000;
    assign weights1[43][227] = 16'b0000000000011110;
    assign weights1[43][228] = 16'b0000000000011010;
    assign weights1[43][229] = 16'b0000000000001100;
    assign weights1[43][230] = 16'b1111111111110110;
    assign weights1[43][231] = 16'b1111111111010011;
    assign weights1[43][232] = 16'b1111111110110100;
    assign weights1[43][233] = 16'b1111111111111011;
    assign weights1[43][234] = 16'b0000000000001000;
    assign weights1[43][235] = 16'b0000000000011101;
    assign weights1[43][236] = 16'b0000000000100010;
    assign weights1[43][237] = 16'b0000000000010100;
    assign weights1[43][238] = 16'b1111111111010111;
    assign weights1[43][239] = 16'b1111111110010000;
    assign weights1[43][240] = 16'b1111111111101111;
    assign weights1[43][241] = 16'b0000000000011011;
    assign weights1[43][242] = 16'b0000000000100111;
    assign weights1[43][243] = 16'b0000000000010100;
    assign weights1[43][244] = 16'b0000000000001001;
    assign weights1[43][245] = 16'b0000000000011110;
    assign weights1[43][246] = 16'b1111111111110010;
    assign weights1[43][247] = 16'b1111111111010011;
    assign weights1[43][248] = 16'b1111111110111100;
    assign weights1[43][249] = 16'b1111111111010110;
    assign weights1[43][250] = 16'b1111111111100011;
    assign weights1[43][251] = 16'b1111111111101100;
    assign weights1[43][252] = 16'b0000000000000110;
    assign weights1[43][253] = 16'b0000000000010110;
    assign weights1[43][254] = 16'b0000000000011110;
    assign weights1[43][255] = 16'b0000000000001000;
    assign weights1[43][256] = 16'b0000000000011000;
    assign weights1[43][257] = 16'b0000000000010101;
    assign weights1[43][258] = 16'b1111111111111010;
    assign weights1[43][259] = 16'b1111111111010010;
    assign weights1[43][260] = 16'b1111111111011011;
    assign weights1[43][261] = 16'b1111111111011111;
    assign weights1[43][262] = 16'b1111111111100001;
    assign weights1[43][263] = 16'b0000000000010010;
    assign weights1[43][264] = 16'b0000000000011100;
    assign weights1[43][265] = 16'b0000000000000110;
    assign weights1[43][266] = 16'b1111111111001100;
    assign weights1[43][267] = 16'b1111111111000110;
    assign weights1[43][268] = 16'b1111111111111001;
    assign weights1[43][269] = 16'b0000000000100001;
    assign weights1[43][270] = 16'b0000000000001101;
    assign weights1[43][271] = 16'b0000000000001111;
    assign weights1[43][272] = 16'b1111111111111110;
    assign weights1[43][273] = 16'b1111111111110100;
    assign weights1[43][274] = 16'b1111111111011101;
    assign weights1[43][275] = 16'b1111111110110111;
    assign weights1[43][276] = 16'b1111111111010101;
    assign weights1[43][277] = 16'b1111111111111011;
    assign weights1[43][278] = 16'b1111111111111111;
    assign weights1[43][279] = 16'b0000000000001010;
    assign weights1[43][280] = 16'b0000000000000001;
    assign weights1[43][281] = 16'b0000000000000000;
    assign weights1[43][282] = 16'b0000000000010111;
    assign weights1[43][283] = 16'b0000000000000101;
    assign weights1[43][284] = 16'b0000000000010011;
    assign weights1[43][285] = 16'b0000000000011110;
    assign weights1[43][286] = 16'b1111111111110010;
    assign weights1[43][287] = 16'b1111111111011100;
    assign weights1[43][288] = 16'b1111111111010001;
    assign weights1[43][289] = 16'b0000000000001001;
    assign weights1[43][290] = 16'b1111111111101110;
    assign weights1[43][291] = 16'b0000000000101011;
    assign weights1[43][292] = 16'b0000000000010000;
    assign weights1[43][293] = 16'b1111111111110010;
    assign weights1[43][294] = 16'b1111111111101000;
    assign weights1[43][295] = 16'b1111111111011110;
    assign weights1[43][296] = 16'b0000000000001110;
    assign weights1[43][297] = 16'b0000000000001111;
    assign weights1[43][298] = 16'b0000000000001100;
    assign weights1[43][299] = 16'b0000000000001011;
    assign weights1[43][300] = 16'b1111111111110000;
    assign weights1[43][301] = 16'b1111111111111110;
    assign weights1[43][302] = 16'b1111111111011000;
    assign weights1[43][303] = 16'b1111111111011000;
    assign weights1[43][304] = 16'b1111111111111011;
    assign weights1[43][305] = 16'b0000000000001110;
    assign weights1[43][306] = 16'b0000000000010010;
    assign weights1[43][307] = 16'b0000000000010111;
    assign weights1[43][308] = 16'b0000000000000101;
    assign weights1[43][309] = 16'b1111111111111111;
    assign weights1[43][310] = 16'b0000000000001001;
    assign weights1[43][311] = 16'b1111111111110010;
    assign weights1[43][312] = 16'b1111111111111001;
    assign weights1[43][313] = 16'b0000000000100011;
    assign weights1[43][314] = 16'b0000000000000101;
    assign weights1[43][315] = 16'b1111111111111110;
    assign weights1[43][316] = 16'b1111111111111011;
    assign weights1[43][317] = 16'b1111111111101111;
    assign weights1[43][318] = 16'b1111111111110110;
    assign weights1[43][319] = 16'b0000000000000000;
    assign weights1[43][320] = 16'b0000000000001001;
    assign weights1[43][321] = 16'b1111111111111100;
    assign weights1[43][322] = 16'b1111111111111011;
    assign weights1[43][323] = 16'b1111111111100101;
    assign weights1[43][324] = 16'b0000000000011000;
    assign weights1[43][325] = 16'b0000000000000110;
    assign weights1[43][326] = 16'b1111111111111010;
    assign weights1[43][327] = 16'b0000000000010000;
    assign weights1[43][328] = 16'b1111111111101110;
    assign weights1[43][329] = 16'b1111111111110011;
    assign weights1[43][330] = 16'b1111111111001000;
    assign weights1[43][331] = 16'b0000000000000001;
    assign weights1[43][332] = 16'b0000000000001011;
    assign weights1[43][333] = 16'b0000000000010001;
    assign weights1[43][334] = 16'b0000000000100010;
    assign weights1[43][335] = 16'b0000000000100110;
    assign weights1[43][336] = 16'b1111111111111011;
    assign weights1[43][337] = 16'b1111111111111100;
    assign weights1[43][338] = 16'b0000000000010000;
    assign weights1[43][339] = 16'b0000000000010101;
    assign weights1[43][340] = 16'b0000000000011001;
    assign weights1[43][341] = 16'b1111111111111011;
    assign weights1[43][342] = 16'b0000000000001100;
    assign weights1[43][343] = 16'b0000000000001101;
    assign weights1[43][344] = 16'b1111111111101111;
    assign weights1[43][345] = 16'b1111111111101001;
    assign weights1[43][346] = 16'b1111111111111110;
    assign weights1[43][347] = 16'b0000000000000111;
    assign weights1[43][348] = 16'b0000000000000011;
    assign weights1[43][349] = 16'b0000000000000011;
    assign weights1[43][350] = 16'b1111111111110110;
    assign weights1[43][351] = 16'b0000000000001000;
    assign weights1[43][352] = 16'b0000000000001010;
    assign weights1[43][353] = 16'b0000000000000001;
    assign weights1[43][354] = 16'b1111111111111110;
    assign weights1[43][355] = 16'b1111111111110110;
    assign weights1[43][356] = 16'b1111111111101100;
    assign weights1[43][357] = 16'b1111111111101110;
    assign weights1[43][358] = 16'b1111111111101110;
    assign weights1[43][359] = 16'b0000000000001001;
    assign weights1[43][360] = 16'b0000000000011111;
    assign weights1[43][361] = 16'b0000000000001000;
    assign weights1[43][362] = 16'b0000000000001001;
    assign weights1[43][363] = 16'b0000000000011011;
    assign weights1[43][364] = 16'b1111111111111001;
    assign weights1[43][365] = 16'b0000000000000110;
    assign weights1[43][366] = 16'b0000000000000110;
    assign weights1[43][367] = 16'b1111111111111111;
    assign weights1[43][368] = 16'b0000000000001111;
    assign weights1[43][369] = 16'b1111111111110100;
    assign weights1[43][370] = 16'b1111111111111100;
    assign weights1[43][371] = 16'b0000000000001101;
    assign weights1[43][372] = 16'b0000000000001100;
    assign weights1[43][373] = 16'b0000000000011001;
    assign weights1[43][374] = 16'b1111111111111111;
    assign weights1[43][375] = 16'b0000000000000100;
    assign weights1[43][376] = 16'b0000000000000110;
    assign weights1[43][377] = 16'b0000000000000100;
    assign weights1[43][378] = 16'b1111111111101111;
    assign weights1[43][379] = 16'b1111111111110011;
    assign weights1[43][380] = 16'b1111111111111000;
    assign weights1[43][381] = 16'b0000000000000100;
    assign weights1[43][382] = 16'b1111111111110111;
    assign weights1[43][383] = 16'b1111111111111001;
    assign weights1[43][384] = 16'b0000000000000111;
    assign weights1[43][385] = 16'b1111111111101101;
    assign weights1[43][386] = 16'b0000000000010000;
    assign weights1[43][387] = 16'b0000000000001000;
    assign weights1[43][388] = 16'b0000000000001111;
    assign weights1[43][389] = 16'b0000000000000011;
    assign weights1[43][390] = 16'b0000000000010111;
    assign weights1[43][391] = 16'b0000000000010110;
    assign weights1[43][392] = 16'b1111111111110001;
    assign weights1[43][393] = 16'b1111111111111111;
    assign weights1[43][394] = 16'b1111111111111100;
    assign weights1[43][395] = 16'b1111111111110011;
    assign weights1[43][396] = 16'b1111111111111111;
    assign weights1[43][397] = 16'b0000000000011001;
    assign weights1[43][398] = 16'b0000000000000001;
    assign weights1[43][399] = 16'b0000000000001001;
    assign weights1[43][400] = 16'b0000000000000100;
    assign weights1[43][401] = 16'b1111111111111100;
    assign weights1[43][402] = 16'b1111111111111011;
    assign weights1[43][403] = 16'b0000000000001111;
    assign weights1[43][404] = 16'b0000000000001100;
    assign weights1[43][405] = 16'b1111111111110110;
    assign weights1[43][406] = 16'b0000000000001111;
    assign weights1[43][407] = 16'b0000000000010111;
    assign weights1[43][408] = 16'b0000000000001100;
    assign weights1[43][409] = 16'b1111111111111011;
    assign weights1[43][410] = 16'b1111111111110011;
    assign weights1[43][411] = 16'b0000000000011000;
    assign weights1[43][412] = 16'b0000000000000010;
    assign weights1[43][413] = 16'b0000000000010010;
    assign weights1[43][414] = 16'b0000000000000000;
    assign weights1[43][415] = 16'b0000000000001111;
    assign weights1[43][416] = 16'b0000000000001110;
    assign weights1[43][417] = 16'b0000000000001110;
    assign weights1[43][418] = 16'b0000000000010100;
    assign weights1[43][419] = 16'b0000000000000000;
    assign weights1[43][420] = 16'b0000000000000100;
    assign weights1[43][421] = 16'b1111111111111000;
    assign weights1[43][422] = 16'b0000000000000100;
    assign weights1[43][423] = 16'b0000000000001000;
    assign weights1[43][424] = 16'b0000000000000101;
    assign weights1[43][425] = 16'b0000000000000100;
    assign weights1[43][426] = 16'b1111111111111110;
    assign weights1[43][427] = 16'b0000000000000011;
    assign weights1[43][428] = 16'b0000000000000010;
    assign weights1[43][429] = 16'b0000000000000111;
    assign weights1[43][430] = 16'b0000000000100011;
    assign weights1[43][431] = 16'b1111111111111111;
    assign weights1[43][432] = 16'b0000000000000110;
    assign weights1[43][433] = 16'b0000000000001111;
    assign weights1[43][434] = 16'b0000000000001011;
    assign weights1[43][435] = 16'b0000000000000100;
    assign weights1[43][436] = 16'b1111111111111010;
    assign weights1[43][437] = 16'b0000000000000001;
    assign weights1[43][438] = 16'b1111111111111001;
    assign weights1[43][439] = 16'b0000000000000100;
    assign weights1[43][440] = 16'b0000000000001110;
    assign weights1[43][441] = 16'b0000000000000111;
    assign weights1[43][442] = 16'b0000000000010111;
    assign weights1[43][443] = 16'b0000000000001010;
    assign weights1[43][444] = 16'b1111111111110011;
    assign weights1[43][445] = 16'b1111111111111111;
    assign weights1[43][446] = 16'b1111111111111010;
    assign weights1[43][447] = 16'b1111111111111111;
    assign weights1[43][448] = 16'b1111111111111010;
    assign weights1[43][449] = 16'b1111111111111010;
    assign weights1[43][450] = 16'b0000000000001011;
    assign weights1[43][451] = 16'b0000000000000010;
    assign weights1[43][452] = 16'b0000000000000100;
    assign weights1[43][453] = 16'b0000000000001001;
    assign weights1[43][454] = 16'b0000000000011101;
    assign weights1[43][455] = 16'b1111111111111010;
    assign weights1[43][456] = 16'b0000000000000111;
    assign weights1[43][457] = 16'b1111111111110111;
    assign weights1[43][458] = 16'b1111111111110111;
    assign weights1[43][459] = 16'b1111111111111000;
    assign weights1[43][460] = 16'b1111111111111011;
    assign weights1[43][461] = 16'b1111111111111111;
    assign weights1[43][462] = 16'b0000000000001001;
    assign weights1[43][463] = 16'b0000000000001111;
    assign weights1[43][464] = 16'b1111111111111110;
    assign weights1[43][465] = 16'b1111111111101011;
    assign weights1[43][466] = 16'b1111111111110111;
    assign weights1[43][467] = 16'b0000000000000100;
    assign weights1[43][468] = 16'b1111111111111010;
    assign weights1[43][469] = 16'b0000000000000111;
    assign weights1[43][470] = 16'b0000000000010011;
    assign weights1[43][471] = 16'b0000000000000111;
    assign weights1[43][472] = 16'b0000000000100111;
    assign weights1[43][473] = 16'b1111111111111010;
    assign weights1[43][474] = 16'b1111111111110011;
    assign weights1[43][475] = 16'b1111111111111011;
    assign weights1[43][476] = 16'b1111111111111011;
    assign weights1[43][477] = 16'b0000000000001000;
    assign weights1[43][478] = 16'b0000000000010100;
    assign weights1[43][479] = 16'b1111111111111110;
    assign weights1[43][480] = 16'b0000000000001100;
    assign weights1[43][481] = 16'b1111111111101010;
    assign weights1[43][482] = 16'b1111111111111101;
    assign weights1[43][483] = 16'b0000000000000010;
    assign weights1[43][484] = 16'b1111111111111101;
    assign weights1[43][485] = 16'b1111111111111001;
    assign weights1[43][486] = 16'b0000000000010010;
    assign weights1[43][487] = 16'b1111111111110111;
    assign weights1[43][488] = 16'b0000000000000001;
    assign weights1[43][489] = 16'b1111111111110011;
    assign weights1[43][490] = 16'b0000000000001111;
    assign weights1[43][491] = 16'b1111111111111001;
    assign weights1[43][492] = 16'b0000000000000110;
    assign weights1[43][493] = 16'b1111111111111101;
    assign weights1[43][494] = 16'b0000000000001010;
    assign weights1[43][495] = 16'b1111111111111110;
    assign weights1[43][496] = 16'b0000000000000110;
    assign weights1[43][497] = 16'b0000000000001011;
    assign weights1[43][498] = 16'b0000000000000011;
    assign weights1[43][499] = 16'b0000000000000001;
    assign weights1[43][500] = 16'b0000000000011110;
    assign weights1[43][501] = 16'b1111111111111010;
    assign weights1[43][502] = 16'b1111111111111001;
    assign weights1[43][503] = 16'b1111111111110111;
    assign weights1[43][504] = 16'b1111111111111110;
    assign weights1[43][505] = 16'b0000000000001011;
    assign weights1[43][506] = 16'b0000000000000011;
    assign weights1[43][507] = 16'b0000000000000001;
    assign weights1[43][508] = 16'b1111111111111111;
    assign weights1[43][509] = 16'b1111111111111101;
    assign weights1[43][510] = 16'b0000000000010001;
    assign weights1[43][511] = 16'b1111111111111101;
    assign weights1[43][512] = 16'b0000000000010110;
    assign weights1[43][513] = 16'b0000000000000000;
    assign weights1[43][514] = 16'b0000000000000001;
    assign weights1[43][515] = 16'b0000000000000011;
    assign weights1[43][516] = 16'b0000000000001110;
    assign weights1[43][517] = 16'b0000000000001010;
    assign weights1[43][518] = 16'b0000000000010001;
    assign weights1[43][519] = 16'b1111111111111111;
    assign weights1[43][520] = 16'b1111111111111100;
    assign weights1[43][521] = 16'b0000000000000111;
    assign weights1[43][522] = 16'b0000000000000111;
    assign weights1[43][523] = 16'b1111111111111011;
    assign weights1[43][524] = 16'b1111111111111001;
    assign weights1[43][525] = 16'b0000000000000110;
    assign weights1[43][526] = 16'b0000000000000000;
    assign weights1[43][527] = 16'b0000000000000100;
    assign weights1[43][528] = 16'b0000000000000111;
    assign weights1[43][529] = 16'b0000000000001100;
    assign weights1[43][530] = 16'b0000000000001100;
    assign weights1[43][531] = 16'b1111111111111001;
    assign weights1[43][532] = 16'b0000000000000001;
    assign weights1[43][533] = 16'b1111111111111110;
    assign weights1[43][534] = 16'b0000000000000111;
    assign weights1[43][535] = 16'b0000000000011000;
    assign weights1[43][536] = 16'b0000000000001010;
    assign weights1[43][537] = 16'b1111111111111100;
    assign weights1[43][538] = 16'b1111111111111100;
    assign weights1[43][539] = 16'b1111111111111111;
    assign weights1[43][540] = 16'b0000000000000111;
    assign weights1[43][541] = 16'b1111111111110100;
    assign weights1[43][542] = 16'b0000000000000011;
    assign weights1[43][543] = 16'b0000000000000001;
    assign weights1[43][544] = 16'b1111111111110100;
    assign weights1[43][545] = 16'b1111111111111000;
    assign weights1[43][546] = 16'b0000000000010110;
    assign weights1[43][547] = 16'b0000000000001100;
    assign weights1[43][548] = 16'b0000000000000101;
    assign weights1[43][549] = 16'b1111111111111100;
    assign weights1[43][550] = 16'b1111111111111011;
    assign weights1[43][551] = 16'b1111111111111000;
    assign weights1[43][552] = 16'b0000000000000111;
    assign weights1[43][553] = 16'b0000000000000001;
    assign weights1[43][554] = 16'b0000000000001101;
    assign weights1[43][555] = 16'b0000000000000010;
    assign weights1[43][556] = 16'b1111111111101110;
    assign weights1[43][557] = 16'b1111111111111110;
    assign weights1[43][558] = 16'b0000000000001111;
    assign weights1[43][559] = 16'b1111111111110110;
    assign weights1[43][560] = 16'b0000000000000111;
    assign weights1[43][561] = 16'b0000000000000011;
    assign weights1[43][562] = 16'b0000000000001000;
    assign weights1[43][563] = 16'b1111111111111110;
    assign weights1[43][564] = 16'b1111111111110100;
    assign weights1[43][565] = 16'b1111111111111100;
    assign weights1[43][566] = 16'b1111111111111010;
    assign weights1[43][567] = 16'b0000000000001101;
    assign weights1[43][568] = 16'b1111111111110110;
    assign weights1[43][569] = 16'b0000000000000001;
    assign weights1[43][570] = 16'b1111111111111110;
    assign weights1[43][571] = 16'b1111111111110011;
    assign weights1[43][572] = 16'b1111111111101110;
    assign weights1[43][573] = 16'b0000000000000000;
    assign weights1[43][574] = 16'b0000000000000011;
    assign weights1[43][575] = 16'b0000000000001010;
    assign weights1[43][576] = 16'b1111111111111100;
    assign weights1[43][577] = 16'b1111111111111101;
    assign weights1[43][578] = 16'b0000000000000000;
    assign weights1[43][579] = 16'b0000000000010011;
    assign weights1[43][580] = 16'b1111111111110010;
    assign weights1[43][581] = 16'b1111111111111111;
    assign weights1[43][582] = 16'b1111111111111000;
    assign weights1[43][583] = 16'b0000000000000100;
    assign weights1[43][584] = 16'b1111111111111111;
    assign weights1[43][585] = 16'b1111111111111111;
    assign weights1[43][586] = 16'b0000000000000001;
    assign weights1[43][587] = 16'b1111111111111001;
    assign weights1[43][588] = 16'b0000000000000011;
    assign weights1[43][589] = 16'b1111111111111011;
    assign weights1[43][590] = 16'b1111111111111110;
    assign weights1[43][591] = 16'b0000000000000111;
    assign weights1[43][592] = 16'b0000000000000111;
    assign weights1[43][593] = 16'b0000000000000010;
    assign weights1[43][594] = 16'b0000000000001011;
    assign weights1[43][595] = 16'b1111111111110110;
    assign weights1[43][596] = 16'b0000000000001101;
    assign weights1[43][597] = 16'b1111111111111001;
    assign weights1[43][598] = 16'b1111111111110100;
    assign weights1[43][599] = 16'b0000000000000010;
    assign weights1[43][600] = 16'b1111111111101111;
    assign weights1[43][601] = 16'b0000000000000111;
    assign weights1[43][602] = 16'b1111111111111101;
    assign weights1[43][603] = 16'b0000000000000011;
    assign weights1[43][604] = 16'b0000000000011000;
    assign weights1[43][605] = 16'b0000000000000100;
    assign weights1[43][606] = 16'b1111111111111100;
    assign weights1[43][607] = 16'b1111111111111100;
    assign weights1[43][608] = 16'b0000000000000000;
    assign weights1[43][609] = 16'b0000000000000010;
    assign weights1[43][610] = 16'b1111111111111010;
    assign weights1[43][611] = 16'b1111111111111100;
    assign weights1[43][612] = 16'b1111111111111010;
    assign weights1[43][613] = 16'b1111111111110101;
    assign weights1[43][614] = 16'b1111111111111110;
    assign weights1[43][615] = 16'b1111111111101111;
    assign weights1[43][616] = 16'b0000000000000001;
    assign weights1[43][617] = 16'b0000000000000000;
    assign weights1[43][618] = 16'b0000000000000110;
    assign weights1[43][619] = 16'b1111111111111011;
    assign weights1[43][620] = 16'b1111111111101111;
    assign weights1[43][621] = 16'b0000000000010000;
    assign weights1[43][622] = 16'b0000000000010010;
    assign weights1[43][623] = 16'b1111111111111011;
    assign weights1[43][624] = 16'b1111111111111001;
    assign weights1[43][625] = 16'b1111111111111011;
    assign weights1[43][626] = 16'b0000000000000110;
    assign weights1[43][627] = 16'b1111111111110100;
    assign weights1[43][628] = 16'b1111111111110101;
    assign weights1[43][629] = 16'b1111111111111011;
    assign weights1[43][630] = 16'b1111111111100010;
    assign weights1[43][631] = 16'b1111111111110000;
    assign weights1[43][632] = 16'b1111111111111100;
    assign weights1[43][633] = 16'b1111111111110000;
    assign weights1[43][634] = 16'b0000000000001101;
    assign weights1[43][635] = 16'b1111111111111100;
    assign weights1[43][636] = 16'b0000000000010001;
    assign weights1[43][637] = 16'b0000000000001101;
    assign weights1[43][638] = 16'b1111111111111001;
    assign weights1[43][639] = 16'b1111111111110100;
    assign weights1[43][640] = 16'b1111111111111111;
    assign weights1[43][641] = 16'b1111111111101011;
    assign weights1[43][642] = 16'b1111111111110101;
    assign weights1[43][643] = 16'b1111111111110101;
    assign weights1[43][644] = 16'b0000000000000010;
    assign weights1[43][645] = 16'b0000000000000101;
    assign weights1[43][646] = 16'b0000000000000100;
    assign weights1[43][647] = 16'b1111111111111001;
    assign weights1[43][648] = 16'b1111111111101101;
    assign weights1[43][649] = 16'b1111111111110111;
    assign weights1[43][650] = 16'b1111111111110111;
    assign weights1[43][651] = 16'b1111111111111100;
    assign weights1[43][652] = 16'b1111111111111100;
    assign weights1[43][653] = 16'b0000000000001001;
    assign weights1[43][654] = 16'b1111111111101000;
    assign weights1[43][655] = 16'b0000000000000000;
    assign weights1[43][656] = 16'b1111111111101111;
    assign weights1[43][657] = 16'b1111111111111001;
    assign weights1[43][658] = 16'b0000000000001000;
    assign weights1[43][659] = 16'b1111111111100010;
    assign weights1[43][660] = 16'b0000000000010110;
    assign weights1[43][661] = 16'b0000000000001000;
    assign weights1[43][662] = 16'b1111111111111001;
    assign weights1[43][663] = 16'b1111111111111010;
    assign weights1[43][664] = 16'b0000000000001011;
    assign weights1[43][665] = 16'b1111111111101000;
    assign weights1[43][666] = 16'b0000000000001000;
    assign weights1[43][667] = 16'b0000000000001011;
    assign weights1[43][668] = 16'b1111111111101110;
    assign weights1[43][669] = 16'b1111111111110110;
    assign weights1[43][670] = 16'b1111111111111000;
    assign weights1[43][671] = 16'b1111111111110010;
    assign weights1[43][672] = 16'b0000000000000001;
    assign weights1[43][673] = 16'b0000000000000000;
    assign weights1[43][674] = 16'b1111111111111001;
    assign weights1[43][675] = 16'b1111111111101101;
    assign weights1[43][676] = 16'b1111111111111010;
    assign weights1[43][677] = 16'b0000000000000101;
    assign weights1[43][678] = 16'b0000000000000001;
    assign weights1[43][679] = 16'b0000000000000011;
    assign weights1[43][680] = 16'b1111111111110000;
    assign weights1[43][681] = 16'b0000000000001011;
    assign weights1[43][682] = 16'b0000000000000111;
    assign weights1[43][683] = 16'b1111111111110101;
    assign weights1[43][684] = 16'b1111111111111000;
    assign weights1[43][685] = 16'b0000000000010101;
    assign weights1[43][686] = 16'b0000000000010101;
    assign weights1[43][687] = 16'b1111111111101110;
    assign weights1[43][688] = 16'b1111111111101010;
    assign weights1[43][689] = 16'b1111111111100101;
    assign weights1[43][690] = 16'b1111111111101101;
    assign weights1[43][691] = 16'b0000000000000011;
    assign weights1[43][692] = 16'b1111111111100111;
    assign weights1[43][693] = 16'b1111111111101111;
    assign weights1[43][694] = 16'b1111111111111011;
    assign weights1[43][695] = 16'b0000000000000100;
    assign weights1[43][696] = 16'b1111111111110110;
    assign weights1[43][697] = 16'b1111111111111100;
    assign weights1[43][698] = 16'b1111111111110111;
    assign weights1[43][699] = 16'b1111111111111010;
    assign weights1[43][700] = 16'b1111111111111111;
    assign weights1[43][701] = 16'b1111111111111010;
    assign weights1[43][702] = 16'b1111111111111111;
    assign weights1[43][703] = 16'b1111111111111100;
    assign weights1[43][704] = 16'b0000000000000110;
    assign weights1[43][705] = 16'b1111111111111001;
    assign weights1[43][706] = 16'b1111111111111101;
    assign weights1[43][707] = 16'b1111111111111110;
    assign weights1[43][708] = 16'b0000000000000111;
    assign weights1[43][709] = 16'b1111111111111111;
    assign weights1[43][710] = 16'b1111111111111111;
    assign weights1[43][711] = 16'b1111111111111000;
    assign weights1[43][712] = 16'b1111111111100110;
    assign weights1[43][713] = 16'b1111111111101110;
    assign weights1[43][714] = 16'b1111111111111010;
    assign weights1[43][715] = 16'b1111111111110101;
    assign weights1[43][716] = 16'b1111111111110011;
    assign weights1[43][717] = 16'b1111111111111110;
    assign weights1[43][718] = 16'b1111111111101001;
    assign weights1[43][719] = 16'b1111111111101010;
    assign weights1[43][720] = 16'b1111111111101100;
    assign weights1[43][721] = 16'b1111111111101111;
    assign weights1[43][722] = 16'b1111111111100000;
    assign weights1[43][723] = 16'b1111111111110001;
    assign weights1[43][724] = 16'b1111111111110010;
    assign weights1[43][725] = 16'b1111111111110100;
    assign weights1[43][726] = 16'b1111111111111111;
    assign weights1[43][727] = 16'b0000000000000000;
    assign weights1[43][728] = 16'b0000000000000000;
    assign weights1[43][729] = 16'b1111111111111110;
    assign weights1[43][730] = 16'b0000000000000010;
    assign weights1[43][731] = 16'b1111111111111111;
    assign weights1[43][732] = 16'b1111111111111011;
    assign weights1[43][733] = 16'b1111111111110011;
    assign weights1[43][734] = 16'b1111111111110001;
    assign weights1[43][735] = 16'b1111111111111010;
    assign weights1[43][736] = 16'b0000000000000000;
    assign weights1[43][737] = 16'b0000000000000100;
    assign weights1[43][738] = 16'b1111111111111010;
    assign weights1[43][739] = 16'b1111111111110110;
    assign weights1[43][740] = 16'b0000000000000100;
    assign weights1[43][741] = 16'b1111111111100100;
    assign weights1[43][742] = 16'b1111111111111001;
    assign weights1[43][743] = 16'b1111111111100110;
    assign weights1[43][744] = 16'b1111111111111001;
    assign weights1[43][745] = 16'b1111111111101110;
    assign weights1[43][746] = 16'b1111111111111111;
    assign weights1[43][747] = 16'b1111111111101101;
    assign weights1[43][748] = 16'b0000000000000000;
    assign weights1[43][749] = 16'b1111111111111000;
    assign weights1[43][750] = 16'b1111111111101101;
    assign weights1[43][751] = 16'b1111111111111001;
    assign weights1[43][752] = 16'b1111111111101110;
    assign weights1[43][753] = 16'b1111111111111011;
    assign weights1[43][754] = 16'b1111111111111111;
    assign weights1[43][755] = 16'b0000000000000001;
    assign weights1[43][756] = 16'b0000000000000000;
    assign weights1[43][757] = 16'b0000000000000001;
    assign weights1[43][758] = 16'b0000000000000100;
    assign weights1[43][759] = 16'b0000000000001000;
    assign weights1[43][760] = 16'b0000000000000100;
    assign weights1[43][761] = 16'b1111111111110001;
    assign weights1[43][762] = 16'b1111111111100110;
    assign weights1[43][763] = 16'b1111111111110001;
    assign weights1[43][764] = 16'b1111111111111000;
    assign weights1[43][765] = 16'b0000000000000010;
    assign weights1[43][766] = 16'b1111111111111101;
    assign weights1[43][767] = 16'b1111111111110000;
    assign weights1[43][768] = 16'b0000000000000011;
    assign weights1[43][769] = 16'b1111111111111001;
    assign weights1[43][770] = 16'b1111111111100011;
    assign weights1[43][771] = 16'b1111111111110001;
    assign weights1[43][772] = 16'b1111111111101111;
    assign weights1[43][773] = 16'b1111111111101111;
    assign weights1[43][774] = 16'b1111111111101010;
    assign weights1[43][775] = 16'b1111111111100100;
    assign weights1[43][776] = 16'b1111111111111010;
    assign weights1[43][777] = 16'b1111111111110000;
    assign weights1[43][778] = 16'b1111111111110101;
    assign weights1[43][779] = 16'b1111111111110111;
    assign weights1[43][780] = 16'b1111111111110011;
    assign weights1[43][781] = 16'b1111111111111100;
    assign weights1[43][782] = 16'b0000000000000001;
    assign weights1[43][783] = 16'b0000000000000001;
    assign weights1[44][0] = 16'b1111111111111111;
    assign weights1[44][1] = 16'b1111111111111111;
    assign weights1[44][2] = 16'b1111111111111101;
    assign weights1[44][3] = 16'b1111111111111101;
    assign weights1[44][4] = 16'b1111111111111011;
    assign weights1[44][5] = 16'b1111111111110111;
    assign weights1[44][6] = 16'b1111111111111000;
    assign weights1[44][7] = 16'b1111111111111001;
    assign weights1[44][8] = 16'b1111111111101111;
    assign weights1[44][9] = 16'b1111111111101110;
    assign weights1[44][10] = 16'b1111111111100111;
    assign weights1[44][11] = 16'b1111111111010011;
    assign weights1[44][12] = 16'b1111111111001010;
    assign weights1[44][13] = 16'b1111111110111000;
    assign weights1[44][14] = 16'b1111111110110000;
    assign weights1[44][15] = 16'b1111111110101001;
    assign weights1[44][16] = 16'b1111111110010011;
    assign weights1[44][17] = 16'b1111111110100110;
    assign weights1[44][18] = 16'b1111111111000000;
    assign weights1[44][19] = 16'b1111111111001110;
    assign weights1[44][20] = 16'b1111111111011001;
    assign weights1[44][21] = 16'b1111111111100011;
    assign weights1[44][22] = 16'b1111111111110000;
    assign weights1[44][23] = 16'b1111111111111100;
    assign weights1[44][24] = 16'b1111111111111111;
    assign weights1[44][25] = 16'b0000000000000000;
    assign weights1[44][26] = 16'b0000000000000000;
    assign weights1[44][27] = 16'b0000000000000000;
    assign weights1[44][28] = 16'b1111111111111111;
    assign weights1[44][29] = 16'b0000000000000000;
    assign weights1[44][30] = 16'b1111111111111010;
    assign weights1[44][31] = 16'b1111111111111110;
    assign weights1[44][32] = 16'b1111111111111010;
    assign weights1[44][33] = 16'b1111111111110011;
    assign weights1[44][34] = 16'b1111111111111100;
    assign weights1[44][35] = 16'b1111111111111011;
    assign weights1[44][36] = 16'b0000000000010011;
    assign weights1[44][37] = 16'b1111111111111110;
    assign weights1[44][38] = 16'b0000000000000011;
    assign weights1[44][39] = 16'b0000000000000110;
    assign weights1[44][40] = 16'b1111111111110110;
    assign weights1[44][41] = 16'b1111111111100000;
    assign weights1[44][42] = 16'b1111111111011010;
    assign weights1[44][43] = 16'b1111111111001000;
    assign weights1[44][44] = 16'b1111111110101010;
    assign weights1[44][45] = 16'b1111111110010111;
    assign weights1[44][46] = 16'b1111111110101000;
    assign weights1[44][47] = 16'b1111111110111000;
    assign weights1[44][48] = 16'b1111111111001001;
    assign weights1[44][49] = 16'b1111111111011011;
    assign weights1[44][50] = 16'b1111111111101100;
    assign weights1[44][51] = 16'b1111111111110100;
    assign weights1[44][52] = 16'b1111111111111100;
    assign weights1[44][53] = 16'b1111111111111100;
    assign weights1[44][54] = 16'b1111111111111110;
    assign weights1[44][55] = 16'b1111111111111111;
    assign weights1[44][56] = 16'b1111111111111110;
    assign weights1[44][57] = 16'b1111111111111011;
    assign weights1[44][58] = 16'b1111111111111101;
    assign weights1[44][59] = 16'b0000000000000001;
    assign weights1[44][60] = 16'b1111111111111000;
    assign weights1[44][61] = 16'b1111111111111000;
    assign weights1[44][62] = 16'b1111111111111111;
    assign weights1[44][63] = 16'b0000000000000001;
    assign weights1[44][64] = 16'b0000000000010100;
    assign weights1[44][65] = 16'b0000000000100000;
    assign weights1[44][66] = 16'b0000000000100100;
    assign weights1[44][67] = 16'b0000000000010000;
    assign weights1[44][68] = 16'b0000000000110001;
    assign weights1[44][69] = 16'b0000000000101001;
    assign weights1[44][70] = 16'b1111111111111100;
    assign weights1[44][71] = 16'b1111111111101100;
    assign weights1[44][72] = 16'b1111111111100011;
    assign weights1[44][73] = 16'b1111111110111100;
    assign weights1[44][74] = 16'b1111111110010100;
    assign weights1[44][75] = 16'b1111111110011010;
    assign weights1[44][76] = 16'b1111111110101001;
    assign weights1[44][77] = 16'b1111111111000101;
    assign weights1[44][78] = 16'b1111111111010111;
    assign weights1[44][79] = 16'b1111111111101101;
    assign weights1[44][80] = 16'b1111111111110001;
    assign weights1[44][81] = 16'b1111111111110111;
    assign weights1[44][82] = 16'b1111111111111010;
    assign weights1[44][83] = 16'b1111111111111111;
    assign weights1[44][84] = 16'b1111111111111110;
    assign weights1[44][85] = 16'b1111111111111111;
    assign weights1[44][86] = 16'b0000000000000010;
    assign weights1[44][87] = 16'b1111111111111100;
    assign weights1[44][88] = 16'b0000000000000101;
    assign weights1[44][89] = 16'b1111111111110011;
    assign weights1[44][90] = 16'b0000000000000010;
    assign weights1[44][91] = 16'b1111111111111111;
    assign weights1[44][92] = 16'b0000000000010000;
    assign weights1[44][93] = 16'b0000000000001011;
    assign weights1[44][94] = 16'b0000000000010011;
    assign weights1[44][95] = 16'b0000000000110011;
    assign weights1[44][96] = 16'b0000000000100110;
    assign weights1[44][97] = 16'b0000000000101110;
    assign weights1[44][98] = 16'b0000000000101001;
    assign weights1[44][99] = 16'b0000000000010001;
    assign weights1[44][100] = 16'b1111111111110100;
    assign weights1[44][101] = 16'b1111111111111100;
    assign weights1[44][102] = 16'b1111111111001011;
    assign weights1[44][103] = 16'b1111111110011010;
    assign weights1[44][104] = 16'b1111111110000110;
    assign weights1[44][105] = 16'b1111111110001111;
    assign weights1[44][106] = 16'b1111111110111100;
    assign weights1[44][107] = 16'b1111111111011100;
    assign weights1[44][108] = 16'b1111111111101010;
    assign weights1[44][109] = 16'b1111111111101110;
    assign weights1[44][110] = 16'b1111111111111000;
    assign weights1[44][111] = 16'b1111111111111110;
    assign weights1[44][112] = 16'b1111111111111110;
    assign weights1[44][113] = 16'b0000000000000101;
    assign weights1[44][114] = 16'b0000000000000010;
    assign weights1[44][115] = 16'b1111111111111001;
    assign weights1[44][116] = 16'b0000000000000011;
    assign weights1[44][117] = 16'b0000000000000000;
    assign weights1[44][118] = 16'b0000000000010001;
    assign weights1[44][119] = 16'b0000000000010000;
    assign weights1[44][120] = 16'b0000000000000001;
    assign weights1[44][121] = 16'b0000000000101010;
    assign weights1[44][122] = 16'b0000000000011010;
    assign weights1[44][123] = 16'b0000000000110111;
    assign weights1[44][124] = 16'b0000000001000110;
    assign weights1[44][125] = 16'b0000000001000100;
    assign weights1[44][126] = 16'b0000000000101001;
    assign weights1[44][127] = 16'b0000000000011001;
    assign weights1[44][128] = 16'b0000000000001111;
    assign weights1[44][129] = 16'b1111111111111110;
    assign weights1[44][130] = 16'b1111111111101010;
    assign weights1[44][131] = 16'b1111111111011110;
    assign weights1[44][132] = 16'b1111111110110011;
    assign weights1[44][133] = 16'b1111111101110100;
    assign weights1[44][134] = 16'b1111111110011101;
    assign weights1[44][135] = 16'b1111111111001101;
    assign weights1[44][136] = 16'b1111111111100001;
    assign weights1[44][137] = 16'b1111111111101000;
    assign weights1[44][138] = 16'b1111111111111010;
    assign weights1[44][139] = 16'b1111111111111110;
    assign weights1[44][140] = 16'b1111111111111010;
    assign weights1[44][141] = 16'b1111111111111011;
    assign weights1[44][142] = 16'b1111111111111010;
    assign weights1[44][143] = 16'b1111111111110010;
    assign weights1[44][144] = 16'b1111111111111010;
    assign weights1[44][145] = 16'b0000000000000100;
    assign weights1[44][146] = 16'b0000000000001010;
    assign weights1[44][147] = 16'b0000000000001110;
    assign weights1[44][148] = 16'b0000000000010011;
    assign weights1[44][149] = 16'b0000000000001100;
    assign weights1[44][150] = 16'b0000000000011001;
    assign weights1[44][151] = 16'b0000000000011100;
    assign weights1[44][152] = 16'b0000000000100011;
    assign weights1[44][153] = 16'b0000000000110000;
    assign weights1[44][154] = 16'b1111111111111110;
    assign weights1[44][155] = 16'b0000000000101000;
    assign weights1[44][156] = 16'b0000000000001001;
    assign weights1[44][157] = 16'b1111111111110111;
    assign weights1[44][158] = 16'b0000000000000001;
    assign weights1[44][159] = 16'b1111111111111111;
    assign weights1[44][160] = 16'b1111111111100100;
    assign weights1[44][161] = 16'b1111111110101100;
    assign weights1[44][162] = 16'b1111111110010110;
    assign weights1[44][163] = 16'b1111111111000001;
    assign weights1[44][164] = 16'b1111111111010100;
    assign weights1[44][165] = 16'b1111111111101000;
    assign weights1[44][166] = 16'b1111111111110111;
    assign weights1[44][167] = 16'b1111111111111011;
    assign weights1[44][168] = 16'b1111111111110100;
    assign weights1[44][169] = 16'b1111111111110100;
    assign weights1[44][170] = 16'b1111111111110000;
    assign weights1[44][171] = 16'b1111111111101011;
    assign weights1[44][172] = 16'b1111111111011001;
    assign weights1[44][173] = 16'b1111111111110110;
    assign weights1[44][174] = 16'b1111111111111100;
    assign weights1[44][175] = 16'b1111111111101001;
    assign weights1[44][176] = 16'b1111111111111111;
    assign weights1[44][177] = 16'b1111111111110111;
    assign weights1[44][178] = 16'b1111111111110010;
    assign weights1[44][179] = 16'b0000000000000011;
    assign weights1[44][180] = 16'b1111111111111001;
    assign weights1[44][181] = 16'b0000000000101010;
    assign weights1[44][182] = 16'b0000000001001000;
    assign weights1[44][183] = 16'b0000000000010110;
    assign weights1[44][184] = 16'b0000000000100101;
    assign weights1[44][185] = 16'b0000000000010111;
    assign weights1[44][186] = 16'b0000000000010111;
    assign weights1[44][187] = 16'b1111111111110110;
    assign weights1[44][188] = 16'b1111111111100111;
    assign weights1[44][189] = 16'b1111111110111010;
    assign weights1[44][190] = 16'b1111111110010110;
    assign weights1[44][191] = 16'b1111111110010010;
    assign weights1[44][192] = 16'b1111111110111110;
    assign weights1[44][193] = 16'b1111111111011101;
    assign weights1[44][194] = 16'b1111111111110001;
    assign weights1[44][195] = 16'b1111111111111100;
    assign weights1[44][196] = 16'b1111111111110101;
    assign weights1[44][197] = 16'b1111111111110101;
    assign weights1[44][198] = 16'b1111111111100101;
    assign weights1[44][199] = 16'b1111111111010001;
    assign weights1[44][200] = 16'b1111111111010010;
    assign weights1[44][201] = 16'b1111111111001100;
    assign weights1[44][202] = 16'b1111111111110010;
    assign weights1[44][203] = 16'b1111111111010011;
    assign weights1[44][204] = 16'b1111111111011110;
    assign weights1[44][205] = 16'b1111111110111011;
    assign weights1[44][206] = 16'b1111111111101000;
    assign weights1[44][207] = 16'b1111111111110000;
    assign weights1[44][208] = 16'b1111111111110110;
    assign weights1[44][209] = 16'b0000000000110011;
    assign weights1[44][210] = 16'b0000000001011101;
    assign weights1[44][211] = 16'b0000000000110011;
    assign weights1[44][212] = 16'b0000000000100100;
    assign weights1[44][213] = 16'b0000000000100000;
    assign weights1[44][214] = 16'b0000000000000110;
    assign weights1[44][215] = 16'b0000000000000010;
    assign weights1[44][216] = 16'b1111111111111011;
    assign weights1[44][217] = 16'b1111111111110110;
    assign weights1[44][218] = 16'b1111111111001011;
    assign weights1[44][219] = 16'b1111111110001011;
    assign weights1[44][220] = 16'b1111111110110111;
    assign weights1[44][221] = 16'b1111111111011110;
    assign weights1[44][222] = 16'b1111111111101011;
    assign weights1[44][223] = 16'b1111111111111011;
    assign weights1[44][224] = 16'b1111111111111010;
    assign weights1[44][225] = 16'b1111111111101110;
    assign weights1[44][226] = 16'b1111111111011110;
    assign weights1[44][227] = 16'b1111111111100100;
    assign weights1[44][228] = 16'b1111111111001010;
    assign weights1[44][229] = 16'b1111111111001111;
    assign weights1[44][230] = 16'b1111111111011001;
    assign weights1[44][231] = 16'b1111111111000101;
    assign weights1[44][232] = 16'b1111111111001101;
    assign weights1[44][233] = 16'b1111111111110000;
    assign weights1[44][234] = 16'b1111111111110100;
    assign weights1[44][235] = 16'b1111111111100101;
    assign weights1[44][236] = 16'b1111111111101001;
    assign weights1[44][237] = 16'b1111111111111101;
    assign weights1[44][238] = 16'b0000000000101001;
    assign weights1[44][239] = 16'b0000000001010100;
    assign weights1[44][240] = 16'b0000000001001000;
    assign weights1[44][241] = 16'b0000000000100010;
    assign weights1[44][242] = 16'b0000000000100000;
    assign weights1[44][243] = 16'b0000000000001111;
    assign weights1[44][244] = 16'b0000000000000001;
    assign weights1[44][245] = 16'b1111111111111010;
    assign weights1[44][246] = 16'b1111111111011000;
    assign weights1[44][247] = 16'b1111111110010110;
    assign weights1[44][248] = 16'b1111111110101010;
    assign weights1[44][249] = 16'b1111111111001100;
    assign weights1[44][250] = 16'b1111111111101100;
    assign weights1[44][251] = 16'b1111111111110100;
    assign weights1[44][252] = 16'b1111111111111011;
    assign weights1[44][253] = 16'b1111111111101100;
    assign weights1[44][254] = 16'b1111111111010111;
    assign weights1[44][255] = 16'b1111111111100000;
    assign weights1[44][256] = 16'b1111111111011001;
    assign weights1[44][257] = 16'b1111111111001001;
    assign weights1[44][258] = 16'b1111111111100100;
    assign weights1[44][259] = 16'b1111111111101011;
    assign weights1[44][260] = 16'b1111111111110101;
    assign weights1[44][261] = 16'b1111111111101011;
    assign weights1[44][262] = 16'b1111111111111001;
    assign weights1[44][263] = 16'b1111111111100101;
    assign weights1[44][264] = 16'b1111111111011011;
    assign weights1[44][265] = 16'b1111111111101111;
    assign weights1[44][266] = 16'b0000000000001011;
    assign weights1[44][267] = 16'b0000000000110001;
    assign weights1[44][268] = 16'b0000000001000101;
    assign weights1[44][269] = 16'b0000000000100000;
    assign weights1[44][270] = 16'b0000000000100010;
    assign weights1[44][271] = 16'b0000000000010001;
    assign weights1[44][272] = 16'b0000000000000101;
    assign weights1[44][273] = 16'b0000000000000101;
    assign weights1[44][274] = 16'b1111111111001111;
    assign weights1[44][275] = 16'b1111111110101110;
    assign weights1[44][276] = 16'b1111111110111001;
    assign weights1[44][277] = 16'b1111111111011010;
    assign weights1[44][278] = 16'b1111111111101110;
    assign weights1[44][279] = 16'b1111111111110101;
    assign weights1[44][280] = 16'b1111111111111101;
    assign weights1[44][281] = 16'b1111111111101110;
    assign weights1[44][282] = 16'b1111111111100000;
    assign weights1[44][283] = 16'b1111111111101011;
    assign weights1[44][284] = 16'b1111111111110100;
    assign weights1[44][285] = 16'b0000000000000000;
    assign weights1[44][286] = 16'b0000000000001100;
    assign weights1[44][287] = 16'b1111111111110010;
    assign weights1[44][288] = 16'b0000000000000100;
    assign weights1[44][289] = 16'b1111111111101100;
    assign weights1[44][290] = 16'b1111111111110100;
    assign weights1[44][291] = 16'b1111111111110101;
    assign weights1[44][292] = 16'b1111111111110110;
    assign weights1[44][293] = 16'b1111111111001111;
    assign weights1[44][294] = 16'b1111111111110101;
    assign weights1[44][295] = 16'b0000000000010100;
    assign weights1[44][296] = 16'b0000000000110111;
    assign weights1[44][297] = 16'b0000000000110110;
    assign weights1[44][298] = 16'b0000000000100010;
    assign weights1[44][299] = 16'b0000000000101000;
    assign weights1[44][300] = 16'b1111111111110011;
    assign weights1[44][301] = 16'b0000000000000011;
    assign weights1[44][302] = 16'b1111111111110100;
    assign weights1[44][303] = 16'b1111111110100100;
    assign weights1[44][304] = 16'b1111111110110110;
    assign weights1[44][305] = 16'b1111111111011010;
    assign weights1[44][306] = 16'b1111111111100101;
    assign weights1[44][307] = 16'b1111111111110110;
    assign weights1[44][308] = 16'b1111111111111100;
    assign weights1[44][309] = 16'b1111111111110111;
    assign weights1[44][310] = 16'b1111111111101101;
    assign weights1[44][311] = 16'b0000000000000100;
    assign weights1[44][312] = 16'b1111111111111110;
    assign weights1[44][313] = 16'b0000000000011010;
    assign weights1[44][314] = 16'b0000000000010000;
    assign weights1[44][315] = 16'b0000000000010111;
    assign weights1[44][316] = 16'b1111111111111111;
    assign weights1[44][317] = 16'b0000000000001010;
    assign weights1[44][318] = 16'b1111111111110111;
    assign weights1[44][319] = 16'b1111111111110010;
    assign weights1[44][320] = 16'b1111111111001011;
    assign weights1[44][321] = 16'b1111111111101111;
    assign weights1[44][322] = 16'b1111111111100111;
    assign weights1[44][323] = 16'b0000000000011100;
    assign weights1[44][324] = 16'b0000000000000111;
    assign weights1[44][325] = 16'b0000000000101111;
    assign weights1[44][326] = 16'b0000000000100010;
    assign weights1[44][327] = 16'b0000000000101100;
    assign weights1[44][328] = 16'b0000000000101100;
    assign weights1[44][329] = 16'b0000000000000111;
    assign weights1[44][330] = 16'b1111111111011101;
    assign weights1[44][331] = 16'b1111111111001001;
    assign weights1[44][332] = 16'b1111111110101011;
    assign weights1[44][333] = 16'b1111111111100010;
    assign weights1[44][334] = 16'b1111111111110101;
    assign weights1[44][335] = 16'b1111111111111000;
    assign weights1[44][336] = 16'b0000000000001001;
    assign weights1[44][337] = 16'b0000000000000000;
    assign weights1[44][338] = 16'b1111111111111010;
    assign weights1[44][339] = 16'b0000000000000110;
    assign weights1[44][340] = 16'b0000000000000111;
    assign weights1[44][341] = 16'b1111111111110111;
    assign weights1[44][342] = 16'b0000000000001100;
    assign weights1[44][343] = 16'b1111111111111000;
    assign weights1[44][344] = 16'b1111111111111011;
    assign weights1[44][345] = 16'b1111111111111101;
    assign weights1[44][346] = 16'b1111111111101000;
    assign weights1[44][347] = 16'b1111111111011101;
    assign weights1[44][348] = 16'b1111111111010111;
    assign weights1[44][349] = 16'b1111111111011111;
    assign weights1[44][350] = 16'b1111111111110001;
    assign weights1[44][351] = 16'b0000000000000111;
    assign weights1[44][352] = 16'b1111111111111111;
    assign weights1[44][353] = 16'b0000000000011110;
    assign weights1[44][354] = 16'b0000000000001101;
    assign weights1[44][355] = 16'b0000000000010011;
    assign weights1[44][356] = 16'b0000000000011110;
    assign weights1[44][357] = 16'b0000000000010010;
    assign weights1[44][358] = 16'b1111111111100110;
    assign weights1[44][359] = 16'b1111111110111110;
    assign weights1[44][360] = 16'b1111111111010111;
    assign weights1[44][361] = 16'b1111111111101101;
    assign weights1[44][362] = 16'b1111111111111110;
    assign weights1[44][363] = 16'b0000000000000100;
    assign weights1[44][364] = 16'b0000000000010101;
    assign weights1[44][365] = 16'b0000000000000110;
    assign weights1[44][366] = 16'b1111111111111011;
    assign weights1[44][367] = 16'b0000000000000000;
    assign weights1[44][368] = 16'b1111111111110111;
    assign weights1[44][369] = 16'b1111111111110001;
    assign weights1[44][370] = 16'b0000000000000011;
    assign weights1[44][371] = 16'b1111111111101001;
    assign weights1[44][372] = 16'b1111111111111001;
    assign weights1[44][373] = 16'b1111111111110001;
    assign weights1[44][374] = 16'b1111111111100011;
    assign weights1[44][375] = 16'b1111111111110001;
    assign weights1[44][376] = 16'b1111111111101111;
    assign weights1[44][377] = 16'b1111111111010011;
    assign weights1[44][378] = 16'b1111111111101011;
    assign weights1[44][379] = 16'b1111111111110111;
    assign weights1[44][380] = 16'b0000000000010110;
    assign weights1[44][381] = 16'b0000000000011000;
    assign weights1[44][382] = 16'b0000000000001111;
    assign weights1[44][383] = 16'b0000000000010111;
    assign weights1[44][384] = 16'b0000000000000010;
    assign weights1[44][385] = 16'b1111111111111011;
    assign weights1[44][386] = 16'b1111111111111010;
    assign weights1[44][387] = 16'b1111111111011110;
    assign weights1[44][388] = 16'b1111111111100000;
    assign weights1[44][389] = 16'b1111111111110001;
    assign weights1[44][390] = 16'b1111111111111000;
    assign weights1[44][391] = 16'b1111111111111100;
    assign weights1[44][392] = 16'b0000000000010000;
    assign weights1[44][393] = 16'b0000000000001111;
    assign weights1[44][394] = 16'b1111111111111111;
    assign weights1[44][395] = 16'b0000000000001010;
    assign weights1[44][396] = 16'b0000000000001000;
    assign weights1[44][397] = 16'b1111111111111011;
    assign weights1[44][398] = 16'b1111111111011110;
    assign weights1[44][399] = 16'b1111111111111010;
    assign weights1[44][400] = 16'b1111111111111000;
    assign weights1[44][401] = 16'b1111111111110111;
    assign weights1[44][402] = 16'b1111111111101100;
    assign weights1[44][403] = 16'b1111111111111101;
    assign weights1[44][404] = 16'b1111111111110001;
    assign weights1[44][405] = 16'b1111111111110100;
    assign weights1[44][406] = 16'b1111111111101111;
    assign weights1[44][407] = 16'b0000000000000001;
    assign weights1[44][408] = 16'b0000000000000010;
    assign weights1[44][409] = 16'b0000000000011111;
    assign weights1[44][410] = 16'b0000000000010100;
    assign weights1[44][411] = 16'b0000000000001010;
    assign weights1[44][412] = 16'b1111111111111001;
    assign weights1[44][413] = 16'b1111111111110010;
    assign weights1[44][414] = 16'b1111111111110111;
    assign weights1[44][415] = 16'b1111111111110010;
    assign weights1[44][416] = 16'b1111111111111101;
    assign weights1[44][417] = 16'b1111111111101011;
    assign weights1[44][418] = 16'b0000000000001010;
    assign weights1[44][419] = 16'b1111111111111101;
    assign weights1[44][420] = 16'b0000000000001011;
    assign weights1[44][421] = 16'b0000000000001111;
    assign weights1[44][422] = 16'b0000000000001010;
    assign weights1[44][423] = 16'b1111111111111101;
    assign weights1[44][424] = 16'b1111111111110110;
    assign weights1[44][425] = 16'b1111111111111111;
    assign weights1[44][426] = 16'b1111111111111011;
    assign weights1[44][427] = 16'b1111111111111001;
    assign weights1[44][428] = 16'b1111111111111100;
    assign weights1[44][429] = 16'b1111111111111100;
    assign weights1[44][430] = 16'b1111111111110100;
    assign weights1[44][431] = 16'b0000000000001011;
    assign weights1[44][432] = 16'b1111111111110110;
    assign weights1[44][433] = 16'b1111111111111100;
    assign weights1[44][434] = 16'b1111111111111001;
    assign weights1[44][435] = 16'b0000000000000001;
    assign weights1[44][436] = 16'b0000000000000011;
    assign weights1[44][437] = 16'b0000000000010100;
    assign weights1[44][438] = 16'b1111111111111111;
    assign weights1[44][439] = 16'b1111111111111010;
    assign weights1[44][440] = 16'b0000000000000101;
    assign weights1[44][441] = 16'b1111111111011101;
    assign weights1[44][442] = 16'b1111111111100110;
    assign weights1[44][443] = 16'b1111111111111001;
    assign weights1[44][444] = 16'b1111111111101001;
    assign weights1[44][445] = 16'b0000000000000101;
    assign weights1[44][446] = 16'b0000000000000111;
    assign weights1[44][447] = 16'b0000000000000001;
    assign weights1[44][448] = 16'b0000000000001110;
    assign weights1[44][449] = 16'b0000000000011000;
    assign weights1[44][450] = 16'b0000000000010001;
    assign weights1[44][451] = 16'b0000000000001001;
    assign weights1[44][452] = 16'b0000000000000010;
    assign weights1[44][453] = 16'b0000000000001011;
    assign weights1[44][454] = 16'b1111111111110011;
    assign weights1[44][455] = 16'b0000000000000011;
    assign weights1[44][456] = 16'b1111111111110001;
    assign weights1[44][457] = 16'b1111111111110010;
    assign weights1[44][458] = 16'b0000000000000011;
    assign weights1[44][459] = 16'b1111111111110011;
    assign weights1[44][460] = 16'b1111111111101110;
    assign weights1[44][461] = 16'b1111111111011010;
    assign weights1[44][462] = 16'b1111111111011111;
    assign weights1[44][463] = 16'b1111111111100101;
    assign weights1[44][464] = 16'b1111111111111011;
    assign weights1[44][465] = 16'b0000000000000110;
    assign weights1[44][466] = 16'b0000000000000000;
    assign weights1[44][467] = 16'b1111111111110110;
    assign weights1[44][468] = 16'b1111111111111100;
    assign weights1[44][469] = 16'b0000000000001100;
    assign weights1[44][470] = 16'b1111111111110110;
    assign weights1[44][471] = 16'b1111111111100010;
    assign weights1[44][472] = 16'b0000000000000000;
    assign weights1[44][473] = 16'b1111111111111110;
    assign weights1[44][474] = 16'b1111111111111111;
    assign weights1[44][475] = 16'b0000000000001010;
    assign weights1[44][476] = 16'b0000000000001111;
    assign weights1[44][477] = 16'b0000000000010100;
    assign weights1[44][478] = 16'b0000000000011100;
    assign weights1[44][479] = 16'b0000000000001111;
    assign weights1[44][480] = 16'b0000000000000110;
    assign weights1[44][481] = 16'b1111111111111110;
    assign weights1[44][482] = 16'b1111111111111110;
    assign weights1[44][483] = 16'b1111111111110100;
    assign weights1[44][484] = 16'b0000000000000001;
    assign weights1[44][485] = 16'b1111111111100001;
    assign weights1[44][486] = 16'b1111111111110111;
    assign weights1[44][487] = 16'b1111111111100010;
    assign weights1[44][488] = 16'b0000000000000010;
    assign weights1[44][489] = 16'b1111111111111100;
    assign weights1[44][490] = 16'b1111111111111100;
    assign weights1[44][491] = 16'b0000000000000100;
    assign weights1[44][492] = 16'b1111111111110111;
    assign weights1[44][493] = 16'b1111111111111110;
    assign weights1[44][494] = 16'b1111111111110011;
    assign weights1[44][495] = 16'b1111111111110010;
    assign weights1[44][496] = 16'b1111111111110111;
    assign weights1[44][497] = 16'b1111111111110100;
    assign weights1[44][498] = 16'b1111111111110001;
    assign weights1[44][499] = 16'b1111111111011100;
    assign weights1[44][500] = 16'b1111111111110101;
    assign weights1[44][501] = 16'b0000000000000000;
    assign weights1[44][502] = 16'b1111111111111101;
    assign weights1[44][503] = 16'b0000000000001100;
    assign weights1[44][504] = 16'b0000000000001110;
    assign weights1[44][505] = 16'b0000000000011010;
    assign weights1[44][506] = 16'b0000000000001001;
    assign weights1[44][507] = 16'b0000000000001000;
    assign weights1[44][508] = 16'b0000000000000100;
    assign weights1[44][509] = 16'b0000000000011100;
    assign weights1[44][510] = 16'b0000000000001011;
    assign weights1[44][511] = 16'b0000000000001100;
    assign weights1[44][512] = 16'b0000000000000000;
    assign weights1[44][513] = 16'b0000000000001110;
    assign weights1[44][514] = 16'b0000000000000101;
    assign weights1[44][515] = 16'b0000000000001011;
    assign weights1[44][516] = 16'b1111111111110100;
    assign weights1[44][517] = 16'b1111111111111000;
    assign weights1[44][518] = 16'b1111111111101000;
    assign weights1[44][519] = 16'b1111111111100000;
    assign weights1[44][520] = 16'b0000000000001001;
    assign weights1[44][521] = 16'b1111111111111111;
    assign weights1[44][522] = 16'b0000000000010010;
    assign weights1[44][523] = 16'b0000000000001011;
    assign weights1[44][524] = 16'b1111111111110111;
    assign weights1[44][525] = 16'b0000000000001001;
    assign weights1[44][526] = 16'b1111111111111000;
    assign weights1[44][527] = 16'b1111111111110110;
    assign weights1[44][528] = 16'b0000000000100010;
    assign weights1[44][529] = 16'b0000000000010100;
    assign weights1[44][530] = 16'b0000000000000110;
    assign weights1[44][531] = 16'b0000000000001001;
    assign weights1[44][532] = 16'b0000000000001100;
    assign weights1[44][533] = 16'b0000000000001110;
    assign weights1[44][534] = 16'b0000000000010000;
    assign weights1[44][535] = 16'b0000000000001110;
    assign weights1[44][536] = 16'b1111111111111010;
    assign weights1[44][537] = 16'b0000000000011001;
    assign weights1[44][538] = 16'b0000000000000011;
    assign weights1[44][539] = 16'b1111111111111111;
    assign weights1[44][540] = 16'b0000000000010000;
    assign weights1[44][541] = 16'b1111111111111000;
    assign weights1[44][542] = 16'b1111111111111001;
    assign weights1[44][543] = 16'b1111111111111000;
    assign weights1[44][544] = 16'b0000000000001110;
    assign weights1[44][545] = 16'b1111111111110100;
    assign weights1[44][546] = 16'b1111111111111100;
    assign weights1[44][547] = 16'b1111111111101011;
    assign weights1[44][548] = 16'b1111111111110101;
    assign weights1[44][549] = 16'b0000000000001111;
    assign weights1[44][550] = 16'b0000000000000010;
    assign weights1[44][551] = 16'b1111111111111010;
    assign weights1[44][552] = 16'b0000000000001101;
    assign weights1[44][553] = 16'b0000000000001010;
    assign weights1[44][554] = 16'b1111111111111011;
    assign weights1[44][555] = 16'b0000000000000110;
    assign weights1[44][556] = 16'b1111111111111100;
    assign weights1[44][557] = 16'b1111111111111110;
    assign weights1[44][558] = 16'b0000000000000110;
    assign weights1[44][559] = 16'b0000000000000100;
    assign weights1[44][560] = 16'b0000000000010010;
    assign weights1[44][561] = 16'b0000000000011011;
    assign weights1[44][562] = 16'b0000000000001001;
    assign weights1[44][563] = 16'b0000000000000001;
    assign weights1[44][564] = 16'b0000000000010111;
    assign weights1[44][565] = 16'b1111111111110011;
    assign weights1[44][566] = 16'b0000000000000000;
    assign weights1[44][567] = 16'b0000000000010111;
    assign weights1[44][568] = 16'b0000000000000000;
    assign weights1[44][569] = 16'b1111111111101100;
    assign weights1[44][570] = 16'b1111111111110111;
    assign weights1[44][571] = 16'b0000000000000001;
    assign weights1[44][572] = 16'b0000000000000000;
    assign weights1[44][573] = 16'b0000000000001000;
    assign weights1[44][574] = 16'b0000000000010000;
    assign weights1[44][575] = 16'b1111111111111001;
    assign weights1[44][576] = 16'b1111111111111000;
    assign weights1[44][577] = 16'b1111111111110110;
    assign weights1[44][578] = 16'b1111111111111110;
    assign weights1[44][579] = 16'b0000000000010011;
    assign weights1[44][580] = 16'b1111111111111011;
    assign weights1[44][581] = 16'b1111111111110101;
    assign weights1[44][582] = 16'b1111111111111100;
    assign weights1[44][583] = 16'b0000000000010011;
    assign weights1[44][584] = 16'b0000000000010111;
    assign weights1[44][585] = 16'b0000000000000001;
    assign weights1[44][586] = 16'b1111111111111000;
    assign weights1[44][587] = 16'b1111111111111110;
    assign weights1[44][588] = 16'b0000000000100000;
    assign weights1[44][589] = 16'b0000000000010011;
    assign weights1[44][590] = 16'b0000000000010100;
    assign weights1[44][591] = 16'b1111111111111110;
    assign weights1[44][592] = 16'b0000000000001100;
    assign weights1[44][593] = 16'b1111111111110111;
    assign weights1[44][594] = 16'b0000000000000111;
    assign weights1[44][595] = 16'b0000000000010001;
    assign weights1[44][596] = 16'b0000000000001100;
    assign weights1[44][597] = 16'b0000000000000000;
    assign weights1[44][598] = 16'b0000000000011001;
    assign weights1[44][599] = 16'b1111111111111101;
    assign weights1[44][600] = 16'b1111111111110000;
    assign weights1[44][601] = 16'b1111111111110101;
    assign weights1[44][602] = 16'b1111111111111010;
    assign weights1[44][603] = 16'b1111111111110000;
    assign weights1[44][604] = 16'b1111111111100101;
    assign weights1[44][605] = 16'b1111111111110010;
    assign weights1[44][606] = 16'b1111111111100110;
    assign weights1[44][607] = 16'b1111111111111111;
    assign weights1[44][608] = 16'b0000000000000010;
    assign weights1[44][609] = 16'b1111111111111001;
    assign weights1[44][610] = 16'b0000000000000011;
    assign weights1[44][611] = 16'b1111111111111000;
    assign weights1[44][612] = 16'b1111111111111110;
    assign weights1[44][613] = 16'b1111111111110011;
    assign weights1[44][614] = 16'b1111111111110110;
    assign weights1[44][615] = 16'b0000000000000101;
    assign weights1[44][616] = 16'b0000000000001110;
    assign weights1[44][617] = 16'b0000000000010000;
    assign weights1[44][618] = 16'b0000000000000010;
    assign weights1[44][619] = 16'b0000000000001000;
    assign weights1[44][620] = 16'b0000000000000001;
    assign weights1[44][621] = 16'b0000000000011110;
    assign weights1[44][622] = 16'b0000000000010100;
    assign weights1[44][623] = 16'b0000000000000010;
    assign weights1[44][624] = 16'b0000000000000001;
    assign weights1[44][625] = 16'b1111111111111010;
    assign weights1[44][626] = 16'b0000000000001111;
    assign weights1[44][627] = 16'b1111111111110101;
    assign weights1[44][628] = 16'b0000000000000110;
    assign weights1[44][629] = 16'b1111111111101101;
    assign weights1[44][630] = 16'b0000000000001110;
    assign weights1[44][631] = 16'b0000000000000111;
    assign weights1[44][632] = 16'b1111111111111000;
    assign weights1[44][633] = 16'b0000000000000111;
    assign weights1[44][634] = 16'b1111111111110111;
    assign weights1[44][635] = 16'b0000000000000000;
    assign weights1[44][636] = 16'b1111111111100011;
    assign weights1[44][637] = 16'b0000000000010010;
    assign weights1[44][638] = 16'b0000000000001111;
    assign weights1[44][639] = 16'b1111111111110110;
    assign weights1[44][640] = 16'b0000000000000000;
    assign weights1[44][641] = 16'b1111111111111111;
    assign weights1[44][642] = 16'b1111111111111101;
    assign weights1[44][643] = 16'b0000000000000011;
    assign weights1[44][644] = 16'b0000000000010011;
    assign weights1[44][645] = 16'b0000000000001100;
    assign weights1[44][646] = 16'b0000000000001100;
    assign weights1[44][647] = 16'b1111111111111011;
    assign weights1[44][648] = 16'b1111111111110101;
    assign weights1[44][649] = 16'b1111111111101010;
    assign weights1[44][650] = 16'b0000000000001101;
    assign weights1[44][651] = 16'b0000000000100101;
    assign weights1[44][652] = 16'b0000000000000111;
    assign weights1[44][653] = 16'b1111111111101100;
    assign weights1[44][654] = 16'b0000000000010100;
    assign weights1[44][655] = 16'b1111111111110101;
    assign weights1[44][656] = 16'b0000000000010000;
    assign weights1[44][657] = 16'b1111111111111110;
    assign weights1[44][658] = 16'b1111111111101000;
    assign weights1[44][659] = 16'b1111111111101011;
    assign weights1[44][660] = 16'b1111111111101101;
    assign weights1[44][661] = 16'b1111111111100100;
    assign weights1[44][662] = 16'b1111111111111000;
    assign weights1[44][663] = 16'b1111111111110010;
    assign weights1[44][664] = 16'b1111111111101100;
    assign weights1[44][665] = 16'b0000000000001010;
    assign weights1[44][666] = 16'b0000000000000110;
    assign weights1[44][667] = 16'b1111111111111101;
    assign weights1[44][668] = 16'b1111111111101011;
    assign weights1[44][669] = 16'b0000000000000011;
    assign weights1[44][670] = 16'b0000000000000100;
    assign weights1[44][671] = 16'b0000000000000110;
    assign weights1[44][672] = 16'b0000000000010010;
    assign weights1[44][673] = 16'b0000000000001110;
    assign weights1[44][674] = 16'b0000000000001011;
    assign weights1[44][675] = 16'b0000000000000001;
    assign weights1[44][676] = 16'b0000000000010011;
    assign weights1[44][677] = 16'b0000000000010110;
    assign weights1[44][678] = 16'b0000000000000011;
    assign weights1[44][679] = 16'b0000000000010001;
    assign weights1[44][680] = 16'b1111111111101001;
    assign weights1[44][681] = 16'b1111111111111011;
    assign weights1[44][682] = 16'b0000000000010010;
    assign weights1[44][683] = 16'b1111111111110110;
    assign weights1[44][684] = 16'b1111111111101110;
    assign weights1[44][685] = 16'b0000000000001101;
    assign weights1[44][686] = 16'b1111111111100111;
    assign weights1[44][687] = 16'b1111111111111100;
    assign weights1[44][688] = 16'b0000000000000111;
    assign weights1[44][689] = 16'b0000000000001111;
    assign weights1[44][690] = 16'b1111111111100110;
    assign weights1[44][691] = 16'b1111111111101110;
    assign weights1[44][692] = 16'b1111111111110111;
    assign weights1[44][693] = 16'b1111111111111111;
    assign weights1[44][694] = 16'b1111111111110001;
    assign weights1[44][695] = 16'b1111111111110111;
    assign weights1[44][696] = 16'b1111111111111001;
    assign weights1[44][697] = 16'b0000000000000111;
    assign weights1[44][698] = 16'b0000000000000011;
    assign weights1[44][699] = 16'b0000000000000011;
    assign weights1[44][700] = 16'b0000000000001010;
    assign weights1[44][701] = 16'b0000000000010101;
    assign weights1[44][702] = 16'b0000000000011001;
    assign weights1[44][703] = 16'b0000000000001000;
    assign weights1[44][704] = 16'b0000000000001010;
    assign weights1[44][705] = 16'b0000000000010001;
    assign weights1[44][706] = 16'b0000000000000100;
    assign weights1[44][707] = 16'b1111111111111101;
    assign weights1[44][708] = 16'b0000000000000010;
    assign weights1[44][709] = 16'b0000000000011001;
    assign weights1[44][710] = 16'b0000000000001110;
    assign weights1[44][711] = 16'b0000000000010111;
    assign weights1[44][712] = 16'b0000000000010101;
    assign weights1[44][713] = 16'b0000000000011010;
    assign weights1[44][714] = 16'b0000000000000011;
    assign weights1[44][715] = 16'b0000000000000000;
    assign weights1[44][716] = 16'b1111111111111110;
    assign weights1[44][717] = 16'b0000000000001110;
    assign weights1[44][718] = 16'b0000000000001010;
    assign weights1[44][719] = 16'b1111111111110100;
    assign weights1[44][720] = 16'b1111111111110010;
    assign weights1[44][721] = 16'b0000000000000111;
    assign weights1[44][722] = 16'b0000000000001010;
    assign weights1[44][723] = 16'b1111111111111000;
    assign weights1[44][724] = 16'b1111111111111101;
    assign weights1[44][725] = 16'b1111111111110111;
    assign weights1[44][726] = 16'b1111111111111111;
    assign weights1[44][727] = 16'b0000000000000001;
    assign weights1[44][728] = 16'b0000000000000101;
    assign weights1[44][729] = 16'b0000000000010010;
    assign weights1[44][730] = 16'b0000000000011000;
    assign weights1[44][731] = 16'b0000000000011001;
    assign weights1[44][732] = 16'b0000000000010101;
    assign weights1[44][733] = 16'b1111111111111000;
    assign weights1[44][734] = 16'b1111111111111100;
    assign weights1[44][735] = 16'b0000000000000110;
    assign weights1[44][736] = 16'b0000000000001010;
    assign weights1[44][737] = 16'b1111111111111001;
    assign weights1[44][738] = 16'b0000000000010110;
    assign weights1[44][739] = 16'b1111111111100111;
    assign weights1[44][740] = 16'b1111111111110011;
    assign weights1[44][741] = 16'b1111111111111101;
    assign weights1[44][742] = 16'b0000000000001111;
    assign weights1[44][743] = 16'b1111111111100010;
    assign weights1[44][744] = 16'b1111111111111101;
    assign weights1[44][745] = 16'b0000000000001001;
    assign weights1[44][746] = 16'b0000000000001001;
    assign weights1[44][747] = 16'b1111111111101111;
    assign weights1[44][748] = 16'b1111111111111001;
    assign weights1[44][749] = 16'b0000000000000101;
    assign weights1[44][750] = 16'b0000000000000110;
    assign weights1[44][751] = 16'b0000000000000010;
    assign weights1[44][752] = 16'b0000000000000000;
    assign weights1[44][753] = 16'b1111111111111011;
    assign weights1[44][754] = 16'b0000000000000000;
    assign weights1[44][755] = 16'b0000000000000010;
    assign weights1[44][756] = 16'b0000000000000001;
    assign weights1[44][757] = 16'b0000000000001011;
    assign weights1[44][758] = 16'b0000000000001010;
    assign weights1[44][759] = 16'b0000000000001111;
    assign weights1[44][760] = 16'b0000000000000011;
    assign weights1[44][761] = 16'b1111111111111001;
    assign weights1[44][762] = 16'b0000000000000101;
    assign weights1[44][763] = 16'b0000000000000111;
    assign weights1[44][764] = 16'b0000000000000110;
    assign weights1[44][765] = 16'b0000000000000100;
    assign weights1[44][766] = 16'b0000000000001111;
    assign weights1[44][767] = 16'b0000000000000010;
    assign weights1[44][768] = 16'b0000000000001111;
    assign weights1[44][769] = 16'b0000000000001000;
    assign weights1[44][770] = 16'b0000000000001001;
    assign weights1[44][771] = 16'b0000000000001111;
    assign weights1[44][772] = 16'b0000000000000011;
    assign weights1[44][773] = 16'b0000000000000000;
    assign weights1[44][774] = 16'b1111111111110101;
    assign weights1[44][775] = 16'b1111111111111101;
    assign weights1[44][776] = 16'b0000000000000000;
    assign weights1[44][777] = 16'b0000000000000000;
    assign weights1[44][778] = 16'b1111111111110100;
    assign weights1[44][779] = 16'b0000000000000000;
    assign weights1[44][780] = 16'b0000000000000001;
    assign weights1[44][781] = 16'b0000000000000000;
    assign weights1[44][782] = 16'b0000000000000011;
    assign weights1[44][783] = 16'b0000000000000010;
    assign weights1[45][0] = 16'b0000000000000000;
    assign weights1[45][1] = 16'b0000000000000000;
    assign weights1[45][2] = 16'b0000000000000000;
    assign weights1[45][3] = 16'b1111111111111111;
    assign weights1[45][4] = 16'b1111111111111111;
    assign weights1[45][5] = 16'b1111111111111001;
    assign weights1[45][6] = 16'b1111111111110101;
    assign weights1[45][7] = 16'b1111111111110100;
    assign weights1[45][8] = 16'b1111111111101110;
    assign weights1[45][9] = 16'b1111111111011101;
    assign weights1[45][10] = 16'b1111111111001011;
    assign weights1[45][11] = 16'b1111111111001010;
    assign weights1[45][12] = 16'b1111111111010000;
    assign weights1[45][13] = 16'b1111111111110010;
    assign weights1[45][14] = 16'b0000000000010001;
    assign weights1[45][15] = 16'b0000000000011001;
    assign weights1[45][16] = 16'b0000000000100111;
    assign weights1[45][17] = 16'b0000000000110000;
    assign weights1[45][18] = 16'b0000000000011110;
    assign weights1[45][19] = 16'b0000000000011110;
    assign weights1[45][20] = 16'b0000000000100001;
    assign weights1[45][21] = 16'b0000000000001001;
    assign weights1[45][22] = 16'b1111111111111111;
    assign weights1[45][23] = 16'b1111111111111101;
    assign weights1[45][24] = 16'b0000000000000001;
    assign weights1[45][25] = 16'b1111111111111110;
    assign weights1[45][26] = 16'b1111111111111101;
    assign weights1[45][27] = 16'b1111111111111100;
    assign weights1[45][28] = 16'b0000000000000000;
    assign weights1[45][29] = 16'b0000000000000000;
    assign weights1[45][30] = 16'b0000000000000000;
    assign weights1[45][31] = 16'b0000000000000001;
    assign weights1[45][32] = 16'b1111111111111011;
    assign weights1[45][33] = 16'b1111111111110101;
    assign weights1[45][34] = 16'b1111111111110100;
    assign weights1[45][35] = 16'b1111111111101000;
    assign weights1[45][36] = 16'b1111111111100000;
    assign weights1[45][37] = 16'b1111111111010101;
    assign weights1[45][38] = 16'b1111111111000111;
    assign weights1[45][39] = 16'b1111111110111111;
    assign weights1[45][40] = 16'b1111111111100101;
    assign weights1[45][41] = 16'b1111111111101100;
    assign weights1[45][42] = 16'b0000000000000110;
    assign weights1[45][43] = 16'b0000000000011010;
    assign weights1[45][44] = 16'b0000000000100101;
    assign weights1[45][45] = 16'b0000000000011011;
    assign weights1[45][46] = 16'b0000000000011101;
    assign weights1[45][47] = 16'b0000000000010010;
    assign weights1[45][48] = 16'b0000000000001110;
    assign weights1[45][49] = 16'b0000000000000111;
    assign weights1[45][50] = 16'b0000000000001001;
    assign weights1[45][51] = 16'b0000000000000100;
    assign weights1[45][52] = 16'b0000000000000000;
    assign weights1[45][53] = 16'b1111111111110110;
    assign weights1[45][54] = 16'b1111111111110110;
    assign weights1[45][55] = 16'b1111111111111100;
    assign weights1[45][56] = 16'b0000000000000000;
    assign weights1[45][57] = 16'b0000000000000000;
    assign weights1[45][58] = 16'b1111111111111110;
    assign weights1[45][59] = 16'b1111111111111111;
    assign weights1[45][60] = 16'b1111111111111011;
    assign weights1[45][61] = 16'b1111111111111000;
    assign weights1[45][62] = 16'b1111111111101010;
    assign weights1[45][63] = 16'b1111111111100001;
    assign weights1[45][64] = 16'b1111111111010001;
    assign weights1[45][65] = 16'b1111111111010011;
    assign weights1[45][66] = 16'b1111111111000000;
    assign weights1[45][67] = 16'b1111111111011101;
    assign weights1[45][68] = 16'b0000000000010001;
    assign weights1[45][69] = 16'b0000000000010110;
    assign weights1[45][70] = 16'b0000000000010110;
    assign weights1[45][71] = 16'b0000000000100000;
    assign weights1[45][72] = 16'b0000000000010111;
    assign weights1[45][73] = 16'b0000000000011010;
    assign weights1[45][74] = 16'b0000000000001011;
    assign weights1[45][75] = 16'b0000000000011100;
    assign weights1[45][76] = 16'b0000000000001111;
    assign weights1[45][77] = 16'b1111111111111101;
    assign weights1[45][78] = 16'b1111111111111000;
    assign weights1[45][79] = 16'b1111111111101111;
    assign weights1[45][80] = 16'b1111111111101011;
    assign weights1[45][81] = 16'b1111111111101111;
    assign weights1[45][82] = 16'b1111111111110010;
    assign weights1[45][83] = 16'b1111111111111000;
    assign weights1[45][84] = 16'b0000000000000000;
    assign weights1[45][85] = 16'b0000000000000000;
    assign weights1[45][86] = 16'b0000000000000000;
    assign weights1[45][87] = 16'b1111111111111011;
    assign weights1[45][88] = 16'b1111111111110101;
    assign weights1[45][89] = 16'b1111111111110000;
    assign weights1[45][90] = 16'b1111111111101011;
    assign weights1[45][91] = 16'b1111111111010111;
    assign weights1[45][92] = 16'b1111111111001100;
    assign weights1[45][93] = 16'b1111111111000011;
    assign weights1[45][94] = 16'b1111111110111010;
    assign weights1[45][95] = 16'b0000000000000010;
    assign weights1[45][96] = 16'b0000000000010001;
    assign weights1[45][97] = 16'b0000000000011010;
    assign weights1[45][98] = 16'b0000000000011000;
    assign weights1[45][99] = 16'b0000000000101011;
    assign weights1[45][100] = 16'b0000000000101011;
    assign weights1[45][101] = 16'b0000000000100111;
    assign weights1[45][102] = 16'b0000000000011000;
    assign weights1[45][103] = 16'b0000000000010011;
    assign weights1[45][104] = 16'b1111111111011100;
    assign weights1[45][105] = 16'b1111111111011000;
    assign weights1[45][106] = 16'b1111111111010101;
    assign weights1[45][107] = 16'b1111111111011000;
    assign weights1[45][108] = 16'b1111111111010001;
    assign weights1[45][109] = 16'b1111111111100011;
    assign weights1[45][110] = 16'b1111111111101000;
    assign weights1[45][111] = 16'b1111111111110101;
    assign weights1[45][112] = 16'b0000000000000000;
    assign weights1[45][113] = 16'b0000000000000000;
    assign weights1[45][114] = 16'b0000000000000000;
    assign weights1[45][115] = 16'b1111111111111010;
    assign weights1[45][116] = 16'b1111111111101111;
    assign weights1[45][117] = 16'b1111111111100100;
    assign weights1[45][118] = 16'b1111111111011010;
    assign weights1[45][119] = 16'b1111111111000111;
    assign weights1[45][120] = 16'b1111111110100110;
    assign weights1[45][121] = 16'b1111111110111110;
    assign weights1[45][122] = 16'b1111111111001010;
    assign weights1[45][123] = 16'b0000000000000101;
    assign weights1[45][124] = 16'b1111111111111010;
    assign weights1[45][125] = 16'b0000000000010100;
    assign weights1[45][126] = 16'b1111111111111101;
    assign weights1[45][127] = 16'b0000000000011001;
    assign weights1[45][128] = 16'b0000000000001110;
    assign weights1[45][129] = 16'b0000000000011111;
    assign weights1[45][130] = 16'b0000000000010000;
    assign weights1[45][131] = 16'b1111111111101101;
    assign weights1[45][132] = 16'b1111111111000100;
    assign weights1[45][133] = 16'b1111111111001110;
    assign weights1[45][134] = 16'b1111111110111000;
    assign weights1[45][135] = 16'b1111111110101001;
    assign weights1[45][136] = 16'b1111111111000001;
    assign weights1[45][137] = 16'b1111111111100000;
    assign weights1[45][138] = 16'b1111111111100110;
    assign weights1[45][139] = 16'b1111111111110101;
    assign weights1[45][140] = 16'b1111111111111111;
    assign weights1[45][141] = 16'b1111111111111011;
    assign weights1[45][142] = 16'b1111111111110110;
    assign weights1[45][143] = 16'b1111111111110100;
    assign weights1[45][144] = 16'b1111111111101011;
    assign weights1[45][145] = 16'b1111111111011011;
    assign weights1[45][146] = 16'b1111111111010100;
    assign weights1[45][147] = 16'b1111111110101001;
    assign weights1[45][148] = 16'b1111111110110100;
    assign weights1[45][149] = 16'b1111111111011010;
    assign weights1[45][150] = 16'b0000000000000100;
    assign weights1[45][151] = 16'b0000000001000010;
    assign weights1[45][152] = 16'b0000000000011010;
    assign weights1[45][153] = 16'b0000000000001000;
    assign weights1[45][154] = 16'b0000000000011001;
    assign weights1[45][155] = 16'b0000000000010110;
    assign weights1[45][156] = 16'b0000000000001010;
    assign weights1[45][157] = 16'b0000000000011101;
    assign weights1[45][158] = 16'b1111111111101101;
    assign weights1[45][159] = 16'b1111111111100011;
    assign weights1[45][160] = 16'b1111111111010100;
    assign weights1[45][161] = 16'b1111111111001000;
    assign weights1[45][162] = 16'b1111111110101010;
    assign weights1[45][163] = 16'b1111111111000011;
    assign weights1[45][164] = 16'b1111111111011010;
    assign weights1[45][165] = 16'b1111111111101010;
    assign weights1[45][166] = 16'b1111111111101111;
    assign weights1[45][167] = 16'b1111111111110100;
    assign weights1[45][168] = 16'b1111111111111110;
    assign weights1[45][169] = 16'b1111111111111001;
    assign weights1[45][170] = 16'b1111111111110010;
    assign weights1[45][171] = 16'b1111111111101011;
    assign weights1[45][172] = 16'b1111111111100011;
    assign weights1[45][173] = 16'b1111111111010100;
    assign weights1[45][174] = 16'b1111111110111110;
    assign weights1[45][175] = 16'b1111111110110000;
    assign weights1[45][176] = 16'b1111111110100000;
    assign weights1[45][177] = 16'b1111111111011010;
    assign weights1[45][178] = 16'b0000000000010100;
    assign weights1[45][179] = 16'b0000000000010100;
    assign weights1[45][180] = 16'b0000000000000001;
    assign weights1[45][181] = 16'b0000000000011101;
    assign weights1[45][182] = 16'b0000000000011101;
    assign weights1[45][183] = 16'b1111111111101111;
    assign weights1[45][184] = 16'b1111111111011101;
    assign weights1[45][185] = 16'b1111111111110100;
    assign weights1[45][186] = 16'b1111111110111101;
    assign weights1[45][187] = 16'b1111111111010110;
    assign weights1[45][188] = 16'b1111111111011010;
    assign weights1[45][189] = 16'b1111111111011101;
    assign weights1[45][190] = 16'b1111111111100110;
    assign weights1[45][191] = 16'b1111111111111001;
    assign weights1[45][192] = 16'b1111111111110110;
    assign weights1[45][193] = 16'b1111111111101000;
    assign weights1[45][194] = 16'b1111111111111101;
    assign weights1[45][195] = 16'b1111111111110000;
    assign weights1[45][196] = 16'b1111111111111110;
    assign weights1[45][197] = 16'b1111111111111010;
    assign weights1[45][198] = 16'b1111111111110110;
    assign weights1[45][199] = 16'b1111111111101101;
    assign weights1[45][200] = 16'b1111111111101110;
    assign weights1[45][201] = 16'b1111111111011010;
    assign weights1[45][202] = 16'b1111111110111111;
    assign weights1[45][203] = 16'b1111111110101011;
    assign weights1[45][204] = 16'b1111111110110001;
    assign weights1[45][205] = 16'b0000000000010110;
    assign weights1[45][206] = 16'b0000000000011101;
    assign weights1[45][207] = 16'b0000000000110010;
    assign weights1[45][208] = 16'b0000000000001101;
    assign weights1[45][209] = 16'b0000000000001111;
    assign weights1[45][210] = 16'b0000000000001110;
    assign weights1[45][211] = 16'b1111111111111101;
    assign weights1[45][212] = 16'b1111111111100111;
    assign weights1[45][213] = 16'b1111111111011010;
    assign weights1[45][214] = 16'b1111111111101000;
    assign weights1[45][215] = 16'b1111111111011110;
    assign weights1[45][216] = 16'b1111111111101101;
    assign weights1[45][217] = 16'b1111111111011110;
    assign weights1[45][218] = 16'b1111111111110011;
    assign weights1[45][219] = 16'b1111111111110001;
    assign weights1[45][220] = 16'b0000000000000110;
    assign weights1[45][221] = 16'b0000000000000100;
    assign weights1[45][222] = 16'b1111111111111101;
    assign weights1[45][223] = 16'b1111111111110111;
    assign weights1[45][224] = 16'b1111111111111101;
    assign weights1[45][225] = 16'b1111111111110110;
    assign weights1[45][226] = 16'b1111111111110001;
    assign weights1[45][227] = 16'b1111111111101001;
    assign weights1[45][228] = 16'b1111111111100111;
    assign weights1[45][229] = 16'b1111111111010011;
    assign weights1[45][230] = 16'b1111111111000001;
    assign weights1[45][231] = 16'b1111111110011001;
    assign weights1[45][232] = 16'b1111111111001100;
    assign weights1[45][233] = 16'b0000000000000111;
    assign weights1[45][234] = 16'b0000000000001010;
    assign weights1[45][235] = 16'b0000000000011101;
    assign weights1[45][236] = 16'b0000000000001111;
    assign weights1[45][237] = 16'b0000000000010101;
    assign weights1[45][238] = 16'b0000000000000111;
    assign weights1[45][239] = 16'b1111111111011010;
    assign weights1[45][240] = 16'b1111111111001111;
    assign weights1[45][241] = 16'b1111111111010010;
    assign weights1[45][242] = 16'b1111111111011001;
    assign weights1[45][243] = 16'b1111111111100001;
    assign weights1[45][244] = 16'b1111111111101111;
    assign weights1[45][245] = 16'b1111111111111011;
    assign weights1[45][246] = 16'b1111111111111101;
    assign weights1[45][247] = 16'b0000000000000101;
    assign weights1[45][248] = 16'b0000000000001110;
    assign weights1[45][249] = 16'b0000000000000000;
    assign weights1[45][250] = 16'b0000000000001000;
    assign weights1[45][251] = 16'b0000000000000000;
    assign weights1[45][252] = 16'b0000000000000000;
    assign weights1[45][253] = 16'b1111111111111100;
    assign weights1[45][254] = 16'b1111111111110011;
    assign weights1[45][255] = 16'b1111111111101010;
    assign weights1[45][256] = 16'b1111111111100101;
    assign weights1[45][257] = 16'b1111111111000110;
    assign weights1[45][258] = 16'b1111111110101001;
    assign weights1[45][259] = 16'b1111111110011100;
    assign weights1[45][260] = 16'b1111111111111001;
    assign weights1[45][261] = 16'b0000000000010001;
    assign weights1[45][262] = 16'b0000000000001110;
    assign weights1[45][263] = 16'b0000000000000100;
    assign weights1[45][264] = 16'b0000000000001111;
    assign weights1[45][265] = 16'b0000000000000111;
    assign weights1[45][266] = 16'b1111111111100100;
    assign weights1[45][267] = 16'b1111111111000100;
    assign weights1[45][268] = 16'b1111111111011101;
    assign weights1[45][269] = 16'b1111111111100101;
    assign weights1[45][270] = 16'b1111111111100001;
    assign weights1[45][271] = 16'b1111111111110010;
    assign weights1[45][272] = 16'b1111111111110010;
    assign weights1[45][273] = 16'b0000000000011101;
    assign weights1[45][274] = 16'b0000000000001011;
    assign weights1[45][275] = 16'b0000000000011001;
    assign weights1[45][276] = 16'b0000000000010001;
    assign weights1[45][277] = 16'b0000000000001010;
    assign weights1[45][278] = 16'b0000000000001011;
    assign weights1[45][279] = 16'b0000000000001000;
    assign weights1[45][280] = 16'b1111111111111110;
    assign weights1[45][281] = 16'b1111111111110110;
    assign weights1[45][282] = 16'b1111111111110010;
    assign weights1[45][283] = 16'b1111111111101100;
    assign weights1[45][284] = 16'b1111111111011010;
    assign weights1[45][285] = 16'b1111111111000101;
    assign weights1[45][286] = 16'b1111111110010111;
    assign weights1[45][287] = 16'b1111111111110010;
    assign weights1[45][288] = 16'b1111111111101001;
    assign weights1[45][289] = 16'b0000000000011001;
    assign weights1[45][290] = 16'b0000000000001011;
    assign weights1[45][291] = 16'b0000000000011110;
    assign weights1[45][292] = 16'b0000000000001001;
    assign weights1[45][293] = 16'b0000000000000111;
    assign weights1[45][294] = 16'b1111111111011010;
    assign weights1[45][295] = 16'b1111111111000101;
    assign weights1[45][296] = 16'b1111111111110101;
    assign weights1[45][297] = 16'b1111111111111111;
    assign weights1[45][298] = 16'b1111111111111111;
    assign weights1[45][299] = 16'b1111111111110100;
    assign weights1[45][300] = 16'b0000000000001100;
    assign weights1[45][301] = 16'b0000000000010100;
    assign weights1[45][302] = 16'b0000000000011001;
    assign weights1[45][303] = 16'b0000000000000100;
    assign weights1[45][304] = 16'b0000000000000011;
    assign weights1[45][305] = 16'b1111111111101011;
    assign weights1[45][306] = 16'b0000000000000111;
    assign weights1[45][307] = 16'b0000000000000100;
    assign weights1[45][308] = 16'b1111111111111111;
    assign weights1[45][309] = 16'b1111111111111010;
    assign weights1[45][310] = 16'b1111111111110011;
    assign weights1[45][311] = 16'b1111111111110010;
    assign weights1[45][312] = 16'b1111111111010110;
    assign weights1[45][313] = 16'b1111111110111101;
    assign weights1[45][314] = 16'b1111111111001100;
    assign weights1[45][315] = 16'b1111111111101100;
    assign weights1[45][316] = 16'b1111111111110110;
    assign weights1[45][317] = 16'b0000000000001010;
    assign weights1[45][318] = 16'b0000000000000010;
    assign weights1[45][319] = 16'b0000000000011110;
    assign weights1[45][320] = 16'b0000000000100100;
    assign weights1[45][321] = 16'b1111111111101100;
    assign weights1[45][322] = 16'b1111111111000001;
    assign weights1[45][323] = 16'b1111111111001011;
    assign weights1[45][324] = 16'b0000000000001000;
    assign weights1[45][325] = 16'b1111111111101000;
    assign weights1[45][326] = 16'b1111111111111100;
    assign weights1[45][327] = 16'b0000000000010011;
    assign weights1[45][328] = 16'b0000000000001100;
    assign weights1[45][329] = 16'b1111111111111100;
    assign weights1[45][330] = 16'b0000000000001111;
    assign weights1[45][331] = 16'b0000000000001011;
    assign weights1[45][332] = 16'b1111111111110001;
    assign weights1[45][333] = 16'b0000000000001010;
    assign weights1[45][334] = 16'b0000000000010011;
    assign weights1[45][335] = 16'b0000000000001001;
    assign weights1[45][336] = 16'b1111111111111111;
    assign weights1[45][337] = 16'b1111111111111011;
    assign weights1[45][338] = 16'b1111111111110100;
    assign weights1[45][339] = 16'b1111111111100111;
    assign weights1[45][340] = 16'b1111111111010010;
    assign weights1[45][341] = 16'b1111111111000111;
    assign weights1[45][342] = 16'b1111111111100101;
    assign weights1[45][343] = 16'b1111111111101110;
    assign weights1[45][344] = 16'b0000000000001011;
    assign weights1[45][345] = 16'b0000000000001110;
    assign weights1[45][346] = 16'b1111111111111110;
    assign weights1[45][347] = 16'b0000000000101110;
    assign weights1[45][348] = 16'b0000000000010010;
    assign weights1[45][349] = 16'b1111111111101111;
    assign weights1[45][350] = 16'b1111111111000010;
    assign weights1[45][351] = 16'b1111111111110001;
    assign weights1[45][352] = 16'b1111111111111101;
    assign weights1[45][353] = 16'b0000000000000000;
    assign weights1[45][354] = 16'b1111111111111110;
    assign weights1[45][355] = 16'b1111111111110101;
    assign weights1[45][356] = 16'b1111111111111001;
    assign weights1[45][357] = 16'b0000000000000010;
    assign weights1[45][358] = 16'b0000000000000001;
    assign weights1[45][359] = 16'b1111111111111111;
    assign weights1[45][360] = 16'b0000000000010001;
    assign weights1[45][361] = 16'b1111111111101100;
    assign weights1[45][362] = 16'b0000000000000000;
    assign weights1[45][363] = 16'b0000000000001100;
    assign weights1[45][364] = 16'b1111111111111110;
    assign weights1[45][365] = 16'b1111111111110101;
    assign weights1[45][366] = 16'b1111111111101111;
    assign weights1[45][367] = 16'b1111111111100001;
    assign weights1[45][368] = 16'b1111111111100100;
    assign weights1[45][369] = 16'b1111111111010100;
    assign weights1[45][370] = 16'b1111111111110100;
    assign weights1[45][371] = 16'b0000000000011001;
    assign weights1[45][372] = 16'b1111111111111011;
    assign weights1[45][373] = 16'b0000000000000001;
    assign weights1[45][374] = 16'b0000000000011000;
    assign weights1[45][375] = 16'b0000000000101000;
    assign weights1[45][376] = 16'b0000000000000110;
    assign weights1[45][377] = 16'b1111111111100100;
    assign weights1[45][378] = 16'b1111111111001101;
    assign weights1[45][379] = 16'b1111111111110111;
    assign weights1[45][380] = 16'b1111111111110111;
    assign weights1[45][381] = 16'b0000000000000010;
    assign weights1[45][382] = 16'b1111111111110101;
    assign weights1[45][383] = 16'b0000000000011011;
    assign weights1[45][384] = 16'b1111111111111101;
    assign weights1[45][385] = 16'b0000000000011111;
    assign weights1[45][386] = 16'b0000000000001101;
    assign weights1[45][387] = 16'b1111111111110000;
    assign weights1[45][388] = 16'b0000000000001111;
    assign weights1[45][389] = 16'b0000000000001011;
    assign weights1[45][390] = 16'b0000000000000110;
    assign weights1[45][391] = 16'b1111111111111111;
    assign weights1[45][392] = 16'b1111111111111000;
    assign weights1[45][393] = 16'b1111111111110100;
    assign weights1[45][394] = 16'b1111111111110000;
    assign weights1[45][395] = 16'b1111111111100000;
    assign weights1[45][396] = 16'b1111111111001011;
    assign weights1[45][397] = 16'b1111111111100111;
    assign weights1[45][398] = 16'b0000000000000110;
    assign weights1[45][399] = 16'b0000000000001100;
    assign weights1[45][400] = 16'b0000000000001011;
    assign weights1[45][401] = 16'b0000000000010000;
    assign weights1[45][402] = 16'b0000000000010110;
    assign weights1[45][403] = 16'b0000000000100110;
    assign weights1[45][404] = 16'b0000000000000011;
    assign weights1[45][405] = 16'b1111111111101010;
    assign weights1[45][406] = 16'b1111111111100101;
    assign weights1[45][407] = 16'b1111111111111010;
    assign weights1[45][408] = 16'b0000000000011010;
    assign weights1[45][409] = 16'b0000000000001000;
    assign weights1[45][410] = 16'b1111111111111001;
    assign weights1[45][411] = 16'b1111111111110000;
    assign weights1[45][412] = 16'b0000000000100001;
    assign weights1[45][413] = 16'b0000000000001011;
    assign weights1[45][414] = 16'b0000000000011001;
    assign weights1[45][415] = 16'b1111111111111100;
    assign weights1[45][416] = 16'b0000000000011001;
    assign weights1[45][417] = 16'b1111111111101011;
    assign weights1[45][418] = 16'b0000000000010100;
    assign weights1[45][419] = 16'b0000000000001000;
    assign weights1[45][420] = 16'b1111111111110100;
    assign weights1[45][421] = 16'b1111111111101111;
    assign weights1[45][422] = 16'b1111111111101010;
    assign weights1[45][423] = 16'b1111111111100000;
    assign weights1[45][424] = 16'b1111111111100101;
    assign weights1[45][425] = 16'b1111111111101101;
    assign weights1[45][426] = 16'b1111111111111100;
    assign weights1[45][427] = 16'b0000000000001001;
    assign weights1[45][428] = 16'b0000000000100110;
    assign weights1[45][429] = 16'b0000000000100001;
    assign weights1[45][430] = 16'b0000000000010111;
    assign weights1[45][431] = 16'b0000000000101110;
    assign weights1[45][432] = 16'b1111111111111101;
    assign weights1[45][433] = 16'b1111111111101010;
    assign weights1[45][434] = 16'b1111111111110110;
    assign weights1[45][435] = 16'b1111111111101000;
    assign weights1[45][436] = 16'b1111111111111100;
    assign weights1[45][437] = 16'b1111111111111011;
    assign weights1[45][438] = 16'b1111111111111110;
    assign weights1[45][439] = 16'b0000000000001101;
    assign weights1[45][440] = 16'b1111111111111111;
    assign weights1[45][441] = 16'b0000000000100100;
    assign weights1[45][442] = 16'b0000000000001111;
    assign weights1[45][443] = 16'b0000000000100011;
    assign weights1[45][444] = 16'b0000000000000111;
    assign weights1[45][445] = 16'b0000000000001110;
    assign weights1[45][446] = 16'b1111111111111101;
    assign weights1[45][447] = 16'b0000000000010011;
    assign weights1[45][448] = 16'b1111111111110101;
    assign weights1[45][449] = 16'b1111111111110000;
    assign weights1[45][450] = 16'b1111111111110001;
    assign weights1[45][451] = 16'b1111111111011110;
    assign weights1[45][452] = 16'b1111111111110010;
    assign weights1[45][453] = 16'b0000000000010101;
    assign weights1[45][454] = 16'b0000000000001111;
    assign weights1[45][455] = 16'b0000000000001110;
    assign weights1[45][456] = 16'b0000000000001110;
    assign weights1[45][457] = 16'b1111111111111100;
    assign weights1[45][458] = 16'b1111111111111010;
    assign weights1[45][459] = 16'b0000000000100010;
    assign weights1[45][460] = 16'b1111111111111000;
    assign weights1[45][461] = 16'b1111111111111000;
    assign weights1[45][462] = 16'b0000000000001001;
    assign weights1[45][463] = 16'b0000000000000100;
    assign weights1[45][464] = 16'b1111111111100010;
    assign weights1[45][465] = 16'b1111111111111000;
    assign weights1[45][466] = 16'b0000000000000010;
    assign weights1[45][467] = 16'b0000000000000101;
    assign weights1[45][468] = 16'b0000000000001101;
    assign weights1[45][469] = 16'b0000000000001010;
    assign weights1[45][470] = 16'b0000000000000100;
    assign weights1[45][471] = 16'b1111111111111010;
    assign weights1[45][472] = 16'b1111111111110000;
    assign weights1[45][473] = 16'b0000000000000100;
    assign weights1[45][474] = 16'b0000000000001011;
    assign weights1[45][475] = 16'b0000000000010000;
    assign weights1[45][476] = 16'b1111111111110111;
    assign weights1[45][477] = 16'b1111111111110001;
    assign weights1[45][478] = 16'b1111111111101110;
    assign weights1[45][479] = 16'b1111111111100011;
    assign weights1[45][480] = 16'b1111111111110111;
    assign weights1[45][481] = 16'b0000000000010001;
    assign weights1[45][482] = 16'b0000000000000101;
    assign weights1[45][483] = 16'b0000000000001001;
    assign weights1[45][484] = 16'b0000000000001100;
    assign weights1[45][485] = 16'b0000000000000110;
    assign weights1[45][486] = 16'b1111111111111100;
    assign weights1[45][487] = 16'b0000000000011011;
    assign weights1[45][488] = 16'b0000000000001010;
    assign weights1[45][489] = 16'b0000000000000101;
    assign weights1[45][490] = 16'b0000000000000000;
    assign weights1[45][491] = 16'b1111111111100111;
    assign weights1[45][492] = 16'b1111111111111010;
    assign weights1[45][493] = 16'b0000000000001111;
    assign weights1[45][494] = 16'b1111111111111110;
    assign weights1[45][495] = 16'b0000000000001010;
    assign weights1[45][496] = 16'b0000000000000100;
    assign weights1[45][497] = 16'b1111111111111111;
    assign weights1[45][498] = 16'b0000000000010001;
    assign weights1[45][499] = 16'b0000000000000010;
    assign weights1[45][500] = 16'b0000000000000010;
    assign weights1[45][501] = 16'b0000000000000111;
    assign weights1[45][502] = 16'b0000000000000111;
    assign weights1[45][503] = 16'b0000000000001100;
    assign weights1[45][504] = 16'b1111111111111101;
    assign weights1[45][505] = 16'b1111111111110001;
    assign weights1[45][506] = 16'b1111111111101110;
    assign weights1[45][507] = 16'b1111111111101010;
    assign weights1[45][508] = 16'b1111111111111101;
    assign weights1[45][509] = 16'b1111111111111001;
    assign weights1[45][510] = 16'b1111111111110100;
    assign weights1[45][511] = 16'b1111111111111110;
    assign weights1[45][512] = 16'b0000000000011001;
    assign weights1[45][513] = 16'b0000000000001011;
    assign weights1[45][514] = 16'b1111111111111111;
    assign weights1[45][515] = 16'b0000000000000010;
    assign weights1[45][516] = 16'b1111111111111100;
    assign weights1[45][517] = 16'b1111111111111010;
    assign weights1[45][518] = 16'b0000000000000100;
    assign weights1[45][519] = 16'b0000000000001010;
    assign weights1[45][520] = 16'b1111111111101111;
    assign weights1[45][521] = 16'b1111111111111000;
    assign weights1[45][522] = 16'b1111111111110100;
    assign weights1[45][523] = 16'b1111111111011100;
    assign weights1[45][524] = 16'b1111111111100111;
    assign weights1[45][525] = 16'b1111111111001101;
    assign weights1[45][526] = 16'b0000000000000100;
    assign weights1[45][527] = 16'b1111111111101010;
    assign weights1[45][528] = 16'b0000000000000010;
    assign weights1[45][529] = 16'b0000000000000001;
    assign weights1[45][530] = 16'b0000000000000110;
    assign weights1[45][531] = 16'b1111111111110101;
    assign weights1[45][532] = 16'b1111111111111111;
    assign weights1[45][533] = 16'b1111111111110100;
    assign weights1[45][534] = 16'b1111111111100111;
    assign weights1[45][535] = 16'b1111111111101000;
    assign weights1[45][536] = 16'b1111111111110001;
    assign weights1[45][537] = 16'b0000000000000011;
    assign weights1[45][538] = 16'b1111111111101011;
    assign weights1[45][539] = 16'b1111111111111011;
    assign weights1[45][540] = 16'b1111111111111110;
    assign weights1[45][541] = 16'b0000000000001000;
    assign weights1[45][542] = 16'b0000000000010001;
    assign weights1[45][543] = 16'b0000000000100000;
    assign weights1[45][544] = 16'b0000000000011000;
    assign weights1[45][545] = 16'b0000000000001110;
    assign weights1[45][546] = 16'b1111111111111100;
    assign weights1[45][547] = 16'b0000000000000001;
    assign weights1[45][548] = 16'b1111111111110001;
    assign weights1[45][549] = 16'b1111111111101000;
    assign weights1[45][550] = 16'b0000000000010101;
    assign weights1[45][551] = 16'b0000000000000110;
    assign weights1[45][552] = 16'b1111111111111101;
    assign weights1[45][553] = 16'b0000000000000101;
    assign weights1[45][554] = 16'b1111111111011100;
    assign weights1[45][555] = 16'b1111111111110110;
    assign weights1[45][556] = 16'b1111111111111100;
    assign weights1[45][557] = 16'b1111111111110010;
    assign weights1[45][558] = 16'b1111111111111001;
    assign weights1[45][559] = 16'b1111111111110111;
    assign weights1[45][560] = 16'b1111111111111010;
    assign weights1[45][561] = 16'b1111111111111001;
    assign weights1[45][562] = 16'b1111111111101000;
    assign weights1[45][563] = 16'b1111111111101010;
    assign weights1[45][564] = 16'b1111111111111110;
    assign weights1[45][565] = 16'b0000000000001001;
    assign weights1[45][566] = 16'b0000000000000111;
    assign weights1[45][567] = 16'b1111111111110001;
    assign weights1[45][568] = 16'b0000000000000101;
    assign weights1[45][569] = 16'b0000000000001001;
    assign weights1[45][570] = 16'b0000000000010111;
    assign weights1[45][571] = 16'b0000000000010001;
    assign weights1[45][572] = 16'b0000000000011111;
    assign weights1[45][573] = 16'b0000000000010100;
    assign weights1[45][574] = 16'b1111111111111101;
    assign weights1[45][575] = 16'b0000000000001010;
    assign weights1[45][576] = 16'b1111111111110011;
    assign weights1[45][577] = 16'b1111111111110111;
    assign weights1[45][578] = 16'b1111111111110010;
    assign weights1[45][579] = 16'b1111111111110111;
    assign weights1[45][580] = 16'b0000000000000001;
    assign weights1[45][581] = 16'b0000000000000100;
    assign weights1[45][582] = 16'b1111111111101101;
    assign weights1[45][583] = 16'b1111111111101011;
    assign weights1[45][584] = 16'b1111111111101111;
    assign weights1[45][585] = 16'b1111111111101100;
    assign weights1[45][586] = 16'b1111111111110011;
    assign weights1[45][587] = 16'b1111111111110001;
    assign weights1[45][588] = 16'b1111111111111011;
    assign weights1[45][589] = 16'b1111111111111000;
    assign weights1[45][590] = 16'b1111111111101101;
    assign weights1[45][591] = 16'b1111111111011111;
    assign weights1[45][592] = 16'b1111111111101001;
    assign weights1[45][593] = 16'b0000000000000010;
    assign weights1[45][594] = 16'b1111111111110111;
    assign weights1[45][595] = 16'b0000000000001001;
    assign weights1[45][596] = 16'b0000000000000001;
    assign weights1[45][597] = 16'b0000000000000110;
    assign weights1[45][598] = 16'b0000000000001110;
    assign weights1[45][599] = 16'b0000000000011001;
    assign weights1[45][600] = 16'b0000000000011011;
    assign weights1[45][601] = 16'b0000000000010011;
    assign weights1[45][602] = 16'b0000000000000111;
    assign weights1[45][603] = 16'b0000000000010110;
    assign weights1[45][604] = 16'b1111111111110011;
    assign weights1[45][605] = 16'b1111111111110110;
    assign weights1[45][606] = 16'b1111111111111111;
    assign weights1[45][607] = 16'b1111111111100100;
    assign weights1[45][608] = 16'b0000000000001100;
    assign weights1[45][609] = 16'b1111111111101010;
    assign weights1[45][610] = 16'b1111111111100111;
    assign weights1[45][611] = 16'b0000000000000100;
    assign weights1[45][612] = 16'b1111111111110100;
    assign weights1[45][613] = 16'b1111111111110110;
    assign weights1[45][614] = 16'b1111111111111000;
    assign weights1[45][615] = 16'b1111111111101110;
    assign weights1[45][616] = 16'b1111111111111000;
    assign weights1[45][617] = 16'b1111111111110110;
    assign weights1[45][618] = 16'b1111111111110010;
    assign weights1[45][619] = 16'b1111111111100101;
    assign weights1[45][620] = 16'b1111111111011111;
    assign weights1[45][621] = 16'b1111111111110011;
    assign weights1[45][622] = 16'b1111111111110011;
    assign weights1[45][623] = 16'b0000000000001100;
    assign weights1[45][624] = 16'b1111111111110001;
    assign weights1[45][625] = 16'b0000000000010011;
    assign weights1[45][626] = 16'b0000000000000100;
    assign weights1[45][627] = 16'b0000000000010000;
    assign weights1[45][628] = 16'b0000000000010100;
    assign weights1[45][629] = 16'b0000000000001010;
    assign weights1[45][630] = 16'b0000000000001000;
    assign weights1[45][631] = 16'b0000000000001010;
    assign weights1[45][632] = 16'b0000000000000001;
    assign weights1[45][633] = 16'b1111111111110000;
    assign weights1[45][634] = 16'b0000000000001100;
    assign weights1[45][635] = 16'b0000000000000111;
    assign weights1[45][636] = 16'b1111111111111010;
    assign weights1[45][637] = 16'b1111111111101101;
    assign weights1[45][638] = 16'b1111111111110110;
    assign weights1[45][639] = 16'b1111111111110000;
    assign weights1[45][640] = 16'b1111111111101111;
    assign weights1[45][641] = 16'b1111111111101111;
    assign weights1[45][642] = 16'b1111111111111000;
    assign weights1[45][643] = 16'b1111111111110101;
    assign weights1[45][644] = 16'b1111111111111101;
    assign weights1[45][645] = 16'b1111111111110111;
    assign weights1[45][646] = 16'b1111111111110000;
    assign weights1[45][647] = 16'b1111111111110111;
    assign weights1[45][648] = 16'b1111111111101101;
    assign weights1[45][649] = 16'b1111111111110001;
    assign weights1[45][650] = 16'b1111111111110010;
    assign weights1[45][651] = 16'b1111111111110010;
    assign weights1[45][652] = 16'b0000000000011111;
    assign weights1[45][653] = 16'b0000000000000100;
    assign weights1[45][654] = 16'b0000000000000111;
    assign weights1[45][655] = 16'b0000000000101000;
    assign weights1[45][656] = 16'b0000000000010110;
    assign weights1[45][657] = 16'b0000000000011011;
    assign weights1[45][658] = 16'b0000000000000100;
    assign weights1[45][659] = 16'b0000000000101011;
    assign weights1[45][660] = 16'b0000000000010000;
    assign weights1[45][661] = 16'b0000000000000000;
    assign weights1[45][662] = 16'b0000000000001010;
    assign weights1[45][663] = 16'b0000000000100000;
    assign weights1[45][664] = 16'b0000000000000001;
    assign weights1[45][665] = 16'b1111111111111010;
    assign weights1[45][666] = 16'b1111111111101111;
    assign weights1[45][667] = 16'b1111111111110110;
    assign weights1[45][668] = 16'b1111111111101001;
    assign weights1[45][669] = 16'b1111111111111001;
    assign weights1[45][670] = 16'b1111111111111001;
    assign weights1[45][671] = 16'b1111111111110101;
    assign weights1[45][672] = 16'b0000000000000000;
    assign weights1[45][673] = 16'b0000000000000001;
    assign weights1[45][674] = 16'b1111111111111001;
    assign weights1[45][675] = 16'b1111111111110010;
    assign weights1[45][676] = 16'b1111111111110101;
    assign weights1[45][677] = 16'b1111111111100110;
    assign weights1[45][678] = 16'b1111111111101000;
    assign weights1[45][679] = 16'b1111111111110110;
    assign weights1[45][680] = 16'b1111111111110001;
    assign weights1[45][681] = 16'b0000000000010100;
    assign weights1[45][682] = 16'b0000000000010101;
    assign weights1[45][683] = 16'b0000000000010011;
    assign weights1[45][684] = 16'b0000000000011010;
    assign weights1[45][685] = 16'b0000000000011010;
    assign weights1[45][686] = 16'b0000000000010000;
    assign weights1[45][687] = 16'b0000000000100011;
    assign weights1[45][688] = 16'b0000000000011100;
    assign weights1[45][689] = 16'b1111111111110001;
    assign weights1[45][690] = 16'b1111111111101010;
    assign weights1[45][691] = 16'b1111111111110010;
    assign weights1[45][692] = 16'b1111111111101001;
    assign weights1[45][693] = 16'b1111111111110111;
    assign weights1[45][694] = 16'b0000000000000110;
    assign weights1[45][695] = 16'b1111111111110111;
    assign weights1[45][696] = 16'b1111111111110101;
    assign weights1[45][697] = 16'b1111111111110101;
    assign weights1[45][698] = 16'b1111111111110111;
    assign weights1[45][699] = 16'b1111111111110100;
    assign weights1[45][700] = 16'b0000000000000000;
    assign weights1[45][701] = 16'b1111111111111111;
    assign weights1[45][702] = 16'b1111111111111100;
    assign weights1[45][703] = 16'b1111111111110101;
    assign weights1[45][704] = 16'b1111111111110001;
    assign weights1[45][705] = 16'b1111111111010111;
    assign weights1[45][706] = 16'b1111111111010111;
    assign weights1[45][707] = 16'b1111111111001110;
    assign weights1[45][708] = 16'b1111111111101110;
    assign weights1[45][709] = 16'b1111111111100010;
    assign weights1[45][710] = 16'b1111111111110001;
    assign weights1[45][711] = 16'b1111111111110010;
    assign weights1[45][712] = 16'b1111111111111010;
    assign weights1[45][713] = 16'b1111111111101101;
    assign weights1[45][714] = 16'b0000000000000000;
    assign weights1[45][715] = 16'b1111111111111101;
    assign weights1[45][716] = 16'b1111111111111001;
    assign weights1[45][717] = 16'b0000000000010010;
    assign weights1[45][718] = 16'b1111111111111101;
    assign weights1[45][719] = 16'b1111111111110101;
    assign weights1[45][720] = 16'b1111111111110101;
    assign weights1[45][721] = 16'b1111111111110011;
    assign weights1[45][722] = 16'b1111111111111010;
    assign weights1[45][723] = 16'b1111111111111101;
    assign weights1[45][724] = 16'b1111111111110001;
    assign weights1[45][725] = 16'b1111111111110110;
    assign weights1[45][726] = 16'b1111111111110100;
    assign weights1[45][727] = 16'b1111111111110110;
    assign weights1[45][728] = 16'b0000000000000000;
    assign weights1[45][729] = 16'b0000000000000001;
    assign weights1[45][730] = 16'b1111111111111100;
    assign weights1[45][731] = 16'b1111111111110101;
    assign weights1[45][732] = 16'b1111111111110001;
    assign weights1[45][733] = 16'b1111111111101110;
    assign weights1[45][734] = 16'b1111111111010011;
    assign weights1[45][735] = 16'b1111111111001111;
    assign weights1[45][736] = 16'b1111111111010001;
    assign weights1[45][737] = 16'b1111111111010111;
    assign weights1[45][738] = 16'b1111111111011011;
    assign weights1[45][739] = 16'b1111111111101011;
    assign weights1[45][740] = 16'b1111111111110001;
    assign weights1[45][741] = 16'b1111111111101011;
    assign weights1[45][742] = 16'b1111111111101011;
    assign weights1[45][743] = 16'b1111111111101001;
    assign weights1[45][744] = 16'b1111111111100110;
    assign weights1[45][745] = 16'b1111111111100100;
    assign weights1[45][746] = 16'b1111111111111110;
    assign weights1[45][747] = 16'b1111111111110000;
    assign weights1[45][748] = 16'b1111111111110000;
    assign weights1[45][749] = 16'b1111111111101010;
    assign weights1[45][750] = 16'b1111111111110001;
    assign weights1[45][751] = 16'b1111111111110011;
    assign weights1[45][752] = 16'b1111111111110011;
    assign weights1[45][753] = 16'b1111111111111001;
    assign weights1[45][754] = 16'b1111111111110111;
    assign weights1[45][755] = 16'b1111111111111010;
    assign weights1[45][756] = 16'b1111111111111111;
    assign weights1[45][757] = 16'b1111111111111110;
    assign weights1[45][758] = 16'b1111111111111000;
    assign weights1[45][759] = 16'b1111111111111001;
    assign weights1[45][760] = 16'b1111111111101101;
    assign weights1[45][761] = 16'b1111111111100101;
    assign weights1[45][762] = 16'b1111111111100111;
    assign weights1[45][763] = 16'b1111111111011100;
    assign weights1[45][764] = 16'b1111111111001111;
    assign weights1[45][765] = 16'b1111111111001011;
    assign weights1[45][766] = 16'b1111111111011011;
    assign weights1[45][767] = 16'b1111111111000101;
    assign weights1[45][768] = 16'b1111111111001000;
    assign weights1[45][769] = 16'b1111111111000011;
    assign weights1[45][770] = 16'b1111111110111100;
    assign weights1[45][771] = 16'b1111111111001101;
    assign weights1[45][772] = 16'b1111111111001011;
    assign weights1[45][773] = 16'b1111111111100000;
    assign weights1[45][774] = 16'b1111111111100000;
    assign weights1[45][775] = 16'b1111111111011110;
    assign weights1[45][776] = 16'b1111111111101011;
    assign weights1[45][777] = 16'b1111111111100110;
    assign weights1[45][778] = 16'b1111111111110001;
    assign weights1[45][779] = 16'b1111111111110011;
    assign weights1[45][780] = 16'b1111111111110110;
    assign weights1[45][781] = 16'b1111111111111101;
    assign weights1[45][782] = 16'b1111111111111100;
    assign weights1[45][783] = 16'b1111111111111101;
    assign weights1[46][0] = 16'b0000000000000000;
    assign weights1[46][1] = 16'b0000000000000000;
    assign weights1[46][2] = 16'b0000000000000000;
    assign weights1[46][3] = 16'b0000000000000000;
    assign weights1[46][4] = 16'b0000000000000000;
    assign weights1[46][5] = 16'b0000000000000001;
    assign weights1[46][6] = 16'b1111111111111111;
    assign weights1[46][7] = 16'b1111111111111000;
    assign weights1[46][8] = 16'b1111111111110100;
    assign weights1[46][9] = 16'b1111111111101101;
    assign weights1[46][10] = 16'b1111111111101101;
    assign weights1[46][11] = 16'b1111111111100111;
    assign weights1[46][12] = 16'b1111111111101000;
    assign weights1[46][13] = 16'b1111111111100110;
    assign weights1[46][14] = 16'b1111111111100011;
    assign weights1[46][15] = 16'b1111111111100000;
    assign weights1[46][16] = 16'b1111111111010110;
    assign weights1[46][17] = 16'b1111111111011101;
    assign weights1[46][18] = 16'b1111111111010101;
    assign weights1[46][19] = 16'b1111111111101000;
    assign weights1[46][20] = 16'b1111111111110011;
    assign weights1[46][21] = 16'b1111111111111110;
    assign weights1[46][22] = 16'b0000000000001010;
    assign weights1[46][23] = 16'b0000000000001000;
    assign weights1[46][24] = 16'b0000000000000001;
    assign weights1[46][25] = 16'b0000000000000110;
    assign weights1[46][26] = 16'b0000000000000111;
    assign weights1[46][27] = 16'b0000000000000000;
    assign weights1[46][28] = 16'b0000000000000000;
    assign weights1[46][29] = 16'b0000000000000000;
    assign weights1[46][30] = 16'b1111111111111110;
    assign weights1[46][31] = 16'b1111111111111110;
    assign weights1[46][32] = 16'b1111111111111100;
    assign weights1[46][33] = 16'b1111111111111110;
    assign weights1[46][34] = 16'b1111111111111011;
    assign weights1[46][35] = 16'b1111111111111010;
    assign weights1[46][36] = 16'b1111111111110100;
    assign weights1[46][37] = 16'b1111111111111110;
    assign weights1[46][38] = 16'b1111111111110101;
    assign weights1[46][39] = 16'b1111111111011101;
    assign weights1[46][40] = 16'b1111111111011110;
    assign weights1[46][41] = 16'b1111111111100100;
    assign weights1[46][42] = 16'b1111111111100010;
    assign weights1[46][43] = 16'b1111111111010001;
    assign weights1[46][44] = 16'b1111111111100011;
    assign weights1[46][45] = 16'b1111111111011000;
    assign weights1[46][46] = 16'b1111111111011110;
    assign weights1[46][47] = 16'b1111111111110011;
    assign weights1[46][48] = 16'b1111111111111001;
    assign weights1[46][49] = 16'b1111111111101111;
    assign weights1[46][50] = 16'b0000000000000011;
    assign weights1[46][51] = 16'b0000000000001000;
    assign weights1[46][52] = 16'b0000000000000010;
    assign weights1[46][53] = 16'b0000000000000101;
    assign weights1[46][54] = 16'b0000000000000101;
    assign weights1[46][55] = 16'b1111111111111110;
    assign weights1[46][56] = 16'b0000000000000000;
    assign weights1[46][57] = 16'b0000000000000000;
    assign weights1[46][58] = 16'b1111111111111111;
    assign weights1[46][59] = 16'b1111111111111110;
    assign weights1[46][60] = 16'b1111111111111011;
    assign weights1[46][61] = 16'b1111111111111001;
    assign weights1[46][62] = 16'b1111111111111001;
    assign weights1[46][63] = 16'b1111111111111110;
    assign weights1[46][64] = 16'b0000000000000010;
    assign weights1[46][65] = 16'b1111111111110101;
    assign weights1[46][66] = 16'b1111111111110100;
    assign weights1[46][67] = 16'b1111111111110111;
    assign weights1[46][68] = 16'b1111111111100110;
    assign weights1[46][69] = 16'b1111111111101100;
    assign weights1[46][70] = 16'b1111111111100011;
    assign weights1[46][71] = 16'b1111111111111001;
    assign weights1[46][72] = 16'b1111111111111000;
    assign weights1[46][73] = 16'b1111111111100010;
    assign weights1[46][74] = 16'b0000000000000101;
    assign weights1[46][75] = 16'b1111111111101110;
    assign weights1[46][76] = 16'b1111111111110100;
    assign weights1[46][77] = 16'b1111111111111101;
    assign weights1[46][78] = 16'b0000000000010000;
    assign weights1[46][79] = 16'b0000000000000100;
    assign weights1[46][80] = 16'b0000000000000000;
    assign weights1[46][81] = 16'b0000000000011011;
    assign weights1[46][82] = 16'b0000000000010110;
    assign weights1[46][83] = 16'b0000000000001110;
    assign weights1[46][84] = 16'b1111111111111110;
    assign weights1[46][85] = 16'b1111111111111110;
    assign weights1[46][86] = 16'b1111111111111101;
    assign weights1[46][87] = 16'b1111111111111010;
    assign weights1[46][88] = 16'b1111111111111001;
    assign weights1[46][89] = 16'b1111111111111111;
    assign weights1[46][90] = 16'b1111111111110010;
    assign weights1[46][91] = 16'b0000000000000001;
    assign weights1[46][92] = 16'b1111111111111010;
    assign weights1[46][93] = 16'b0000000000000100;
    assign weights1[46][94] = 16'b1111111111101001;
    assign weights1[46][95] = 16'b0000000000000100;
    assign weights1[46][96] = 16'b1111111111101100;
    assign weights1[46][97] = 16'b1111111111111001;
    assign weights1[46][98] = 16'b1111111111111101;
    assign weights1[46][99] = 16'b0000000000000100;
    assign weights1[46][100] = 16'b0000000000000100;
    assign weights1[46][101] = 16'b1111111111111001;
    assign weights1[46][102] = 16'b0000000000011000;
    assign weights1[46][103] = 16'b0000000000101001;
    assign weights1[46][104] = 16'b0000000000011101;
    assign weights1[46][105] = 16'b0000000000011100;
    assign weights1[46][106] = 16'b0000000000010100;
    assign weights1[46][107] = 16'b0000000000010100;
    assign weights1[46][108] = 16'b1111111111111101;
    assign weights1[46][109] = 16'b0000000000010110;
    assign weights1[46][110] = 16'b0000000000101000;
    assign weights1[46][111] = 16'b0000000000011011;
    assign weights1[46][112] = 16'b1111111111111110;
    assign weights1[46][113] = 16'b1111111111111110;
    assign weights1[46][114] = 16'b0000000000000001;
    assign weights1[46][115] = 16'b1111111111111111;
    assign weights1[46][116] = 16'b1111111111101111;
    assign weights1[46][117] = 16'b1111111111110011;
    assign weights1[46][118] = 16'b1111111111110111;
    assign weights1[46][119] = 16'b1111111111111011;
    assign weights1[46][120] = 16'b1111111111111000;
    assign weights1[46][121] = 16'b1111111111110101;
    assign weights1[46][122] = 16'b1111111111101110;
    assign weights1[46][123] = 16'b1111111111111110;
    assign weights1[46][124] = 16'b1111111111110010;
    assign weights1[46][125] = 16'b1111111111110001;
    assign weights1[46][126] = 16'b1111111111111101;
    assign weights1[46][127] = 16'b0000000000000111;
    assign weights1[46][128] = 16'b1111111111111100;
    assign weights1[46][129] = 16'b0000000000010001;
    assign weights1[46][130] = 16'b0000000000011100;
    assign weights1[46][131] = 16'b0000000000011111;
    assign weights1[46][132] = 16'b1111111111110110;
    assign weights1[46][133] = 16'b0000000000010100;
    assign weights1[46][134] = 16'b0000000000010011;
    assign weights1[46][135] = 16'b0000000000011111;
    assign weights1[46][136] = 16'b0000000000100110;
    assign weights1[46][137] = 16'b0000000000010010;
    assign weights1[46][138] = 16'b0000000000011011;
    assign weights1[46][139] = 16'b0000000000100100;
    assign weights1[46][140] = 16'b1111111111111001;
    assign weights1[46][141] = 16'b1111111111111011;
    assign weights1[46][142] = 16'b1111111111111000;
    assign weights1[46][143] = 16'b1111111111110110;
    assign weights1[46][144] = 16'b1111111111101111;
    assign weights1[46][145] = 16'b1111111111011110;
    assign weights1[46][146] = 16'b1111111111111101;
    assign weights1[46][147] = 16'b1111111111100000;
    assign weights1[46][148] = 16'b0000000000001000;
    assign weights1[46][149] = 16'b1111111111111010;
    assign weights1[46][150] = 16'b0000000000010010;
    assign weights1[46][151] = 16'b0000000000000001;
    assign weights1[46][152] = 16'b1111111111111100;
    assign weights1[46][153] = 16'b0000000000001001;
    assign weights1[46][154] = 16'b0000000000001000;
    assign weights1[46][155] = 16'b0000000000000100;
    assign weights1[46][156] = 16'b0000000000100011;
    assign weights1[46][157] = 16'b0000000000001000;
    assign weights1[46][158] = 16'b0000000000011011;
    assign weights1[46][159] = 16'b0000000000001000;
    assign weights1[46][160] = 16'b0000000000011010;
    assign weights1[46][161] = 16'b0000000000100001;
    assign weights1[46][162] = 16'b0000000000101001;
    assign weights1[46][163] = 16'b0000000000110110;
    assign weights1[46][164] = 16'b0000000000101001;
    assign weights1[46][165] = 16'b0000000000100010;
    assign weights1[46][166] = 16'b0000000000010111;
    assign weights1[46][167] = 16'b0000000000101110;
    assign weights1[46][168] = 16'b1111111111111010;
    assign weights1[46][169] = 16'b1111111111110101;
    assign weights1[46][170] = 16'b1111111111111000;
    assign weights1[46][171] = 16'b1111111111111010;
    assign weights1[46][172] = 16'b1111111111100010;
    assign weights1[46][173] = 16'b1111111111101010;
    assign weights1[46][174] = 16'b1111111111101111;
    assign weights1[46][175] = 16'b0000000000010110;
    assign weights1[46][176] = 16'b1111111111110111;
    assign weights1[46][177] = 16'b0000000000000011;
    assign weights1[46][178] = 16'b1111111111110101;
    assign weights1[46][179] = 16'b0000000000000100;
    assign weights1[46][180] = 16'b0000000000001011;
    assign weights1[46][181] = 16'b1111111111111111;
    assign weights1[46][182] = 16'b0000000000010000;
    assign weights1[46][183] = 16'b0000000000000100;
    assign weights1[46][184] = 16'b1111111111110111;
    assign weights1[46][185] = 16'b0000000000000101;
    assign weights1[46][186] = 16'b0000000000000110;
    assign weights1[46][187] = 16'b0000000000100110;
    assign weights1[46][188] = 16'b0000000000100111;
    assign weights1[46][189] = 16'b0000000000011100;
    assign weights1[46][190] = 16'b0000000000011000;
    assign weights1[46][191] = 16'b0000000000101100;
    assign weights1[46][192] = 16'b0000000001011110;
    assign weights1[46][193] = 16'b0000000000101110;
    assign weights1[46][194] = 16'b0000000000101110;
    assign weights1[46][195] = 16'b0000000000100100;
    assign weights1[46][196] = 16'b1111111111111100;
    assign weights1[46][197] = 16'b1111111111110111;
    assign weights1[46][198] = 16'b1111111111101000;
    assign weights1[46][199] = 16'b0000000000000010;
    assign weights1[46][200] = 16'b1111111111110011;
    assign weights1[46][201] = 16'b1111111111111110;
    assign weights1[46][202] = 16'b0000000000000100;
    assign weights1[46][203] = 16'b0000000000001101;
    assign weights1[46][204] = 16'b1111111111110011;
    assign weights1[46][205] = 16'b1111111111110101;
    assign weights1[46][206] = 16'b0000000000001100;
    assign weights1[46][207] = 16'b1111111111111110;
    assign weights1[46][208] = 16'b0000000000001100;
    assign weights1[46][209] = 16'b0000000000000100;
    assign weights1[46][210] = 16'b0000000000011101;
    assign weights1[46][211] = 16'b0000000000010011;
    assign weights1[46][212] = 16'b0000000000101000;
    assign weights1[46][213] = 16'b0000000000110010;
    assign weights1[46][214] = 16'b0000000000110111;
    assign weights1[46][215] = 16'b0000000000111111;
    assign weights1[46][216] = 16'b0000000001010101;
    assign weights1[46][217] = 16'b0000000001001000;
    assign weights1[46][218] = 16'b0000000001000011;
    assign weights1[46][219] = 16'b0000000001101010;
    assign weights1[46][220] = 16'b0000000001010011;
    assign weights1[46][221] = 16'b0000000000100101;
    assign weights1[46][222] = 16'b0000000000011000;
    assign weights1[46][223] = 16'b1111111111111011;
    assign weights1[46][224] = 16'b1111111111111101;
    assign weights1[46][225] = 16'b1111111111110000;
    assign weights1[46][226] = 16'b1111111111110011;
    assign weights1[46][227] = 16'b0000000000000101;
    assign weights1[46][228] = 16'b1111111111100010;
    assign weights1[46][229] = 16'b1111111111111010;
    assign weights1[46][230] = 16'b1111111111110111;
    assign weights1[46][231] = 16'b1111111111111100;
    assign weights1[46][232] = 16'b1111111111110111;
    assign weights1[46][233] = 16'b0000000000000001;
    assign weights1[46][234] = 16'b1111111111111110;
    assign weights1[46][235] = 16'b0000000000010000;
    assign weights1[46][236] = 16'b0000000000001111;
    assign weights1[46][237] = 16'b0000000000010100;
    assign weights1[46][238] = 16'b0000000000011000;
    assign weights1[46][239] = 16'b0000000000001111;
    assign weights1[46][240] = 16'b0000000000101010;
    assign weights1[46][241] = 16'b0000000000101000;
    assign weights1[46][242] = 16'b0000000000100110;
    assign weights1[46][243] = 16'b0000000000110000;
    assign weights1[46][244] = 16'b0000000001000100;
    assign weights1[46][245] = 16'b0000000000110000;
    assign weights1[46][246] = 16'b0000000000010111;
    assign weights1[46][247] = 16'b0000000001000010;
    assign weights1[46][248] = 16'b0000000000010101;
    assign weights1[46][249] = 16'b1111111111001011;
    assign weights1[46][250] = 16'b1111111111001000;
    assign weights1[46][251] = 16'b1111111111000101;
    assign weights1[46][252] = 16'b1111111111110100;
    assign weights1[46][253] = 16'b1111111111111001;
    assign weights1[46][254] = 16'b0000000000001100;
    assign weights1[46][255] = 16'b1111111111111100;
    assign weights1[46][256] = 16'b1111111111111011;
    assign weights1[46][257] = 16'b1111111111101000;
    assign weights1[46][258] = 16'b1111111111111100;
    assign weights1[46][259] = 16'b1111111111110100;
    assign weights1[46][260] = 16'b0000000000000001;
    assign weights1[46][261] = 16'b1111111111111101;
    assign weights1[46][262] = 16'b0000000000000011;
    assign weights1[46][263] = 16'b1111111111110100;
    assign weights1[46][264] = 16'b1111111111110110;
    assign weights1[46][265] = 16'b1111111111101111;
    assign weights1[46][266] = 16'b1111111111011111;
    assign weights1[46][267] = 16'b1111111111010011;
    assign weights1[46][268] = 16'b1111111110111010;
    assign weights1[46][269] = 16'b1111111111000001;
    assign weights1[46][270] = 16'b1111111110101000;
    assign weights1[46][271] = 16'b1111111110100000;
    assign weights1[46][272] = 16'b1111111110000010;
    assign weights1[46][273] = 16'b1111111110000111;
    assign weights1[46][274] = 16'b1111111110010000;
    assign weights1[46][275] = 16'b1111111101101010;
    assign weights1[46][276] = 16'b1111111101110010;
    assign weights1[46][277] = 16'b1111111110101000;
    assign weights1[46][278] = 16'b1111111110100010;
    assign weights1[46][279] = 16'b1111111110100000;
    assign weights1[46][280] = 16'b1111111111110110;
    assign weights1[46][281] = 16'b1111111111110101;
    assign weights1[46][282] = 16'b0000000000000010;
    assign weights1[46][283] = 16'b1111111111111011;
    assign weights1[46][284] = 16'b1111111111111001;
    assign weights1[46][285] = 16'b1111111111101111;
    assign weights1[46][286] = 16'b1111111111111000;
    assign weights1[46][287] = 16'b0000000000000101;
    assign weights1[46][288] = 16'b1111111111101110;
    assign weights1[46][289] = 16'b1111111111111111;
    assign weights1[46][290] = 16'b1111111111110011;
    assign weights1[46][291] = 16'b1111111111110101;
    assign weights1[46][292] = 16'b1111111111001011;
    assign weights1[46][293] = 16'b1111111111001110;
    assign weights1[46][294] = 16'b1111111110110101;
    assign weights1[46][295] = 16'b1111111110100010;
    assign weights1[46][296] = 16'b1111111101110110;
    assign weights1[46][297] = 16'b1111111100011100;
    assign weights1[46][298] = 16'b1111111011101101;
    assign weights1[46][299] = 16'b1111111011001111;
    assign weights1[46][300] = 16'b1111111100000011;
    assign weights1[46][301] = 16'b1111111100100001;
    assign weights1[46][302] = 16'b1111111100110011;
    assign weights1[46][303] = 16'b1111111101010100;
    assign weights1[46][304] = 16'b1111111101001000;
    assign weights1[46][305] = 16'b1111111110000001;
    assign weights1[46][306] = 16'b1111111110011001;
    assign weights1[46][307] = 16'b1111111110010100;
    assign weights1[46][308] = 16'b1111111111111010;
    assign weights1[46][309] = 16'b0000000000000001;
    assign weights1[46][310] = 16'b1111111111111000;
    assign weights1[46][311] = 16'b1111111111110110;
    assign weights1[46][312] = 16'b0000000000001110;
    assign weights1[46][313] = 16'b0000000000000001;
    assign weights1[46][314] = 16'b0000000000001000;
    assign weights1[46][315] = 16'b0000000000001100;
    assign weights1[46][316] = 16'b1111111111101111;
    assign weights1[46][317] = 16'b1111111111101001;
    assign weights1[46][318] = 16'b1111111111110000;
    assign weights1[46][319] = 16'b1111111111101011;
    assign weights1[46][320] = 16'b1111111111110101;
    assign weights1[46][321] = 16'b1111111111011011;
    assign weights1[46][322] = 16'b1111111111110000;
    assign weights1[46][323] = 16'b1111111111110101;
    assign weights1[46][324] = 16'b1111111111101110;
    assign weights1[46][325] = 16'b1111111111101001;
    assign weights1[46][326] = 16'b1111111111000110;
    assign weights1[46][327] = 16'b1111111110000101;
    assign weights1[46][328] = 16'b1111111100110110;
    assign weights1[46][329] = 16'b1111111100100000;
    assign weights1[46][330] = 16'b1111111100110011;
    assign weights1[46][331] = 16'b1111111101000010;
    assign weights1[46][332] = 16'b1111111101010100;
    assign weights1[46][333] = 16'b1111111101111100;
    assign weights1[46][334] = 16'b1111111110101000;
    assign weights1[46][335] = 16'b1111111110011011;
    assign weights1[46][336] = 16'b0000000000000010;
    assign weights1[46][337] = 16'b1111111111111001;
    assign weights1[46][338] = 16'b1111111111111110;
    assign weights1[46][339] = 16'b0000000000000101;
    assign weights1[46][340] = 16'b1111111111110000;
    assign weights1[46][341] = 16'b0000000000000001;
    assign weights1[46][342] = 16'b1111111111101110;
    assign weights1[46][343] = 16'b1111111111110011;
    assign weights1[46][344] = 16'b0000000000010000;
    assign weights1[46][345] = 16'b1111111111110101;
    assign weights1[46][346] = 16'b1111111111110110;
    assign weights1[46][347] = 16'b1111111111111101;
    assign weights1[46][348] = 16'b0000000000000100;
    assign weights1[46][349] = 16'b0000000000000011;
    assign weights1[46][350] = 16'b0000000000000010;
    assign weights1[46][351] = 16'b1111111111111101;
    assign weights1[46][352] = 16'b0000000000010011;
    assign weights1[46][353] = 16'b0000000000010110;
    assign weights1[46][354] = 16'b0000000000010000;
    assign weights1[46][355] = 16'b1111111111111111;
    assign weights1[46][356] = 16'b1111111111100001;
    assign weights1[46][357] = 16'b1111111110110000;
    assign weights1[46][358] = 16'b1111111101111110;
    assign weights1[46][359] = 16'b1111111101111011;
    assign weights1[46][360] = 16'b1111111101101100;
    assign weights1[46][361] = 16'b1111111101111011;
    assign weights1[46][362] = 16'b1111111110011111;
    assign weights1[46][363] = 16'b1111111110010110;
    assign weights1[46][364] = 16'b1111111111111111;
    assign weights1[46][365] = 16'b0000000000000000;
    assign weights1[46][366] = 16'b0000000000001010;
    assign weights1[46][367] = 16'b1111111111111000;
    assign weights1[46][368] = 16'b0000000000000110;
    assign weights1[46][369] = 16'b1111111111110101;
    assign weights1[46][370] = 16'b0000000000010010;
    assign weights1[46][371] = 16'b1111111111111010;
    assign weights1[46][372] = 16'b1111111111101101;
    assign weights1[46][373] = 16'b1111111111110111;
    assign weights1[46][374] = 16'b0000000000000010;
    assign weights1[46][375] = 16'b0000000000000000;
    assign weights1[46][376] = 16'b0000000000001100;
    assign weights1[46][377] = 16'b0000000000000010;
    assign weights1[46][378] = 16'b1111111111111100;
    assign weights1[46][379] = 16'b0000000000000110;
    assign weights1[46][380] = 16'b1111111111110001;
    assign weights1[46][381] = 16'b0000000000010100;
    assign weights1[46][382] = 16'b1111111111111100;
    assign weights1[46][383] = 16'b0000000000001111;
    assign weights1[46][384] = 16'b0000000000010100;
    assign weights1[46][385] = 16'b0000000000000101;
    assign weights1[46][386] = 16'b0000000000010101;
    assign weights1[46][387] = 16'b1111111111010001;
    assign weights1[46][388] = 16'b1111111111011000;
    assign weights1[46][389] = 16'b1111111110111001;
    assign weights1[46][390] = 16'b1111111110100111;
    assign weights1[46][391] = 16'b1111111110100101;
    assign weights1[46][392] = 16'b1111111111110111;
    assign weights1[46][393] = 16'b0000000000000111;
    assign weights1[46][394] = 16'b0000000000010000;
    assign weights1[46][395] = 16'b0000000000000010;
    assign weights1[46][396] = 16'b0000000000010001;
    assign weights1[46][397] = 16'b1111111111101001;
    assign weights1[46][398] = 16'b0000000000011001;
    assign weights1[46][399] = 16'b0000000000010000;
    assign weights1[46][400] = 16'b0000000000010011;
    assign weights1[46][401] = 16'b1111111111111111;
    assign weights1[46][402] = 16'b0000000000000001;
    assign weights1[46][403] = 16'b0000000000001110;
    assign weights1[46][404] = 16'b1111111111111101;
    assign weights1[46][405] = 16'b0000000000001010;
    assign weights1[46][406] = 16'b1111111111111111;
    assign weights1[46][407] = 16'b0000000000001010;
    assign weights1[46][408] = 16'b0000000000001001;
    assign weights1[46][409] = 16'b1111111111111010;
    assign weights1[46][410] = 16'b0000000000010000;
    assign weights1[46][411] = 16'b0000000000010001;
    assign weights1[46][412] = 16'b0000000000100000;
    assign weights1[46][413] = 16'b0000000000010001;
    assign weights1[46][414] = 16'b0000000000011101;
    assign weights1[46][415] = 16'b0000000000100100;
    assign weights1[46][416] = 16'b0000000000100010;
    assign weights1[46][417] = 16'b1111111111110110;
    assign weights1[46][418] = 16'b1111111111100000;
    assign weights1[46][419] = 16'b1111111111010011;
    assign weights1[46][420] = 16'b1111111111111101;
    assign weights1[46][421] = 16'b0000000000001011;
    assign weights1[46][422] = 16'b0000000000000010;
    assign weights1[46][423] = 16'b0000000000000010;
    assign weights1[46][424] = 16'b0000000000010110;
    assign weights1[46][425] = 16'b0000000000001101;
    assign weights1[46][426] = 16'b0000000000000101;
    assign weights1[46][427] = 16'b1111111111110100;
    assign weights1[46][428] = 16'b0000000000010100;
    assign weights1[46][429] = 16'b1111111111111011;
    assign weights1[46][430] = 16'b0000000000001111;
    assign weights1[46][431] = 16'b0000000000000001;
    assign weights1[46][432] = 16'b1111111111110100;
    assign weights1[46][433] = 16'b1111111111111111;
    assign weights1[46][434] = 16'b1111111111101011;
    assign weights1[46][435] = 16'b0000000000001001;
    assign weights1[46][436] = 16'b0000000000000111;
    assign weights1[46][437] = 16'b0000000000000111;
    assign weights1[46][438] = 16'b0000000000001001;
    assign weights1[46][439] = 16'b0000000000000000;
    assign weights1[46][440] = 16'b0000000000011010;
    assign weights1[46][441] = 16'b0000000000010101;
    assign weights1[46][442] = 16'b0000000000000001;
    assign weights1[46][443] = 16'b0000000000101001;
    assign weights1[46][444] = 16'b0000000000011011;
    assign weights1[46][445] = 16'b0000000000000110;
    assign weights1[46][446] = 16'b0000000000000001;
    assign weights1[46][447] = 16'b1111111111110110;
    assign weights1[46][448] = 16'b1111111111111110;
    assign weights1[46][449] = 16'b0000000000010000;
    assign weights1[46][450] = 16'b0000000000001111;
    assign weights1[46][451] = 16'b1111111111111010;
    assign weights1[46][452] = 16'b0000000000000001;
    assign weights1[46][453] = 16'b1111111111111100;
    assign weights1[46][454] = 16'b1111111111111101;
    assign weights1[46][455] = 16'b0000000000001010;
    assign weights1[46][456] = 16'b1111111111111010;
    assign weights1[46][457] = 16'b0000000000001001;
    assign weights1[46][458] = 16'b0000000000000011;
    assign weights1[46][459] = 16'b0000000000000100;
    assign weights1[46][460] = 16'b1111111111111100;
    assign weights1[46][461] = 16'b0000000000000110;
    assign weights1[46][462] = 16'b0000000000001100;
    assign weights1[46][463] = 16'b0000000000000101;
    assign weights1[46][464] = 16'b1111111111111110;
    assign weights1[46][465] = 16'b0000000000010110;
    assign weights1[46][466] = 16'b0000000000000001;
    assign weights1[46][467] = 16'b0000000000000101;
    assign weights1[46][468] = 16'b1111111111111110;
    assign weights1[46][469] = 16'b0000000000001011;
    assign weights1[46][470] = 16'b0000000000100000;
    assign weights1[46][471] = 16'b0000000000001010;
    assign weights1[46][472] = 16'b0000000000010001;
    assign weights1[46][473] = 16'b1111111111111011;
    assign weights1[46][474] = 16'b0000000000000110;
    assign weights1[46][475] = 16'b0000000000000100;
    assign weights1[46][476] = 16'b0000000000000100;
    assign weights1[46][477] = 16'b1111111111111100;
    assign weights1[46][478] = 16'b1111111111111010;
    assign weights1[46][479] = 16'b1111111111111110;
    assign weights1[46][480] = 16'b1111111111110011;
    assign weights1[46][481] = 16'b0000000000001101;
    assign weights1[46][482] = 16'b1111111111111010;
    assign weights1[46][483] = 16'b0000000000000011;
    assign weights1[46][484] = 16'b0000000000010100;
    assign weights1[46][485] = 16'b1111111111110011;
    assign weights1[46][486] = 16'b0000000000000100;
    assign weights1[46][487] = 16'b0000000000000111;
    assign weights1[46][488] = 16'b1111111111111010;
    assign weights1[46][489] = 16'b0000000000000000;
    assign weights1[46][490] = 16'b1111111111110010;
    assign weights1[46][491] = 16'b1111111111111000;
    assign weights1[46][492] = 16'b1111111111111011;
    assign weights1[46][493] = 16'b1111111111111010;
    assign weights1[46][494] = 16'b0000000000010100;
    assign weights1[46][495] = 16'b0000000000000011;
    assign weights1[46][496] = 16'b0000000000001110;
    assign weights1[46][497] = 16'b1111111111101110;
    assign weights1[46][498] = 16'b1111111111111111;
    assign weights1[46][499] = 16'b0000000000000101;
    assign weights1[46][500] = 16'b0000000000010010;
    assign weights1[46][501] = 16'b1111111111111101;
    assign weights1[46][502] = 16'b0000000000010000;
    assign weights1[46][503] = 16'b1111111111110101;
    assign weights1[46][504] = 16'b1111111111111111;
    assign weights1[46][505] = 16'b1111111111110101;
    assign weights1[46][506] = 16'b1111111111111101;
    assign weights1[46][507] = 16'b0000000000010010;
    assign weights1[46][508] = 16'b0000000000000100;
    assign weights1[46][509] = 16'b1111111111111111;
    assign weights1[46][510] = 16'b0000000000000001;
    assign weights1[46][511] = 16'b0000000000000011;
    assign weights1[46][512] = 16'b1111111111110111;
    assign weights1[46][513] = 16'b0000000000000110;
    assign weights1[46][514] = 16'b0000000000000000;
    assign weights1[46][515] = 16'b1111111111111000;
    assign weights1[46][516] = 16'b0000000000001001;
    assign weights1[46][517] = 16'b0000000000001110;
    assign weights1[46][518] = 16'b1111111111110100;
    assign weights1[46][519] = 16'b0000000000000111;
    assign weights1[46][520] = 16'b0000000000001010;
    assign weights1[46][521] = 16'b1111111111111111;
    assign weights1[46][522] = 16'b1111111111111100;
    assign weights1[46][523] = 16'b0000000000011001;
    assign weights1[46][524] = 16'b0000000000000101;
    assign weights1[46][525] = 16'b1111111111111101;
    assign weights1[46][526] = 16'b0000000000000110;
    assign weights1[46][527] = 16'b0000000000001010;
    assign weights1[46][528] = 16'b1111111111111000;
    assign weights1[46][529] = 16'b0000000000000110;
    assign weights1[46][530] = 16'b0000000000000011;
    assign weights1[46][531] = 16'b1111111111111000;
    assign weights1[46][532] = 16'b1111111111111000;
    assign weights1[46][533] = 16'b0000000000000011;
    assign weights1[46][534] = 16'b0000000000000100;
    assign weights1[46][535] = 16'b1111111111110000;
    assign weights1[46][536] = 16'b0000000000000110;
    assign weights1[46][537] = 16'b0000000000001100;
    assign weights1[46][538] = 16'b1111111111111001;
    assign weights1[46][539] = 16'b1111111111101100;
    assign weights1[46][540] = 16'b0000000000010001;
    assign weights1[46][541] = 16'b0000000000000001;
    assign weights1[46][542] = 16'b0000000000000000;
    assign weights1[46][543] = 16'b1111111111110101;
    assign weights1[46][544] = 16'b0000000000011100;
    assign weights1[46][545] = 16'b1111111111110110;
    assign weights1[46][546] = 16'b0000000000010010;
    assign weights1[46][547] = 16'b0000000000000100;
    assign weights1[46][548] = 16'b0000000000000011;
    assign weights1[46][549] = 16'b0000000000001000;
    assign weights1[46][550] = 16'b0000000000000110;
    assign weights1[46][551] = 16'b0000000000000000;
    assign weights1[46][552] = 16'b1111111111111110;
    assign weights1[46][553] = 16'b0000000000000110;
    assign weights1[46][554] = 16'b0000000000010011;
    assign weights1[46][555] = 16'b1111111111101111;
    assign weights1[46][556] = 16'b0000000000011010;
    assign weights1[46][557] = 16'b0000000000000110;
    assign weights1[46][558] = 16'b0000000000001011;
    assign weights1[46][559] = 16'b0000000000010000;
    assign weights1[46][560] = 16'b1111111111111111;
    assign weights1[46][561] = 16'b1111111111111011;
    assign weights1[46][562] = 16'b1111111111111110;
    assign weights1[46][563] = 16'b1111111111111101;
    assign weights1[46][564] = 16'b1111111111110001;
    assign weights1[46][565] = 16'b0000000000000101;
    assign weights1[46][566] = 16'b0000000000000001;
    assign weights1[46][567] = 16'b1111111111101011;
    assign weights1[46][568] = 16'b1111111111111010;
    assign weights1[46][569] = 16'b0000000000000010;
    assign weights1[46][570] = 16'b1111111111111001;
    assign weights1[46][571] = 16'b0000000000010100;
    assign weights1[46][572] = 16'b1111111111111111;
    assign weights1[46][573] = 16'b1111111111110011;
    assign weights1[46][574] = 16'b1111111111111111;
    assign weights1[46][575] = 16'b0000000000001000;
    assign weights1[46][576] = 16'b1111111111111111;
    assign weights1[46][577] = 16'b0000000000001010;
    assign weights1[46][578] = 16'b1111111111111100;
    assign weights1[46][579] = 16'b1111111111101011;
    assign weights1[46][580] = 16'b0000000000001000;
    assign weights1[46][581] = 16'b0000000000001110;
    assign weights1[46][582] = 16'b0000000000000011;
    assign weights1[46][583] = 16'b0000000000010001;
    assign weights1[46][584] = 16'b1111111111110111;
    assign weights1[46][585] = 16'b0000000000010000;
    assign weights1[46][586] = 16'b0000000000001011;
    assign weights1[46][587] = 16'b0000000000001110;
    assign weights1[46][588] = 16'b1111111111111111;
    assign weights1[46][589] = 16'b0000000000001001;
    assign weights1[46][590] = 16'b0000000000001111;
    assign weights1[46][591] = 16'b0000000000010011;
    assign weights1[46][592] = 16'b0000000000010001;
    assign weights1[46][593] = 16'b0000000000010001;
    assign weights1[46][594] = 16'b1111111111111100;
    assign weights1[46][595] = 16'b0000000000010111;
    assign weights1[46][596] = 16'b1111111111110010;
    assign weights1[46][597] = 16'b0000000000001010;
    assign weights1[46][598] = 16'b0000000000001101;
    assign weights1[46][599] = 16'b0000000000000000;
    assign weights1[46][600] = 16'b0000000000000110;
    assign weights1[46][601] = 16'b0000000000010111;
    assign weights1[46][602] = 16'b1111111111111010;
    assign weights1[46][603] = 16'b0000000000001110;
    assign weights1[46][604] = 16'b0000000000001101;
    assign weights1[46][605] = 16'b0000000000010000;
    assign weights1[46][606] = 16'b0000000000000110;
    assign weights1[46][607] = 16'b0000000000001111;
    assign weights1[46][608] = 16'b1111111111111100;
    assign weights1[46][609] = 16'b1111111111110100;
    assign weights1[46][610] = 16'b0000000000011010;
    assign weights1[46][611] = 16'b0000000000011101;
    assign weights1[46][612] = 16'b0000000000000001;
    assign weights1[46][613] = 16'b0000000000011110;
    assign weights1[46][614] = 16'b0000000000000000;
    assign weights1[46][615] = 16'b0000000000000010;
    assign weights1[46][616] = 16'b1111111111110100;
    assign weights1[46][617] = 16'b1111111111111111;
    assign weights1[46][618] = 16'b0000000000001011;
    assign weights1[46][619] = 16'b1111111111111111;
    assign weights1[46][620] = 16'b1111111111111001;
    assign weights1[46][621] = 16'b1111111111111001;
    assign weights1[46][622] = 16'b1111111111111110;
    assign weights1[46][623] = 16'b1111111111111110;
    assign weights1[46][624] = 16'b0000000000001001;
    assign weights1[46][625] = 16'b1111111111101101;
    assign weights1[46][626] = 16'b0000000000010000;
    assign weights1[46][627] = 16'b1111111111110000;
    assign weights1[46][628] = 16'b0000000000001100;
    assign weights1[46][629] = 16'b1111111111111100;
    assign weights1[46][630] = 16'b0000000000000110;
    assign weights1[46][631] = 16'b0000000000000100;
    assign weights1[46][632] = 16'b1111111111111010;
    assign weights1[46][633] = 16'b1111111111111110;
    assign weights1[46][634] = 16'b0000000000011000;
    assign weights1[46][635] = 16'b1111111111110110;
    assign weights1[46][636] = 16'b0000000000010010;
    assign weights1[46][637] = 16'b1111111111110010;
    assign weights1[46][638] = 16'b0000000000010001;
    assign weights1[46][639] = 16'b0000000000001101;
    assign weights1[46][640] = 16'b1111111111111101;
    assign weights1[46][641] = 16'b0000000000001011;
    assign weights1[46][642] = 16'b1111111111111101;
    assign weights1[46][643] = 16'b0000000000000111;
    assign weights1[46][644] = 16'b1111111111111100;
    assign weights1[46][645] = 16'b1111111111111010;
    assign weights1[46][646] = 16'b1111111111110001;
    assign weights1[46][647] = 16'b1111111111101111;
    assign weights1[46][648] = 16'b1111111111111010;
    assign weights1[46][649] = 16'b0000000000000011;
    assign weights1[46][650] = 16'b1111111111101011;
    assign weights1[46][651] = 16'b1111111111111100;
    assign weights1[46][652] = 16'b1111111111111110;
    assign weights1[46][653] = 16'b0000000000001111;
    assign weights1[46][654] = 16'b1111111111110001;
    assign weights1[46][655] = 16'b1111111111101101;
    assign weights1[46][656] = 16'b1111111111111100;
    assign weights1[46][657] = 16'b1111111111110101;
    assign weights1[46][658] = 16'b0000000000001000;
    assign weights1[46][659] = 16'b0000000000000110;
    assign weights1[46][660] = 16'b0000000000001010;
    assign weights1[46][661] = 16'b1111111111111010;
    assign weights1[46][662] = 16'b1111111111111110;
    assign weights1[46][663] = 16'b0000000000001101;
    assign weights1[46][664] = 16'b0000000000001010;
    assign weights1[46][665] = 16'b0000000000000011;
    assign weights1[46][666] = 16'b1111111111111111;
    assign weights1[46][667] = 16'b0000000000001101;
    assign weights1[46][668] = 16'b0000000000001101;
    assign weights1[46][669] = 16'b0000000000000010;
    assign weights1[46][670] = 16'b0000000000000110;
    assign weights1[46][671] = 16'b1111111111111100;
    assign weights1[46][672] = 16'b1111111111111010;
    assign weights1[46][673] = 16'b0000000000000001;
    assign weights1[46][674] = 16'b1111111111111010;
    assign weights1[46][675] = 16'b0000000000000010;
    assign weights1[46][676] = 16'b1111111111111010;
    assign weights1[46][677] = 16'b0000000000010100;
    assign weights1[46][678] = 16'b0000000000000000;
    assign weights1[46][679] = 16'b0000000000001010;
    assign weights1[46][680] = 16'b1111111111101011;
    assign weights1[46][681] = 16'b0000000000001110;
    assign weights1[46][682] = 16'b1111111111111000;
    assign weights1[46][683] = 16'b0000000000000111;
    assign weights1[46][684] = 16'b0000000000000100;
    assign weights1[46][685] = 16'b1111111111110000;
    assign weights1[46][686] = 16'b1111111111111010;
    assign weights1[46][687] = 16'b0000000000000101;
    assign weights1[46][688] = 16'b1111111111110001;
    assign weights1[46][689] = 16'b0000000000000101;
    assign weights1[46][690] = 16'b1111111111111100;
    assign weights1[46][691] = 16'b1111111111110000;
    assign weights1[46][692] = 16'b0000000000001010;
    assign weights1[46][693] = 16'b0000000000000000;
    assign weights1[46][694] = 16'b1111111111111111;
    assign weights1[46][695] = 16'b0000000000000110;
    assign weights1[46][696] = 16'b0000000000000111;
    assign weights1[46][697] = 16'b1111111111111000;
    assign weights1[46][698] = 16'b1111111111111101;
    assign weights1[46][699] = 16'b1111111111111100;
    assign weights1[46][700] = 16'b1111111111111011;
    assign weights1[46][701] = 16'b0000000000000000;
    assign weights1[46][702] = 16'b1111111111111111;
    assign weights1[46][703] = 16'b0000000000000101;
    assign weights1[46][704] = 16'b1111111111111111;
    assign weights1[46][705] = 16'b0000000000000100;
    assign weights1[46][706] = 16'b0000000000000010;
    assign weights1[46][707] = 16'b0000000000000011;
    assign weights1[46][708] = 16'b1111111111111001;
    assign weights1[46][709] = 16'b0000000000010100;
    assign weights1[46][710] = 16'b1111111111110111;
    assign weights1[46][711] = 16'b1111111111110000;
    assign weights1[46][712] = 16'b0000000000010100;
    assign weights1[46][713] = 16'b0000000000000000;
    assign weights1[46][714] = 16'b0000000000001011;
    assign weights1[46][715] = 16'b0000000000001110;
    assign weights1[46][716] = 16'b0000000000000101;
    assign weights1[46][717] = 16'b0000000000010001;
    assign weights1[46][718] = 16'b0000000000001100;
    assign weights1[46][719] = 16'b1111111111111000;
    assign weights1[46][720] = 16'b0000000000011001;
    assign weights1[46][721] = 16'b0000000000000111;
    assign weights1[46][722] = 16'b0000000000001111;
    assign weights1[46][723] = 16'b0000000000001011;
    assign weights1[46][724] = 16'b0000000000000000;
    assign weights1[46][725] = 16'b1111111111111100;
    assign weights1[46][726] = 16'b1111111111110111;
    assign weights1[46][727] = 16'b1111111111111011;
    assign weights1[46][728] = 16'b1111111111111111;
    assign weights1[46][729] = 16'b1111111111111110;
    assign weights1[46][730] = 16'b1111111111111101;
    assign weights1[46][731] = 16'b1111111111111000;
    assign weights1[46][732] = 16'b1111111111110111;
    assign weights1[46][733] = 16'b1111111111100111;
    assign weights1[46][734] = 16'b1111111111101010;
    assign weights1[46][735] = 16'b1111111111111001;
    assign weights1[46][736] = 16'b0000000000000011;
    assign weights1[46][737] = 16'b0000000000000001;
    assign weights1[46][738] = 16'b1111111111111111;
    assign weights1[46][739] = 16'b0000000000000111;
    assign weights1[46][740] = 16'b1111111111110111;
    assign weights1[46][741] = 16'b0000000000000011;
    assign weights1[46][742] = 16'b1111111111110010;
    assign weights1[46][743] = 16'b1111111111110000;
    assign weights1[46][744] = 16'b1111111111111010;
    assign weights1[46][745] = 16'b1111111111111010;
    assign weights1[46][746] = 16'b0000000000001010;
    assign weights1[46][747] = 16'b0000000000001000;
    assign weights1[46][748] = 16'b1111111111111010;
    assign weights1[46][749] = 16'b1111111111110010;
    assign weights1[46][750] = 16'b1111111111111010;
    assign weights1[46][751] = 16'b1111111111111010;
    assign weights1[46][752] = 16'b0000000000001000;
    assign weights1[46][753] = 16'b0000000000000001;
    assign weights1[46][754] = 16'b0000000000000001;
    assign weights1[46][755] = 16'b0000000000000000;
    assign weights1[46][756] = 16'b1111111111111111;
    assign weights1[46][757] = 16'b1111111111111101;
    assign weights1[46][758] = 16'b1111111111111101;
    assign weights1[46][759] = 16'b1111111111111010;
    assign weights1[46][760] = 16'b1111111111111110;
    assign weights1[46][761] = 16'b0000000000000001;
    assign weights1[46][762] = 16'b1111111111111100;
    assign weights1[46][763] = 16'b1111111111110010;
    assign weights1[46][764] = 16'b1111111111101100;
    assign weights1[46][765] = 16'b0000000000000000;
    assign weights1[46][766] = 16'b1111111111101001;
    assign weights1[46][767] = 16'b1111111111111011;
    assign weights1[46][768] = 16'b1111111111110100;
    assign weights1[46][769] = 16'b1111111111101110;
    assign weights1[46][770] = 16'b1111111111110100;
    assign weights1[46][771] = 16'b0000000000000101;
    assign weights1[46][772] = 16'b1111111111111011;
    assign weights1[46][773] = 16'b1111111111111001;
    assign weights1[46][774] = 16'b1111111111101001;
    assign weights1[46][775] = 16'b1111111111101100;
    assign weights1[46][776] = 16'b1111111111111010;
    assign weights1[46][777] = 16'b1111111111100010;
    assign weights1[46][778] = 16'b1111111111111000;
    assign weights1[46][779] = 16'b0000000000000110;
    assign weights1[46][780] = 16'b0000000000000110;
    assign weights1[46][781] = 16'b0000000000000000;
    assign weights1[46][782] = 16'b0000000000000010;
    assign weights1[46][783] = 16'b0000000000000000;
    assign weights1[47][0] = 16'b0000000000000000;
    assign weights1[47][1] = 16'b0000000000000000;
    assign weights1[47][2] = 16'b0000000000000011;
    assign weights1[47][3] = 16'b0000000000000100;
    assign weights1[47][4] = 16'b0000000000001001;
    assign weights1[47][5] = 16'b0000000000001110;
    assign weights1[47][6] = 16'b0000000000001101;
    assign weights1[47][7] = 16'b0000000000001111;
    assign weights1[47][8] = 16'b0000000000011000;
    assign weights1[47][9] = 16'b0000000000100000;
    assign weights1[47][10] = 16'b0000000000100001;
    assign weights1[47][11] = 16'b0000000000010111;
    assign weights1[47][12] = 16'b0000000000000001;
    assign weights1[47][13] = 16'b0000000000001110;
    assign weights1[47][14] = 16'b0000000000010011;
    assign weights1[47][15] = 16'b0000000000010000;
    assign weights1[47][16] = 16'b0000000000010110;
    assign weights1[47][17] = 16'b0000000000000100;
    assign weights1[47][18] = 16'b0000000000000100;
    assign weights1[47][19] = 16'b1111111111111100;
    assign weights1[47][20] = 16'b0000000000000000;
    assign weights1[47][21] = 16'b0000000000001001;
    assign weights1[47][22] = 16'b0000000000000001;
    assign weights1[47][23] = 16'b1111111111111010;
    assign weights1[47][24] = 16'b0000000000000001;
    assign weights1[47][25] = 16'b0000000000001111;
    assign weights1[47][26] = 16'b0000000000000111;
    assign weights1[47][27] = 16'b1111111111111100;
    assign weights1[47][28] = 16'b0000000000000000;
    assign weights1[47][29] = 16'b0000000000000011;
    assign weights1[47][30] = 16'b0000000000001000;
    assign weights1[47][31] = 16'b0000000000001010;
    assign weights1[47][32] = 16'b0000000000011011;
    assign weights1[47][33] = 16'b0000000000011101;
    assign weights1[47][34] = 16'b0000000000100000;
    assign weights1[47][35] = 16'b0000000000100010;
    assign weights1[47][36] = 16'b0000000000011011;
    assign weights1[47][37] = 16'b0000000000001101;
    assign weights1[47][38] = 16'b0000000000011100;
    assign weights1[47][39] = 16'b0000000000000010;
    assign weights1[47][40] = 16'b0000000000000101;
    assign weights1[47][41] = 16'b0000000000001000;
    assign weights1[47][42] = 16'b1111111111111001;
    assign weights1[47][43] = 16'b1111111111111100;
    assign weights1[47][44] = 16'b0000000000001001;
    assign weights1[47][45] = 16'b0000000000000100;
    assign weights1[47][46] = 16'b0000000000000101;
    assign weights1[47][47] = 16'b1111111111110011;
    assign weights1[47][48] = 16'b1111111111111111;
    assign weights1[47][49] = 16'b1111111111110010;
    assign weights1[47][50] = 16'b1111111111111010;
    assign weights1[47][51] = 16'b1111111111110100;
    assign weights1[47][52] = 16'b0000000000000110;
    assign weights1[47][53] = 16'b0000000000001010;
    assign weights1[47][54] = 16'b0000000000010010;
    assign weights1[47][55] = 16'b0000000000000011;
    assign weights1[47][56] = 16'b0000000000000010;
    assign weights1[47][57] = 16'b0000000000001000;
    assign weights1[47][58] = 16'b0000000000000001;
    assign weights1[47][59] = 16'b0000000000010000;
    assign weights1[47][60] = 16'b0000000000011010;
    assign weights1[47][61] = 16'b0000000000010100;
    assign weights1[47][62] = 16'b0000000000010101;
    assign weights1[47][63] = 16'b0000000000100011;
    assign weights1[47][64] = 16'b0000000000010000;
    assign weights1[47][65] = 16'b0000000000011110;
    assign weights1[47][66] = 16'b0000000000001011;
    assign weights1[47][67] = 16'b0000000000001111;
    assign weights1[47][68] = 16'b0000000000010000;
    assign weights1[47][69] = 16'b0000000000011010;
    assign weights1[47][70] = 16'b0000000000000011;
    assign weights1[47][71] = 16'b0000000000000101;
    assign weights1[47][72] = 16'b1111111111111111;
    assign weights1[47][73] = 16'b0000000000000101;
    assign weights1[47][74] = 16'b0000000000000010;
    assign weights1[47][75] = 16'b1111111111111010;
    assign weights1[47][76] = 16'b1111111111111101;
    assign weights1[47][77] = 16'b0000000000000101;
    assign weights1[47][78] = 16'b0000000000000010;
    assign weights1[47][79] = 16'b1111111111111111;
    assign weights1[47][80] = 16'b0000000000000010;
    assign weights1[47][81] = 16'b1111111111111100;
    assign weights1[47][82] = 16'b0000000000000000;
    assign weights1[47][83] = 16'b1111111111111101;
    assign weights1[47][84] = 16'b0000000000000011;
    assign weights1[47][85] = 16'b0000000000001010;
    assign weights1[47][86] = 16'b0000000000000001;
    assign weights1[47][87] = 16'b0000000000010000;
    assign weights1[47][88] = 16'b0000000000001111;
    assign weights1[47][89] = 16'b0000000000010011;
    assign weights1[47][90] = 16'b0000000000010001;
    assign weights1[47][91] = 16'b0000000000011100;
    assign weights1[47][92] = 16'b0000000000001111;
    assign weights1[47][93] = 16'b0000000000000111;
    assign weights1[47][94] = 16'b0000000000001100;
    assign weights1[47][95] = 16'b0000000000000111;
    assign weights1[47][96] = 16'b0000000000001110;
    assign weights1[47][97] = 16'b0000000000000111;
    assign weights1[47][98] = 16'b1111111111111011;
    assign weights1[47][99] = 16'b0000000000011000;
    assign weights1[47][100] = 16'b0000000000001100;
    assign weights1[47][101] = 16'b1111111111110110;
    assign weights1[47][102] = 16'b0000000000000110;
    assign weights1[47][103] = 16'b0000000000001100;
    assign weights1[47][104] = 16'b0000000000001010;
    assign weights1[47][105] = 16'b0000000000000001;
    assign weights1[47][106] = 16'b0000000000000001;
    assign weights1[47][107] = 16'b1111111111110100;
    assign weights1[47][108] = 16'b0000000000000000;
    assign weights1[47][109] = 16'b1111111111111001;
    assign weights1[47][110] = 16'b0000000000001011;
    assign weights1[47][111] = 16'b0000000000001100;
    assign weights1[47][112] = 16'b0000000000000110;
    assign weights1[47][113] = 16'b0000000000000111;
    assign weights1[47][114] = 16'b0000000000000111;
    assign weights1[47][115] = 16'b1111111111111001;
    assign weights1[47][116] = 16'b1111111111110010;
    assign weights1[47][117] = 16'b0000000000000010;
    assign weights1[47][118] = 16'b0000000000001000;
    assign weights1[47][119] = 16'b0000000000010011;
    assign weights1[47][120] = 16'b0000000000001010;
    assign weights1[47][121] = 16'b0000000000010101;
    assign weights1[47][122] = 16'b0000000000011000;
    assign weights1[47][123] = 16'b0000000000110000;
    assign weights1[47][124] = 16'b0000000000001100;
    assign weights1[47][125] = 16'b0000000000010011;
    assign weights1[47][126] = 16'b0000000000010100;
    assign weights1[47][127] = 16'b1111111111110100;
    assign weights1[47][128] = 16'b0000000000011010;
    assign weights1[47][129] = 16'b1111111111111110;
    assign weights1[47][130] = 16'b0000000000000101;
    assign weights1[47][131] = 16'b1111111111110111;
    assign weights1[47][132] = 16'b0000000000000011;
    assign weights1[47][133] = 16'b1111111111111010;
    assign weights1[47][134] = 16'b1111111111111101;
    assign weights1[47][135] = 16'b0000000000001001;
    assign weights1[47][136] = 16'b0000000000001001;
    assign weights1[47][137] = 16'b0000000000001011;
    assign weights1[47][138] = 16'b0000000000000011;
    assign weights1[47][139] = 16'b0000000000000101;
    assign weights1[47][140] = 16'b0000000000000101;
    assign weights1[47][141] = 16'b0000000000001001;
    assign weights1[47][142] = 16'b0000000000000001;
    assign weights1[47][143] = 16'b1111111111101110;
    assign weights1[47][144] = 16'b1111111111111011;
    assign weights1[47][145] = 16'b0000000000001010;
    assign weights1[47][146] = 16'b0000000000001010;
    assign weights1[47][147] = 16'b1111111111110100;
    assign weights1[47][148] = 16'b0000000000011011;
    assign weights1[47][149] = 16'b0000000000010001;
    assign weights1[47][150] = 16'b0000000000000110;
    assign weights1[47][151] = 16'b0000000000000110;
    assign weights1[47][152] = 16'b0000000000011000;
    assign weights1[47][153] = 16'b0000000000011101;
    assign weights1[47][154] = 16'b0000000000010010;
    assign weights1[47][155] = 16'b0000000000001101;
    assign weights1[47][156] = 16'b0000000000010011;
    assign weights1[47][157] = 16'b0000000000011001;
    assign weights1[47][158] = 16'b0000000000001100;
    assign weights1[47][159] = 16'b0000000000000010;
    assign weights1[47][160] = 16'b0000000000000110;
    assign weights1[47][161] = 16'b0000000000001111;
    assign weights1[47][162] = 16'b0000000000001101;
    assign weights1[47][163] = 16'b0000000000000010;
    assign weights1[47][164] = 16'b1111111111111000;
    assign weights1[47][165] = 16'b0000000000000001;
    assign weights1[47][166] = 16'b0000000000001001;
    assign weights1[47][167] = 16'b0000000000000010;
    assign weights1[47][168] = 16'b0000000000000101;
    assign weights1[47][169] = 16'b1111111111111010;
    assign weights1[47][170] = 16'b1111111111110010;
    assign weights1[47][171] = 16'b1111111111101100;
    assign weights1[47][172] = 16'b1111111111101000;
    assign weights1[47][173] = 16'b1111111111101000;
    assign weights1[47][174] = 16'b0000000000000000;
    assign weights1[47][175] = 16'b1111111111101111;
    assign weights1[47][176] = 16'b1111111111101100;
    assign weights1[47][177] = 16'b1111111111110000;
    assign weights1[47][178] = 16'b1111111111101100;
    assign weights1[47][179] = 16'b1111111111111001;
    assign weights1[47][180] = 16'b1111111111111011;
    assign weights1[47][181] = 16'b0000000000001001;
    assign weights1[47][182] = 16'b0000000000000011;
    assign weights1[47][183] = 16'b0000000000001010;
    assign weights1[47][184] = 16'b0000000000000011;
    assign weights1[47][185] = 16'b1111111111110111;
    assign weights1[47][186] = 16'b0000000000010001;
    assign weights1[47][187] = 16'b0000000000000110;
    assign weights1[47][188] = 16'b0000000000001010;
    assign weights1[47][189] = 16'b0000000000000100;
    assign weights1[47][190] = 16'b0000000000001010;
    assign weights1[47][191] = 16'b0000000000001100;
    assign weights1[47][192] = 16'b0000000000010001;
    assign weights1[47][193] = 16'b0000000000000100;
    assign weights1[47][194] = 16'b0000000000000001;
    assign weights1[47][195] = 16'b0000000000001001;
    assign weights1[47][196] = 16'b1111111111110101;
    assign weights1[47][197] = 16'b1111111111100101;
    assign weights1[47][198] = 16'b1111111111100100;
    assign weights1[47][199] = 16'b1111111111011011;
    assign weights1[47][200] = 16'b1111111111011101;
    assign weights1[47][201] = 16'b1111111111001010;
    assign weights1[47][202] = 16'b1111111111100000;
    assign weights1[47][203] = 16'b1111111111011000;
    assign weights1[47][204] = 16'b1111111111100011;
    assign weights1[47][205] = 16'b1111111111101100;
    assign weights1[47][206] = 16'b1111111111101011;
    assign weights1[47][207] = 16'b1111111111101000;
    assign weights1[47][208] = 16'b1111111111100111;
    assign weights1[47][209] = 16'b1111111111101011;
    assign weights1[47][210] = 16'b1111111111110101;
    assign weights1[47][211] = 16'b1111111111101001;
    assign weights1[47][212] = 16'b0000000000000010;
    assign weights1[47][213] = 16'b1111111111110100;
    assign weights1[47][214] = 16'b1111111111111100;
    assign weights1[47][215] = 16'b1111111111111010;
    assign weights1[47][216] = 16'b1111111111111110;
    assign weights1[47][217] = 16'b1111111111111001;
    assign weights1[47][218] = 16'b1111111111111011;
    assign weights1[47][219] = 16'b1111111111111011;
    assign weights1[47][220] = 16'b1111111111110111;
    assign weights1[47][221] = 16'b0000000000000000;
    assign weights1[47][222] = 16'b0000000000001110;
    assign weights1[47][223] = 16'b0000000000001110;
    assign weights1[47][224] = 16'b1111111111110001;
    assign weights1[47][225] = 16'b1111111111011000;
    assign weights1[47][226] = 16'b1111111111011011;
    assign weights1[47][227] = 16'b1111111111010011;
    assign weights1[47][228] = 16'b1111111111001111;
    assign weights1[47][229] = 16'b1111111111010011;
    assign weights1[47][230] = 16'b1111111111011001;
    assign weights1[47][231] = 16'b1111111111101011;
    assign weights1[47][232] = 16'b1111111111010101;
    assign weights1[47][233] = 16'b1111111111101111;
    assign weights1[47][234] = 16'b1111111111111110;
    assign weights1[47][235] = 16'b1111111111110100;
    assign weights1[47][236] = 16'b1111111111100001;
    assign weights1[47][237] = 16'b0000000000001110;
    assign weights1[47][238] = 16'b1111111111110001;
    assign weights1[47][239] = 16'b0000000000001100;
    assign weights1[47][240] = 16'b1111111111101011;
    assign weights1[47][241] = 16'b0000000000000001;
    assign weights1[47][242] = 16'b0000000000000010;
    assign weights1[47][243] = 16'b1111111111101000;
    assign weights1[47][244] = 16'b0000000000000100;
    assign weights1[47][245] = 16'b1111111111111001;
    assign weights1[47][246] = 16'b0000000000010010;
    assign weights1[47][247] = 16'b0000000000000110;
    assign weights1[47][248] = 16'b1111111111101110;
    assign weights1[47][249] = 16'b0000000000000010;
    assign weights1[47][250] = 16'b1111111111111001;
    assign weights1[47][251] = 16'b0000000000000111;
    assign weights1[47][252] = 16'b1111111111100110;
    assign weights1[47][253] = 16'b1111111111010011;
    assign weights1[47][254] = 16'b1111111111010110;
    assign weights1[47][255] = 16'b1111111111010111;
    assign weights1[47][256] = 16'b1111111111101100;
    assign weights1[47][257] = 16'b1111111111110010;
    assign weights1[47][258] = 16'b0000000000000010;
    assign weights1[47][259] = 16'b0000000000000110;
    assign weights1[47][260] = 16'b1111111111101110;
    assign weights1[47][261] = 16'b1111111111110000;
    assign weights1[47][262] = 16'b1111111111111110;
    assign weights1[47][263] = 16'b0000000000001111;
    assign weights1[47][264] = 16'b0000000000000101;
    assign weights1[47][265] = 16'b0000000000001110;
    assign weights1[47][266] = 16'b0000000000001010;
    assign weights1[47][267] = 16'b0000000000000100;
    assign weights1[47][268] = 16'b0000000000010001;
    assign weights1[47][269] = 16'b0000000000000101;
    assign weights1[47][270] = 16'b0000000000000110;
    assign weights1[47][271] = 16'b1111111111111000;
    assign weights1[47][272] = 16'b1111111111110100;
    assign weights1[47][273] = 16'b1111111111111010;
    assign weights1[47][274] = 16'b1111111111101101;
    assign weights1[47][275] = 16'b1111111111111101;
    assign weights1[47][276] = 16'b1111111111111010;
    assign weights1[47][277] = 16'b0000000000000001;
    assign weights1[47][278] = 16'b0000000000000011;
    assign weights1[47][279] = 16'b0000000000000101;
    assign weights1[47][280] = 16'b1111111111011110;
    assign weights1[47][281] = 16'b1111111111000101;
    assign weights1[47][282] = 16'b1111111111000101;
    assign weights1[47][283] = 16'b1111111111001100;
    assign weights1[47][284] = 16'b1111111111011111;
    assign weights1[47][285] = 16'b1111111111111101;
    assign weights1[47][286] = 16'b0000000000000000;
    assign weights1[47][287] = 16'b0000000000010011;
    assign weights1[47][288] = 16'b0000000000000110;
    assign weights1[47][289] = 16'b0000000000100101;
    assign weights1[47][290] = 16'b0000000000001111;
    assign weights1[47][291] = 16'b0000000000010101;
    assign weights1[47][292] = 16'b0000000000100101;
    assign weights1[47][293] = 16'b0000000000011100;
    assign weights1[47][294] = 16'b0000000000001101;
    assign weights1[47][295] = 16'b0000000000010010;
    assign weights1[47][296] = 16'b1111111111111100;
    assign weights1[47][297] = 16'b0000000000001011;
    assign weights1[47][298] = 16'b0000000000001000;
    assign weights1[47][299] = 16'b0000000000000101;
    assign weights1[47][300] = 16'b0000000000001001;
    assign weights1[47][301] = 16'b0000000000010000;
    assign weights1[47][302] = 16'b1111111111111110;
    assign weights1[47][303] = 16'b0000000000000100;
    assign weights1[47][304] = 16'b1111111111111110;
    assign weights1[47][305] = 16'b1111111111110111;
    assign weights1[47][306] = 16'b1111111111110011;
    assign weights1[47][307] = 16'b0000000000000000;
    assign weights1[47][308] = 16'b1111111111100000;
    assign weights1[47][309] = 16'b1111111111000101;
    assign weights1[47][310] = 16'b1111111110110100;
    assign weights1[47][311] = 16'b1111111110101001;
    assign weights1[47][312] = 16'b1111111110111010;
    assign weights1[47][313] = 16'b1111111111000111;
    assign weights1[47][314] = 16'b1111111111101001;
    assign weights1[47][315] = 16'b0000000000000100;
    assign weights1[47][316] = 16'b0000000000111010;
    assign weights1[47][317] = 16'b0000000000100010;
    assign weights1[47][318] = 16'b0000000000110110;
    assign weights1[47][319] = 16'b0000000000100011;
    assign weights1[47][320] = 16'b0000000000100111;
    assign weights1[47][321] = 16'b0000000000011011;
    assign weights1[47][322] = 16'b0000000000011110;
    assign weights1[47][323] = 16'b0000000000010111;
    assign weights1[47][324] = 16'b0000000000010111;
    assign weights1[47][325] = 16'b0000000000011010;
    assign weights1[47][326] = 16'b0000000000000011;
    assign weights1[47][327] = 16'b0000000000001001;
    assign weights1[47][328] = 16'b0000000000001000;
    assign weights1[47][329] = 16'b0000000000001010;
    assign weights1[47][330] = 16'b1111111111111101;
    assign weights1[47][331] = 16'b0000000000010001;
    assign weights1[47][332] = 16'b1111111111111100;
    assign weights1[47][333] = 16'b1111111111101011;
    assign weights1[47][334] = 16'b0000000000000101;
    assign weights1[47][335] = 16'b1111111111111100;
    assign weights1[47][336] = 16'b1111111111011010;
    assign weights1[47][337] = 16'b1111111111000000;
    assign weights1[47][338] = 16'b1111111110011101;
    assign weights1[47][339] = 16'b1111111110101000;
    assign weights1[47][340] = 16'b1111111110001001;
    assign weights1[47][341] = 16'b1111111110000010;
    assign weights1[47][342] = 16'b1111111101111110;
    assign weights1[47][343] = 16'b1111111110110100;
    assign weights1[47][344] = 16'b1111111111011100;
    assign weights1[47][345] = 16'b1111111111111110;
    assign weights1[47][346] = 16'b0000000000100000;
    assign weights1[47][347] = 16'b0000000000100101;
    assign weights1[47][348] = 16'b0000000000101010;
    assign weights1[47][349] = 16'b0000000000101111;
    assign weights1[47][350] = 16'b0000000000010011;
    assign weights1[47][351] = 16'b0000000000010010;
    assign weights1[47][352] = 16'b0000000000000111;
    assign weights1[47][353] = 16'b0000000000000000;
    assign weights1[47][354] = 16'b0000000000000010;
    assign weights1[47][355] = 16'b1111111111101111;
    assign weights1[47][356] = 16'b1111111111110111;
    assign weights1[47][357] = 16'b1111111111110110;
    assign weights1[47][358] = 16'b1111111111101101;
    assign weights1[47][359] = 16'b1111111111110110;
    assign weights1[47][360] = 16'b1111111111110110;
    assign weights1[47][361] = 16'b1111111111101110;
    assign weights1[47][362] = 16'b1111111111111010;
    assign weights1[47][363] = 16'b1111111111111100;
    assign weights1[47][364] = 16'b1111111111011111;
    assign weights1[47][365] = 16'b1111111111000010;
    assign weights1[47][366] = 16'b1111111110101111;
    assign weights1[47][367] = 16'b1111111110001111;
    assign weights1[47][368] = 16'b1111111110000010;
    assign weights1[47][369] = 16'b1111111101010111;
    assign weights1[47][370] = 16'b1111111100110110;
    assign weights1[47][371] = 16'b1111111100101101;
    assign weights1[47][372] = 16'b1111111100100000;
    assign weights1[47][373] = 16'b1111111101110101;
    assign weights1[47][374] = 16'b1111111110110100;
    assign weights1[47][375] = 16'b1111111111010100;
    assign weights1[47][376] = 16'b1111111111110111;
    assign weights1[47][377] = 16'b0000000000010000;
    assign weights1[47][378] = 16'b1111111111111011;
    assign weights1[47][379] = 16'b0000000000001001;
    assign weights1[47][380] = 16'b1111111111110000;
    assign weights1[47][381] = 16'b1111111111111110;
    assign weights1[47][382] = 16'b1111111111110100;
    assign weights1[47][383] = 16'b0000000000001011;
    assign weights1[47][384] = 16'b1111111111110101;
    assign weights1[47][385] = 16'b1111111111111001;
    assign weights1[47][386] = 16'b0000000000000101;
    assign weights1[47][387] = 16'b1111111111110000;
    assign weights1[47][388] = 16'b1111111111111011;
    assign weights1[47][389] = 16'b1111111111111111;
    assign weights1[47][390] = 16'b1111111111111101;
    assign weights1[47][391] = 16'b1111111111100111;
    assign weights1[47][392] = 16'b1111111111110111;
    assign weights1[47][393] = 16'b1111111111100100;
    assign weights1[47][394] = 16'b1111111111010110;
    assign weights1[47][395] = 16'b1111111111000110;
    assign weights1[47][396] = 16'b1111111110111110;
    assign weights1[47][397] = 16'b1111111110011111;
    assign weights1[47][398] = 16'b1111111101110011;
    assign weights1[47][399] = 16'b1111111101001010;
    assign weights1[47][400] = 16'b1111111100001001;
    assign weights1[47][401] = 16'b1111111011101110;
    assign weights1[47][402] = 16'b1111111011110100;
    assign weights1[47][403] = 16'b1111111100010000;
    assign weights1[47][404] = 16'b1111111101011000;
    assign weights1[47][405] = 16'b1111111110011000;
    assign weights1[47][406] = 16'b1111111110110001;
    assign weights1[47][407] = 16'b1111111111001110;
    assign weights1[47][408] = 16'b1111111111011111;
    assign weights1[47][409] = 16'b1111111111100111;
    assign weights1[47][410] = 16'b1111111111010101;
    assign weights1[47][411] = 16'b1111111111101000;
    assign weights1[47][412] = 16'b1111111111111111;
    assign weights1[47][413] = 16'b0000000000000011;
    assign weights1[47][414] = 16'b1111111111111111;
    assign weights1[47][415] = 16'b1111111111111011;
    assign weights1[47][416] = 16'b0000000000010000;
    assign weights1[47][417] = 16'b0000000000001100;
    assign weights1[47][418] = 16'b1111111111110010;
    assign weights1[47][419] = 16'b1111111111101100;
    assign weights1[47][420] = 16'b0000000000010000;
    assign weights1[47][421] = 16'b1111111111110100;
    assign weights1[47][422] = 16'b0000000000010001;
    assign weights1[47][423] = 16'b0000000000000010;
    assign weights1[47][424] = 16'b0000000000000010;
    assign weights1[47][425] = 16'b1111111111111010;
    assign weights1[47][426] = 16'b0000000000001010;
    assign weights1[47][427] = 16'b1111111111010001;
    assign weights1[47][428] = 16'b1111111111000100;
    assign weights1[47][429] = 16'b1111111110010101;
    assign weights1[47][430] = 16'b1111111101011111;
    assign weights1[47][431] = 16'b1111111101001001;
    assign weights1[47][432] = 16'b1111111101011011;
    assign weights1[47][433] = 16'b1111111101100011;
    assign weights1[47][434] = 16'b1111111110010000;
    assign weights1[47][435] = 16'b1111111110010101;
    assign weights1[47][436] = 16'b1111111111000000;
    assign weights1[47][437] = 16'b1111111110111000;
    assign weights1[47][438] = 16'b1111111111110100;
    assign weights1[47][439] = 16'b1111111111110111;
    assign weights1[47][440] = 16'b1111111111101111;
    assign weights1[47][441] = 16'b1111111111111101;
    assign weights1[47][442] = 16'b0000000000000100;
    assign weights1[47][443] = 16'b1111111111111001;
    assign weights1[47][444] = 16'b0000000000000111;
    assign weights1[47][445] = 16'b0000000000010101;
    assign weights1[47][446] = 16'b0000000000010001;
    assign weights1[47][447] = 16'b1111111111101111;
    assign weights1[47][448] = 16'b0000000000011101;
    assign weights1[47][449] = 16'b0000000000010011;
    assign weights1[47][450] = 16'b0000000000100101;
    assign weights1[47][451] = 16'b0000000000010111;
    assign weights1[47][452] = 16'b0000000000111011;
    assign weights1[47][453] = 16'b0000000000100100;
    assign weights1[47][454] = 16'b0000000000101010;
    assign weights1[47][455] = 16'b0000000001000011;
    assign weights1[47][456] = 16'b0000000000101001;
    assign weights1[47][457] = 16'b0000000000101001;
    assign weights1[47][458] = 16'b0000000000001101;
    assign weights1[47][459] = 16'b0000000000001110;
    assign weights1[47][460] = 16'b1111111111110100;
    assign weights1[47][461] = 16'b1111111111110101;
    assign weights1[47][462] = 16'b1111111111011110;
    assign weights1[47][463] = 16'b1111111111100000;
    assign weights1[47][464] = 16'b1111111111010100;
    assign weights1[47][465] = 16'b1111111111011011;
    assign weights1[47][466] = 16'b1111111111101001;
    assign weights1[47][467] = 16'b1111111111110000;
    assign weights1[47][468] = 16'b1111111111111011;
    assign weights1[47][469] = 16'b1111111111110010;
    assign weights1[47][470] = 16'b0000000000000010;
    assign weights1[47][471] = 16'b0000000000000000;
    assign weights1[47][472] = 16'b0000000000001000;
    assign weights1[47][473] = 16'b0000000000000000;
    assign weights1[47][474] = 16'b1111111111111100;
    assign weights1[47][475] = 16'b1111111111110011;
    assign weights1[47][476] = 16'b0000000000100010;
    assign weights1[47][477] = 16'b0000000000100110;
    assign weights1[47][478] = 16'b0000000000100111;
    assign weights1[47][479] = 16'b0000000000101000;
    assign weights1[47][480] = 16'b0000000000101110;
    assign weights1[47][481] = 16'b0000000000111000;
    assign weights1[47][482] = 16'b0000000000110110;
    assign weights1[47][483] = 16'b0000000001000001;
    assign weights1[47][484] = 16'b0000000001011110;
    assign weights1[47][485] = 16'b0000000001000001;
    assign weights1[47][486] = 16'b0000000001001110;
    assign weights1[47][487] = 16'b0000000001010001;
    assign weights1[47][488] = 16'b0000000000101010;
    assign weights1[47][489] = 16'b0000000000100100;
    assign weights1[47][490] = 16'b1111111111111110;
    assign weights1[47][491] = 16'b0000000000001011;
    assign weights1[47][492] = 16'b0000000000000100;
    assign weights1[47][493] = 16'b0000000000001100;
    assign weights1[47][494] = 16'b1111111111101111;
    assign weights1[47][495] = 16'b0000000000001001;
    assign weights1[47][496] = 16'b1111111111101000;
    assign weights1[47][497] = 16'b1111111111110001;
    assign weights1[47][498] = 16'b1111111111110110;
    assign weights1[47][499] = 16'b1111111111111010;
    assign weights1[47][500] = 16'b1111111111110000;
    assign weights1[47][501] = 16'b1111111111110101;
    assign weights1[47][502] = 16'b1111111111101110;
    assign weights1[47][503] = 16'b1111111111111011;
    assign weights1[47][504] = 16'b0000000000101000;
    assign weights1[47][505] = 16'b0000000000011100;
    assign weights1[47][506] = 16'b0000000000101110;
    assign weights1[47][507] = 16'b0000000000111110;
    assign weights1[47][508] = 16'b0000000000100000;
    assign weights1[47][509] = 16'b1111111111111111;
    assign weights1[47][510] = 16'b0000000000110011;
    assign weights1[47][511] = 16'b0000000000101100;
    assign weights1[47][512] = 16'b0000000000100011;
    assign weights1[47][513] = 16'b0000000000101100;
    assign weights1[47][514] = 16'b0000000000101101;
    assign weights1[47][515] = 16'b0000000000110011;
    assign weights1[47][516] = 16'b0000000000101010;
    assign weights1[47][517] = 16'b0000000000001111;
    assign weights1[47][518] = 16'b0000000000010011;
    assign weights1[47][519] = 16'b0000000000011100;
    assign weights1[47][520] = 16'b1111111111111000;
    assign weights1[47][521] = 16'b0000000000000010;
    assign weights1[47][522] = 16'b1111111111110101;
    assign weights1[47][523] = 16'b1111111111110000;
    assign weights1[47][524] = 16'b1111111111110110;
    assign weights1[47][525] = 16'b1111111111111110;
    assign weights1[47][526] = 16'b1111111111111100;
    assign weights1[47][527] = 16'b1111111111111001;
    assign weights1[47][528] = 16'b0000000000001110;
    assign weights1[47][529] = 16'b0000000000000010;
    assign weights1[47][530] = 16'b1111111111110000;
    assign weights1[47][531] = 16'b0000000000001010;
    assign weights1[47][532] = 16'b0000000000001011;
    assign weights1[47][533] = 16'b0000000000000101;
    assign weights1[47][534] = 16'b0000000000011000;
    assign weights1[47][535] = 16'b0000000000101110;
    assign weights1[47][536] = 16'b0000000000011000;
    assign weights1[47][537] = 16'b0000000000001101;
    assign weights1[47][538] = 16'b0000000000100110;
    assign weights1[47][539] = 16'b0000000000011000;
    assign weights1[47][540] = 16'b0000000000001010;
    assign weights1[47][541] = 16'b0000000000011010;
    assign weights1[47][542] = 16'b0000000000100001;
    assign weights1[47][543] = 16'b0000000000011001;
    assign weights1[47][544] = 16'b0000000000100010;
    assign weights1[47][545] = 16'b0000000000011111;
    assign weights1[47][546] = 16'b0000000000010011;
    assign weights1[47][547] = 16'b0000000000001011;
    assign weights1[47][548] = 16'b0000000000010100;
    assign weights1[47][549] = 16'b0000000000010011;
    assign weights1[47][550] = 16'b0000000000000111;
    assign weights1[47][551] = 16'b0000000000001001;
    assign weights1[47][552] = 16'b1111111111110111;
    assign weights1[47][553] = 16'b1111111111111100;
    assign weights1[47][554] = 16'b1111111111011111;
    assign weights1[47][555] = 16'b1111111111110101;
    assign weights1[47][556] = 16'b1111111111100111;
    assign weights1[47][557] = 16'b1111111111101000;
    assign weights1[47][558] = 16'b1111111111110001;
    assign weights1[47][559] = 16'b1111111111111111;
    assign weights1[47][560] = 16'b0000000000000010;
    assign weights1[47][561] = 16'b0000000000001000;
    assign weights1[47][562] = 16'b0000000000000111;
    assign weights1[47][563] = 16'b1111111111111000;
    assign weights1[47][564] = 16'b1111111111001101;
    assign weights1[47][565] = 16'b0000000000000100;
    assign weights1[47][566] = 16'b1111111111111000;
    assign weights1[47][567] = 16'b0000000000011101;
    assign weights1[47][568] = 16'b0000000000101111;
    assign weights1[47][569] = 16'b0000000000000100;
    assign weights1[47][570] = 16'b0000000000000111;
    assign weights1[47][571] = 16'b0000000000000110;
    assign weights1[47][572] = 16'b0000000000001110;
    assign weights1[47][573] = 16'b0000000000010101;
    assign weights1[47][574] = 16'b0000000000000110;
    assign weights1[47][575] = 16'b0000000000010010;
    assign weights1[47][576] = 16'b0000000000010000;
    assign weights1[47][577] = 16'b1111111111111001;
    assign weights1[47][578] = 16'b0000000000000101;
    assign weights1[47][579] = 16'b0000000000001101;
    assign weights1[47][580] = 16'b0000000000001000;
    assign weights1[47][581] = 16'b0000000000001001;
    assign weights1[47][582] = 16'b0000000000001001;
    assign weights1[47][583] = 16'b1111111111110010;
    assign weights1[47][584] = 16'b1111111111110001;
    assign weights1[47][585] = 16'b1111111111110011;
    assign weights1[47][586] = 16'b1111111111111100;
    assign weights1[47][587] = 16'b1111111111111010;
    assign weights1[47][588] = 16'b0000000000000100;
    assign weights1[47][589] = 16'b0000000000000101;
    assign weights1[47][590] = 16'b0000000000001101;
    assign weights1[47][591] = 16'b1111111111101101;
    assign weights1[47][592] = 16'b1111111111100011;
    assign weights1[47][593] = 16'b1111111111100101;
    assign weights1[47][594] = 16'b1111111111100001;
    assign weights1[47][595] = 16'b1111111111111000;
    assign weights1[47][596] = 16'b0000000000000001;
    assign weights1[47][597] = 16'b1111111111111101;
    assign weights1[47][598] = 16'b1111111111101111;
    assign weights1[47][599] = 16'b0000000000000000;
    assign weights1[47][600] = 16'b0000000000000100;
    assign weights1[47][601] = 16'b1111111111110110;
    assign weights1[47][602] = 16'b1111111111110101;
    assign weights1[47][603] = 16'b1111111111111110;
    assign weights1[47][604] = 16'b1111111111110010;
    assign weights1[47][605] = 16'b0000000000011010;
    assign weights1[47][606] = 16'b1111111111111110;
    assign weights1[47][607] = 16'b0000000000001000;
    assign weights1[47][608] = 16'b1111111111110101;
    assign weights1[47][609] = 16'b1111111111111111;
    assign weights1[47][610] = 16'b1111111111110110;
    assign weights1[47][611] = 16'b0000000000000010;
    assign weights1[47][612] = 16'b0000000000000110;
    assign weights1[47][613] = 16'b0000000000000000;
    assign weights1[47][614] = 16'b0000000000000001;
    assign weights1[47][615] = 16'b1111111111111011;
    assign weights1[47][616] = 16'b1111111111111000;
    assign weights1[47][617] = 16'b0000000000000011;
    assign weights1[47][618] = 16'b0000000000001100;
    assign weights1[47][619] = 16'b0000000000001110;
    assign weights1[47][620] = 16'b1111111111101101;
    assign weights1[47][621] = 16'b1111111111100011;
    assign weights1[47][622] = 16'b1111111111101110;
    assign weights1[47][623] = 16'b1111111111101111;
    assign weights1[47][624] = 16'b1111111111110001;
    assign weights1[47][625] = 16'b0000000000000000;
    assign weights1[47][626] = 16'b1111111111111110;
    assign weights1[47][627] = 16'b1111111111110100;
    assign weights1[47][628] = 16'b1111111111110111;
    assign weights1[47][629] = 16'b0000000000001001;
    assign weights1[47][630] = 16'b0000000000000000;
    assign weights1[47][631] = 16'b0000000000011000;
    assign weights1[47][632] = 16'b0000000000001000;
    assign weights1[47][633] = 16'b1111111111111011;
    assign weights1[47][634] = 16'b1111111111110110;
    assign weights1[47][635] = 16'b1111111111110101;
    assign weights1[47][636] = 16'b1111111111111010;
    assign weights1[47][637] = 16'b0000000000001001;
    assign weights1[47][638] = 16'b0000000000001001;
    assign weights1[47][639] = 16'b0000000000001011;
    assign weights1[47][640] = 16'b0000000000000100;
    assign weights1[47][641] = 16'b0000000000001101;
    assign weights1[47][642] = 16'b0000000000000011;
    assign weights1[47][643] = 16'b0000000000000110;
    assign weights1[47][644] = 16'b1111111111111101;
    assign weights1[47][645] = 16'b0000000000000011;
    assign weights1[47][646] = 16'b0000000000000101;
    assign weights1[47][647] = 16'b0000000000000100;
    assign weights1[47][648] = 16'b1111111111110010;
    assign weights1[47][649] = 16'b1111111111101001;
    assign weights1[47][650] = 16'b1111111111011111;
    assign weights1[47][651] = 16'b1111111111000011;
    assign weights1[47][652] = 16'b1111111111100011;
    assign weights1[47][653] = 16'b1111111111101001;
    assign weights1[47][654] = 16'b1111111111110100;
    assign weights1[47][655] = 16'b0000000000000100;
    assign weights1[47][656] = 16'b0000000000000100;
    assign weights1[47][657] = 16'b1111111111111101;
    assign weights1[47][658] = 16'b1111111111100101;
    assign weights1[47][659] = 16'b1111111111101101;
    assign weights1[47][660] = 16'b0000000000000000;
    assign weights1[47][661] = 16'b1111111111110011;
    assign weights1[47][662] = 16'b1111111111111011;
    assign weights1[47][663] = 16'b0000000000100010;
    assign weights1[47][664] = 16'b0000000000001101;
    assign weights1[47][665] = 16'b0000000000010001;
    assign weights1[47][666] = 16'b0000000000011010;
    assign weights1[47][667] = 16'b0000000000010010;
    assign weights1[47][668] = 16'b0000000000011011;
    assign weights1[47][669] = 16'b0000000000011101;
    assign weights1[47][670] = 16'b0000000000000101;
    assign weights1[47][671] = 16'b0000000000000100;
    assign weights1[47][672] = 16'b0000000000000000;
    assign weights1[47][673] = 16'b1111111111111101;
    assign weights1[47][674] = 16'b0000000000000111;
    assign weights1[47][675] = 16'b1111111111111101;
    assign weights1[47][676] = 16'b1111111111111110;
    assign weights1[47][677] = 16'b0000000000000100;
    assign weights1[47][678] = 16'b1111111111101011;
    assign weights1[47][679] = 16'b1111111111011010;
    assign weights1[47][680] = 16'b1111111111001101;
    assign weights1[47][681] = 16'b1111111111001111;
    assign weights1[47][682] = 16'b1111111111001101;
    assign weights1[47][683] = 16'b1111111111011100;
    assign weights1[47][684] = 16'b1111111111011010;
    assign weights1[47][685] = 16'b1111111111100100;
    assign weights1[47][686] = 16'b1111111111111010;
    assign weights1[47][687] = 16'b1111111111101100;
    assign weights1[47][688] = 16'b1111111111110010;
    assign weights1[47][689] = 16'b1111111111111001;
    assign weights1[47][690] = 16'b0000000000011000;
    assign weights1[47][691] = 16'b0000000000010001;
    assign weights1[47][692] = 16'b1111111111111101;
    assign weights1[47][693] = 16'b0000000000001101;
    assign weights1[47][694] = 16'b0000000000001100;
    assign weights1[47][695] = 16'b0000000000001000;
    assign weights1[47][696] = 16'b0000000000100011;
    assign weights1[47][697] = 16'b0000000000010110;
    assign weights1[47][698] = 16'b0000000000001110;
    assign weights1[47][699] = 16'b0000000000000010;
    assign weights1[47][700] = 16'b1111111111111111;
    assign weights1[47][701] = 16'b1111111111111100;
    assign weights1[47][702] = 16'b0000000000000110;
    assign weights1[47][703] = 16'b1111111111111100;
    assign weights1[47][704] = 16'b0000000000001110;
    assign weights1[47][705] = 16'b1111111111110101;
    assign weights1[47][706] = 16'b1111111111111000;
    assign weights1[47][707] = 16'b1111111111111110;
    assign weights1[47][708] = 16'b1111111111110100;
    assign weights1[47][709] = 16'b0000000000000110;
    assign weights1[47][710] = 16'b1111111111101011;
    assign weights1[47][711] = 16'b1111111111101111;
    assign weights1[47][712] = 16'b1111111111111010;
    assign weights1[47][713] = 16'b1111111111101110;
    assign weights1[47][714] = 16'b1111111111110110;
    assign weights1[47][715] = 16'b0000000000001110;
    assign weights1[47][716] = 16'b1111111111111100;
    assign weights1[47][717] = 16'b0000000000001101;
    assign weights1[47][718] = 16'b1111111111111101;
    assign weights1[47][719] = 16'b0000000000000111;
    assign weights1[47][720] = 16'b0000000000001000;
    assign weights1[47][721] = 16'b0000000000000000;
    assign weights1[47][722] = 16'b0000000000001010;
    assign weights1[47][723] = 16'b0000000000001110;
    assign weights1[47][724] = 16'b0000000000010001;
    assign weights1[47][725] = 16'b0000000000001100;
    assign weights1[47][726] = 16'b1111111111111111;
    assign weights1[47][727] = 16'b0000000000000001;
    assign weights1[47][728] = 16'b0000000000000110;
    assign weights1[47][729] = 16'b0000000000000100;
    assign weights1[47][730] = 16'b0000000000000100;
    assign weights1[47][731] = 16'b0000000000000011;
    assign weights1[47][732] = 16'b0000000000001111;
    assign weights1[47][733] = 16'b1111111111110111;
    assign weights1[47][734] = 16'b0000000000011110;
    assign weights1[47][735] = 16'b0000000000000111;
    assign weights1[47][736] = 16'b0000000000011000;
    assign weights1[47][737] = 16'b0000000000100010;
    assign weights1[47][738] = 16'b0000000000101100;
    assign weights1[47][739] = 16'b0000000000110010;
    assign weights1[47][740] = 16'b0000000000010100;
    assign weights1[47][741] = 16'b0000000000010110;
    assign weights1[47][742] = 16'b0000000000010001;
    assign weights1[47][743] = 16'b0000000000010101;
    assign weights1[47][744] = 16'b0000000000001000;
    assign weights1[47][745] = 16'b0000000000001011;
    assign weights1[47][746] = 16'b0000000000010101;
    assign weights1[47][747] = 16'b1111111111110100;
    assign weights1[47][748] = 16'b1111111111110111;
    assign weights1[47][749] = 16'b0000000000001110;
    assign weights1[47][750] = 16'b0000000000011000;
    assign weights1[47][751] = 16'b0000000000000110;
    assign weights1[47][752] = 16'b0000000000000010;
    assign weights1[47][753] = 16'b0000000000000011;
    assign weights1[47][754] = 16'b0000000000000000;
    assign weights1[47][755] = 16'b1111111111111111;
    assign weights1[47][756] = 16'b0000000000000100;
    assign weights1[47][757] = 16'b0000000000000010;
    assign weights1[47][758] = 16'b0000000000000100;
    assign weights1[47][759] = 16'b0000000000010011;
    assign weights1[47][760] = 16'b0000000000011000;
    assign weights1[47][761] = 16'b0000000000010111;
    assign weights1[47][762] = 16'b0000000000101101;
    assign weights1[47][763] = 16'b0000000000101011;
    assign weights1[47][764] = 16'b0000000000100100;
    assign weights1[47][765] = 16'b0000000000101011;
    assign weights1[47][766] = 16'b0000000000100110;
    assign weights1[47][767] = 16'b0000000000010110;
    assign weights1[47][768] = 16'b0000000000011111;
    assign weights1[47][769] = 16'b0000000000011101;
    assign weights1[47][770] = 16'b0000000000011111;
    assign weights1[47][771] = 16'b0000000000011000;
    assign weights1[47][772] = 16'b0000000000001101;
    assign weights1[47][773] = 16'b0000000000011001;
    assign weights1[47][774] = 16'b0000000000001101;
    assign weights1[47][775] = 16'b0000000000000111;
    assign weights1[47][776] = 16'b0000000000001010;
    assign weights1[47][777] = 16'b0000000000011010;
    assign weights1[47][778] = 16'b0000000000010001;
    assign weights1[47][779] = 16'b0000000000001000;
    assign weights1[47][780] = 16'b0000000000000001;
    assign weights1[47][781] = 16'b0000000000000001;
    assign weights1[47][782] = 16'b1111111111111111;
    assign weights1[47][783] = 16'b0000000000000000;
    assign weights1[48][0] = 16'b1111111111111111;
    assign weights1[48][1] = 16'b1111111111111110;
    assign weights1[48][2] = 16'b1111111111111110;
    assign weights1[48][3] = 16'b1111111111111100;
    assign weights1[48][4] = 16'b1111111111111110;
    assign weights1[48][5] = 16'b1111111111111101;
    assign weights1[48][6] = 16'b0000000000000101;
    assign weights1[48][7] = 16'b0000000000010011;
    assign weights1[48][8] = 16'b0000000000000110;
    assign weights1[48][9] = 16'b0000000000000111;
    assign weights1[48][10] = 16'b1111111111111010;
    assign weights1[48][11] = 16'b0000000000000010;
    assign weights1[48][12] = 16'b1111111111111100;
    assign weights1[48][13] = 16'b1111111111111110;
    assign weights1[48][14] = 16'b1111111111111001;
    assign weights1[48][15] = 16'b1111111111111000;
    assign weights1[48][16] = 16'b1111111111101111;
    assign weights1[48][17] = 16'b1111111111110111;
    assign weights1[48][18] = 16'b1111111111111011;
    assign weights1[48][19] = 16'b1111111111111011;
    assign weights1[48][20] = 16'b0000000000000000;
    assign weights1[48][21] = 16'b0000000000000101;
    assign weights1[48][22] = 16'b0000000000000010;
    assign weights1[48][23] = 16'b0000000000000001;
    assign weights1[48][24] = 16'b0000000000000000;
    assign weights1[48][25] = 16'b1111111111111000;
    assign weights1[48][26] = 16'b1111111111111101;
    assign weights1[48][27] = 16'b0000000000000000;
    assign weights1[48][28] = 16'b0000000000000001;
    assign weights1[48][29] = 16'b1111111111111111;
    assign weights1[48][30] = 16'b1111111111111100;
    assign weights1[48][31] = 16'b1111111111111011;
    assign weights1[48][32] = 16'b0000000000000011;
    assign weights1[48][33] = 16'b0000000000000010;
    assign weights1[48][34] = 16'b0000000000000100;
    assign weights1[48][35] = 16'b0000000000001100;
    assign weights1[48][36] = 16'b0000000000010000;
    assign weights1[48][37] = 16'b0000000000001011;
    assign weights1[48][38] = 16'b1111111111110100;
    assign weights1[48][39] = 16'b0000000000000000;
    assign weights1[48][40] = 16'b1111111111111100;
    assign weights1[48][41] = 16'b1111111111100110;
    assign weights1[48][42] = 16'b0000000000000110;
    assign weights1[48][43] = 16'b1111111111111001;
    assign weights1[48][44] = 16'b1111111111101011;
    assign weights1[48][45] = 16'b1111111111110000;
    assign weights1[48][46] = 16'b0000000000000111;
    assign weights1[48][47] = 16'b0000000000000100;
    assign weights1[48][48] = 16'b1111111111111101;
    assign weights1[48][49] = 16'b1111111111111111;
    assign weights1[48][50] = 16'b0000000000001100;
    assign weights1[48][51] = 16'b0000000000001000;
    assign weights1[48][52] = 16'b1111111111110100;
    assign weights1[48][53] = 16'b1111111111110100;
    assign weights1[48][54] = 16'b1111111111111100;
    assign weights1[48][55] = 16'b0000000000000000;
    assign weights1[48][56] = 16'b1111111111111111;
    assign weights1[48][57] = 16'b1111111111111110;
    assign weights1[48][58] = 16'b1111111111111010;
    assign weights1[48][59] = 16'b0000000000001000;
    assign weights1[48][60] = 16'b0000000000000001;
    assign weights1[48][61] = 16'b0000000000000000;
    assign weights1[48][62] = 16'b1111111111111011;
    assign weights1[48][63] = 16'b0000000000001100;
    assign weights1[48][64] = 16'b0000000000000101;
    assign weights1[48][65] = 16'b1111111111111101;
    assign weights1[48][66] = 16'b0000000000000111;
    assign weights1[48][67] = 16'b1111111111111010;
    assign weights1[48][68] = 16'b1111111111111011;
    assign weights1[48][69] = 16'b1111111111100111;
    assign weights1[48][70] = 16'b1111111111101001;
    assign weights1[48][71] = 16'b1111111111110001;
    assign weights1[48][72] = 16'b0000000000000100;
    assign weights1[48][73] = 16'b0000000000000010;
    assign weights1[48][74] = 16'b0000000000001100;
    assign weights1[48][75] = 16'b1111111111101000;
    assign weights1[48][76] = 16'b0000000000001000;
    assign weights1[48][77] = 16'b1111111111111101;
    assign weights1[48][78] = 16'b0000000000000001;
    assign weights1[48][79] = 16'b1111111111111101;
    assign weights1[48][80] = 16'b1111111111110101;
    assign weights1[48][81] = 16'b1111111111110101;
    assign weights1[48][82] = 16'b1111111111111111;
    assign weights1[48][83] = 16'b1111111111111111;
    assign weights1[48][84] = 16'b1111111111111101;
    assign weights1[48][85] = 16'b1111111111111100;
    assign weights1[48][86] = 16'b0000000000000001;
    assign weights1[48][87] = 16'b0000000000000000;
    assign weights1[48][88] = 16'b1111111111111101;
    assign weights1[48][89] = 16'b0000000000001010;
    assign weights1[48][90] = 16'b0000000000000001;
    assign weights1[48][91] = 16'b1111111111110110;
    assign weights1[48][92] = 16'b1111111111110100;
    assign weights1[48][93] = 16'b1111111111111101;
    assign weights1[48][94] = 16'b1111111111011111;
    assign weights1[48][95] = 16'b0000000000000100;
    assign weights1[48][96] = 16'b1111111111110111;
    assign weights1[48][97] = 16'b0000000000000010;
    assign weights1[48][98] = 16'b0000000000010000;
    assign weights1[48][99] = 16'b0000000000000010;
    assign weights1[48][100] = 16'b0000000000001001;
    assign weights1[48][101] = 16'b1111111111111010;
    assign weights1[48][102] = 16'b0000000000010001;
    assign weights1[48][103] = 16'b0000000000001000;
    assign weights1[48][104] = 16'b0000000000010011;
    assign weights1[48][105] = 16'b0000000000001100;
    assign weights1[48][106] = 16'b0000000000000001;
    assign weights1[48][107] = 16'b1111111111111101;
    assign weights1[48][108] = 16'b0000000000000101;
    assign weights1[48][109] = 16'b0000000000001101;
    assign weights1[48][110] = 16'b0000000000001010;
    assign weights1[48][111] = 16'b0000000000000101;
    assign weights1[48][112] = 16'b1111111111111011;
    assign weights1[48][113] = 16'b1111111111111011;
    assign weights1[48][114] = 16'b1111111111111101;
    assign weights1[48][115] = 16'b0000000000000101;
    assign weights1[48][116] = 16'b1111111111111010;
    assign weights1[48][117] = 16'b0000000000001010;
    assign weights1[48][118] = 16'b0000000000001000;
    assign weights1[48][119] = 16'b0000000000000100;
    assign weights1[48][120] = 16'b1111111111111110;
    assign weights1[48][121] = 16'b0000000000000110;
    assign weights1[48][122] = 16'b1111111111111101;
    assign weights1[48][123] = 16'b1111111111111001;
    assign weights1[48][124] = 16'b1111111111111110;
    assign weights1[48][125] = 16'b1111111111111100;
    assign weights1[48][126] = 16'b1111111111101010;
    assign weights1[48][127] = 16'b0000000000000001;
    assign weights1[48][128] = 16'b1111111111111000;
    assign weights1[48][129] = 16'b0000000000000001;
    assign weights1[48][130] = 16'b0000000000001100;
    assign weights1[48][131] = 16'b0000000000001000;
    assign weights1[48][132] = 16'b1111111111101111;
    assign weights1[48][133] = 16'b1111111111111101;
    assign weights1[48][134] = 16'b1111111111110111;
    assign weights1[48][135] = 16'b0000000000001010;
    assign weights1[48][136] = 16'b1111111111110101;
    assign weights1[48][137] = 16'b1111111111111110;
    assign weights1[48][138] = 16'b0000000000000100;
    assign weights1[48][139] = 16'b1111111111111101;
    assign weights1[48][140] = 16'b1111111111111010;
    assign weights1[48][141] = 16'b1111111111110110;
    assign weights1[48][142] = 16'b0000000000001010;
    assign weights1[48][143] = 16'b1111111111110111;
    assign weights1[48][144] = 16'b0000000000000011;
    assign weights1[48][145] = 16'b1111111111110111;
    assign weights1[48][146] = 16'b1111111111100101;
    assign weights1[48][147] = 16'b1111111111111100;
    assign weights1[48][148] = 16'b1111111111101111;
    assign weights1[48][149] = 16'b0000000000010010;
    assign weights1[48][150] = 16'b0000000000100001;
    assign weights1[48][151] = 16'b1111111111111100;
    assign weights1[48][152] = 16'b1111111111101111;
    assign weights1[48][153] = 16'b1111111111110100;
    assign weights1[48][154] = 16'b0000000000000001;
    assign weights1[48][155] = 16'b1111111111100001;
    assign weights1[48][156] = 16'b0000000000000001;
    assign weights1[48][157] = 16'b1111111111110100;
    assign weights1[48][158] = 16'b1111111111111111;
    assign weights1[48][159] = 16'b1111111111111001;
    assign weights1[48][160] = 16'b0000000000001010;
    assign weights1[48][161] = 16'b1111111111111000;
    assign weights1[48][162] = 16'b1111111111111110;
    assign weights1[48][163] = 16'b1111111111110100;
    assign weights1[48][164] = 16'b1111111111100101;
    assign weights1[48][165] = 16'b0000000000010010;
    assign weights1[48][166] = 16'b0000000000000001;
    assign weights1[48][167] = 16'b1111111111111110;
    assign weights1[48][168] = 16'b0000000000000000;
    assign weights1[48][169] = 16'b1111111111111100;
    assign weights1[48][170] = 16'b0000000000001010;
    assign weights1[48][171] = 16'b0000000000000000;
    assign weights1[48][172] = 16'b1111111111111101;
    assign weights1[48][173] = 16'b0000000000000011;
    assign weights1[48][174] = 16'b1111111111111000;
    assign weights1[48][175] = 16'b0000000000001010;
    assign weights1[48][176] = 16'b1111111111110111;
    assign weights1[48][177] = 16'b1111111111100011;
    assign weights1[48][178] = 16'b1111111111111001;
    assign weights1[48][179] = 16'b1111111111011101;
    assign weights1[48][180] = 16'b1111111111111010;
    assign weights1[48][181] = 16'b1111111111110111;
    assign weights1[48][182] = 16'b1111111111111110;
    assign weights1[48][183] = 16'b0000000000001001;
    assign weights1[48][184] = 16'b1111111111110100;
    assign weights1[48][185] = 16'b1111111111111001;
    assign weights1[48][186] = 16'b0000000000000010;
    assign weights1[48][187] = 16'b1111111111111001;
    assign weights1[48][188] = 16'b1111111111111111;
    assign weights1[48][189] = 16'b1111111111111010;
    assign weights1[48][190] = 16'b1111111111111100;
    assign weights1[48][191] = 16'b0000000000001100;
    assign weights1[48][192] = 16'b0000000000000101;
    assign weights1[48][193] = 16'b1111111111111100;
    assign weights1[48][194] = 16'b1111111111111111;
    assign weights1[48][195] = 16'b0000000000000011;
    assign weights1[48][196] = 16'b1111111111110110;
    assign weights1[48][197] = 16'b1111111111110110;
    assign weights1[48][198] = 16'b0000000000001000;
    assign weights1[48][199] = 16'b1111111111110001;
    assign weights1[48][200] = 16'b0000000000010001;
    assign weights1[48][201] = 16'b0000000000001000;
    assign weights1[48][202] = 16'b0000000000000111;
    assign weights1[48][203] = 16'b1111111111101010;
    assign weights1[48][204] = 16'b0000000000000100;
    assign weights1[48][205] = 16'b1111111111110111;
    assign weights1[48][206] = 16'b1111111111111010;
    assign weights1[48][207] = 16'b0000000000001010;
    assign weights1[48][208] = 16'b1111111111110100;
    assign weights1[48][209] = 16'b1111111111111111;
    assign weights1[48][210] = 16'b1111111111111010;
    assign weights1[48][211] = 16'b1111111111110100;
    assign weights1[48][212] = 16'b0000000000000010;
    assign weights1[48][213] = 16'b0000000000000100;
    assign weights1[48][214] = 16'b1111111111110101;
    assign weights1[48][215] = 16'b0000000000000110;
    assign weights1[48][216] = 16'b1111111111110101;
    assign weights1[48][217] = 16'b1111111111110101;
    assign weights1[48][218] = 16'b0000000000001110;
    assign weights1[48][219] = 16'b1111111111111100;
    assign weights1[48][220] = 16'b1111111111110101;
    assign weights1[48][221] = 16'b1111111111101111;
    assign weights1[48][222] = 16'b0000000000000001;
    assign weights1[48][223] = 16'b0000000000000010;
    assign weights1[48][224] = 16'b1111111111111001;
    assign weights1[48][225] = 16'b1111111111110100;
    assign weights1[48][226] = 16'b1111111111110101;
    assign weights1[48][227] = 16'b0000000000000010;
    assign weights1[48][228] = 16'b0000000000001101;
    assign weights1[48][229] = 16'b1111111111111010;
    assign weights1[48][230] = 16'b0000000000000010;
    assign weights1[48][231] = 16'b1111111111111111;
    assign weights1[48][232] = 16'b1111111111110111;
    assign weights1[48][233] = 16'b0000000000010000;
    assign weights1[48][234] = 16'b1111111111110111;
    assign weights1[48][235] = 16'b1111111111101111;
    assign weights1[48][236] = 16'b0000000000001000;
    assign weights1[48][237] = 16'b1111111111110111;
    assign weights1[48][238] = 16'b0000000000010101;
    assign weights1[48][239] = 16'b0000000000001111;
    assign weights1[48][240] = 16'b1111111111111101;
    assign weights1[48][241] = 16'b0000000000000011;
    assign weights1[48][242] = 16'b1111111111110111;
    assign weights1[48][243] = 16'b1111111111111101;
    assign weights1[48][244] = 16'b0000000000001111;
    assign weights1[48][245] = 16'b1111111111010100;
    assign weights1[48][246] = 16'b0000000000000110;
    assign weights1[48][247] = 16'b1111111111111011;
    assign weights1[48][248] = 16'b1111111111101110;
    assign weights1[48][249] = 16'b1111111111110001;
    assign weights1[48][250] = 16'b1111111111111010;
    assign weights1[48][251] = 16'b1111111111111101;
    assign weights1[48][252] = 16'b1111111111111100;
    assign weights1[48][253] = 16'b0000000000000001;
    assign weights1[48][254] = 16'b1111111111111111;
    assign weights1[48][255] = 16'b1111111111111011;
    assign weights1[48][256] = 16'b1111111111110100;
    assign weights1[48][257] = 16'b1111111111111100;
    assign weights1[48][258] = 16'b1111111111111110;
    assign weights1[48][259] = 16'b0000000000000100;
    assign weights1[48][260] = 16'b0000000000000001;
    assign weights1[48][261] = 16'b1111111111111110;
    assign weights1[48][262] = 16'b1111111111111100;
    assign weights1[48][263] = 16'b1111111111111011;
    assign weights1[48][264] = 16'b1111111111110101;
    assign weights1[48][265] = 16'b1111111111111101;
    assign weights1[48][266] = 16'b1111111111100010;
    assign weights1[48][267] = 16'b1111111111111101;
    assign weights1[48][268] = 16'b1111111111111111;
    assign weights1[48][269] = 16'b1111111111101100;
    assign weights1[48][270] = 16'b1111111111111100;
    assign weights1[48][271] = 16'b1111111111110111;
    assign weights1[48][272] = 16'b0000000000000010;
    assign weights1[48][273] = 16'b1111111111101101;
    assign weights1[48][274] = 16'b0000000000010101;
    assign weights1[48][275] = 16'b1111111111110011;
    assign weights1[48][276] = 16'b1111111111111010;
    assign weights1[48][277] = 16'b0000000000000001;
    assign weights1[48][278] = 16'b1111111111101111;
    assign weights1[48][279] = 16'b0000000000000000;
    assign weights1[48][280] = 16'b1111111111111010;
    assign weights1[48][281] = 16'b0000000000011000;
    assign weights1[48][282] = 16'b0000000000000001;
    assign weights1[48][283] = 16'b0000000000000001;
    assign weights1[48][284] = 16'b1111111111110110;
    assign weights1[48][285] = 16'b1111111111110010;
    assign weights1[48][286] = 16'b0000000000000101;
    assign weights1[48][287] = 16'b1111111111110000;
    assign weights1[48][288] = 16'b1111111111111010;
    assign weights1[48][289] = 16'b1111111111110000;
    assign weights1[48][290] = 16'b1111111111111000;
    assign weights1[48][291] = 16'b1111111111110111;
    assign weights1[48][292] = 16'b0000000000001000;
    assign weights1[48][293] = 16'b1111111111111101;
    assign weights1[48][294] = 16'b1111111111111011;
    assign weights1[48][295] = 16'b1111111111101110;
    assign weights1[48][296] = 16'b1111111111111110;
    assign weights1[48][297] = 16'b1111111111111110;
    assign weights1[48][298] = 16'b0000000000000001;
    assign weights1[48][299] = 16'b1111111111101111;
    assign weights1[48][300] = 16'b0000000000000101;
    assign weights1[48][301] = 16'b1111111111111100;
    assign weights1[48][302] = 16'b1111111111101111;
    assign weights1[48][303] = 16'b1111111111101011;
    assign weights1[48][304] = 16'b1111111111101110;
    assign weights1[48][305] = 16'b1111111111010100;
    assign weights1[48][306] = 16'b1111111111110111;
    assign weights1[48][307] = 16'b1111111111101011;
    assign weights1[48][308] = 16'b1111111111110111;
    assign weights1[48][309] = 16'b1111111111111110;
    assign weights1[48][310] = 16'b1111111111110101;
    assign weights1[48][311] = 16'b1111111111111110;
    assign weights1[48][312] = 16'b1111111111111111;
    assign weights1[48][313] = 16'b1111111111101010;
    assign weights1[48][314] = 16'b0000000000000110;
    assign weights1[48][315] = 16'b1111111111111010;
    assign weights1[48][316] = 16'b1111111111111100;
    assign weights1[48][317] = 16'b1111111111101000;
    assign weights1[48][318] = 16'b0000000000000110;
    assign weights1[48][319] = 16'b1111111111110111;
    assign weights1[48][320] = 16'b1111111111111010;
    assign weights1[48][321] = 16'b0000000000000000;
    assign weights1[48][322] = 16'b0000000000000010;
    assign weights1[48][323] = 16'b0000000000000001;
    assign weights1[48][324] = 16'b1111111111101011;
    assign weights1[48][325] = 16'b1111111111111111;
    assign weights1[48][326] = 16'b1111111111101111;
    assign weights1[48][327] = 16'b1111111111111110;
    assign weights1[48][328] = 16'b1111111111011011;
    assign weights1[48][329] = 16'b1111111111100110;
    assign weights1[48][330] = 16'b1111111111100000;
    assign weights1[48][331] = 16'b1111111111011001;
    assign weights1[48][332] = 16'b1111111111001111;
    assign weights1[48][333] = 16'b1111111111101011;
    assign weights1[48][334] = 16'b1111111111110101;
    assign weights1[48][335] = 16'b1111111111100001;
    assign weights1[48][336] = 16'b1111111111110100;
    assign weights1[48][337] = 16'b1111111111111011;
    assign weights1[48][338] = 16'b1111111111101011;
    assign weights1[48][339] = 16'b0000000000000110;
    assign weights1[48][340] = 16'b1111111111101111;
    assign weights1[48][341] = 16'b1111111111111001;
    assign weights1[48][342] = 16'b1111111111111011;
    assign weights1[48][343] = 16'b0000000000000011;
    assign weights1[48][344] = 16'b1111111111111101;
    assign weights1[48][345] = 16'b0000000000001000;
    assign weights1[48][346] = 16'b0000000000000110;
    assign weights1[48][347] = 16'b0000000000001011;
    assign weights1[48][348] = 16'b0000000000010010;
    assign weights1[48][349] = 16'b1111111111111010;
    assign weights1[48][350] = 16'b1111111111111101;
    assign weights1[48][351] = 16'b0000000000000000;
    assign weights1[48][352] = 16'b0000000000000000;
    assign weights1[48][353] = 16'b1111111111101110;
    assign weights1[48][354] = 16'b1111111111101101;
    assign weights1[48][355] = 16'b1111111111110011;
    assign weights1[48][356] = 16'b1111111111110010;
    assign weights1[48][357] = 16'b0000000000000101;
    assign weights1[48][358] = 16'b0000000000000100;
    assign weights1[48][359] = 16'b1111111111110000;
    assign weights1[48][360] = 16'b1111111111101101;
    assign weights1[48][361] = 16'b1111111111100100;
    assign weights1[48][362] = 16'b1111111111101010;
    assign weights1[48][363] = 16'b1111111111101001;
    assign weights1[48][364] = 16'b1111111111110111;
    assign weights1[48][365] = 16'b0000000000001011;
    assign weights1[48][366] = 16'b1111111111101101;
    assign weights1[48][367] = 16'b0000000000000011;
    assign weights1[48][368] = 16'b1111111111110001;
    assign weights1[48][369] = 16'b0000000000000101;
    assign weights1[48][370] = 16'b1111111111111000;
    assign weights1[48][371] = 16'b1111111111111000;
    assign weights1[48][372] = 16'b1111111111110110;
    assign weights1[48][373] = 16'b0000000000000000;
    assign weights1[48][374] = 16'b1111111111111011;
    assign weights1[48][375] = 16'b1111111111110010;
    assign weights1[48][376] = 16'b1111111111111110;
    assign weights1[48][377] = 16'b1111111111111111;
    assign weights1[48][378] = 16'b0000000000000101;
    assign weights1[48][379] = 16'b1111111111111101;
    assign weights1[48][380] = 16'b1111111111101011;
    assign weights1[48][381] = 16'b0000000000001001;
    assign weights1[48][382] = 16'b1111111111110100;
    assign weights1[48][383] = 16'b1111111111100110;
    assign weights1[48][384] = 16'b1111111111110111;
    assign weights1[48][385] = 16'b1111111111101100;
    assign weights1[48][386] = 16'b1111111111011100;
    assign weights1[48][387] = 16'b1111111111110100;
    assign weights1[48][388] = 16'b1111111111110011;
    assign weights1[48][389] = 16'b1111111111101111;
    assign weights1[48][390] = 16'b1111111111101110;
    assign weights1[48][391] = 16'b1111111111101000;
    assign weights1[48][392] = 16'b0000000000000001;
    assign weights1[48][393] = 16'b0000000000000101;
    assign weights1[48][394] = 16'b1111111111110110;
    assign weights1[48][395] = 16'b0000000000000100;
    assign weights1[48][396] = 16'b1111111111101110;
    assign weights1[48][397] = 16'b1111111111110011;
    assign weights1[48][398] = 16'b0000000000000011;
    assign weights1[48][399] = 16'b0000000000000010;
    assign weights1[48][400] = 16'b0000000000000010;
    assign weights1[48][401] = 16'b0000000000000100;
    assign weights1[48][402] = 16'b0000000000000010;
    assign weights1[48][403] = 16'b1111111111110100;
    assign weights1[48][404] = 16'b0000000000000001;
    assign weights1[48][405] = 16'b1111111111110110;
    assign weights1[48][406] = 16'b1111111111110010;
    assign weights1[48][407] = 16'b1111111111111011;
    assign weights1[48][408] = 16'b1111111111110100;
    assign weights1[48][409] = 16'b1111111111110111;
    assign weights1[48][410] = 16'b0000000000010110;
    assign weights1[48][411] = 16'b1111111111110100;
    assign weights1[48][412] = 16'b1111111111101001;
    assign weights1[48][413] = 16'b0000000000001010;
    assign weights1[48][414] = 16'b0000000000000011;
    assign weights1[48][415] = 16'b0000000000000011;
    assign weights1[48][416] = 16'b0000000000001101;
    assign weights1[48][417] = 16'b0000000000000000;
    assign weights1[48][418] = 16'b0000000000000010;
    assign weights1[48][419] = 16'b1111111111111010;
    assign weights1[48][420] = 16'b0000000000000000;
    assign weights1[48][421] = 16'b0000000000001001;
    assign weights1[48][422] = 16'b0000000000000111;
    assign weights1[48][423] = 16'b0000000000000011;
    assign weights1[48][424] = 16'b0000000000000100;
    assign weights1[48][425] = 16'b0000000000001111;
    assign weights1[48][426] = 16'b0000000000000100;
    assign weights1[48][427] = 16'b0000000000000000;
    assign weights1[48][428] = 16'b1111111111111100;
    assign weights1[48][429] = 16'b1111111111101111;
    assign weights1[48][430] = 16'b0000000000000111;
    assign weights1[48][431] = 16'b1111111111101011;
    assign weights1[48][432] = 16'b1111111111110000;
    assign weights1[48][433] = 16'b1111111111100100;
    assign weights1[48][434] = 16'b0000000000000000;
    assign weights1[48][435] = 16'b1111111111110110;
    assign weights1[48][436] = 16'b1111111111110011;
    assign weights1[48][437] = 16'b0000000000001100;
    assign weights1[48][438] = 16'b1111111111101010;
    assign weights1[48][439] = 16'b0000000000001010;
    assign weights1[48][440] = 16'b1111111111111101;
    assign weights1[48][441] = 16'b1111111111111000;
    assign weights1[48][442] = 16'b1111111111101011;
    assign weights1[48][443] = 16'b0000000000010000;
    assign weights1[48][444] = 16'b0000000000001100;
    assign weights1[48][445] = 16'b0000000000011000;
    assign weights1[48][446] = 16'b0000000000001011;
    assign weights1[48][447] = 16'b0000000000001000;
    assign weights1[48][448] = 16'b0000000000000100;
    assign weights1[48][449] = 16'b0000000000000001;
    assign weights1[48][450] = 16'b0000000000000111;
    assign weights1[48][451] = 16'b1111111111101110;
    assign weights1[48][452] = 16'b1111111111111100;
    assign weights1[48][453] = 16'b0000000000010111;
    assign weights1[48][454] = 16'b0000000000000100;
    assign weights1[48][455] = 16'b1111111111110111;
    assign weights1[48][456] = 16'b0000000000000101;
    assign weights1[48][457] = 16'b0000000000001010;
    assign weights1[48][458] = 16'b1111111111111111;
    assign weights1[48][459] = 16'b0000000000000101;
    assign weights1[48][460] = 16'b1111111111110011;
    assign weights1[48][461] = 16'b1111111111111010;
    assign weights1[48][462] = 16'b1111111111111101;
    assign weights1[48][463] = 16'b1111111111111010;
    assign weights1[48][464] = 16'b1111111111110100;
    assign weights1[48][465] = 16'b0000000000000010;
    assign weights1[48][466] = 16'b1111111111110000;
    assign weights1[48][467] = 16'b0000000000001100;
    assign weights1[48][468] = 16'b1111111111111010;
    assign weights1[48][469] = 16'b0000000000000101;
    assign weights1[48][470] = 16'b0000000000010010;
    assign weights1[48][471] = 16'b0000000000010101;
    assign weights1[48][472] = 16'b0000000000111100;
    assign weights1[48][473] = 16'b0000000000100000;
    assign weights1[48][474] = 16'b0000000000001100;
    assign weights1[48][475] = 16'b0000000000000100;
    assign weights1[48][476] = 16'b0000000000000100;
    assign weights1[48][477] = 16'b1111111111111000;
    assign weights1[48][478] = 16'b0000000000000101;
    assign weights1[48][479] = 16'b1111111111111000;
    assign weights1[48][480] = 16'b0000000000000101;
    assign weights1[48][481] = 16'b0000000000010000;
    assign weights1[48][482] = 16'b0000000000000010;
    assign weights1[48][483] = 16'b1111111111100100;
    assign weights1[48][484] = 16'b1111111111111010;
    assign weights1[48][485] = 16'b1111111111100111;
    assign weights1[48][486] = 16'b0000000000000001;
    assign weights1[48][487] = 16'b1111111111111000;
    assign weights1[48][488] = 16'b1111111111110111;
    assign weights1[48][489] = 16'b1111111111111011;
    assign weights1[48][490] = 16'b1111111111011101;
    assign weights1[48][491] = 16'b1111111111110011;
    assign weights1[48][492] = 16'b1111111111010100;
    assign weights1[48][493] = 16'b1111111111100111;
    assign weights1[48][494] = 16'b1111111111111011;
    assign weights1[48][495] = 16'b0000000000000110;
    assign weights1[48][496] = 16'b1111111111111111;
    assign weights1[48][497] = 16'b0000000000011110;
    assign weights1[48][498] = 16'b0000000000101100;
    assign weights1[48][499] = 16'b0000000000001100;
    assign weights1[48][500] = 16'b0000000000011100;
    assign weights1[48][501] = 16'b0000000000110101;
    assign weights1[48][502] = 16'b0000000000100001;
    assign weights1[48][503] = 16'b0000000000001000;
    assign weights1[48][504] = 16'b0000000000001011;
    assign weights1[48][505] = 16'b1111111111111010;
    assign weights1[48][506] = 16'b0000000000000010;
    assign weights1[48][507] = 16'b1111111111111101;
    assign weights1[48][508] = 16'b1111111111111111;
    assign weights1[48][509] = 16'b1111111111110001;
    assign weights1[48][510] = 16'b1111111111011010;
    assign weights1[48][511] = 16'b0000000000000010;
    assign weights1[48][512] = 16'b0000000000001001;
    assign weights1[48][513] = 16'b1111111111101001;
    assign weights1[48][514] = 16'b1111111111110100;
    assign weights1[48][515] = 16'b1111111111101110;
    assign weights1[48][516] = 16'b1111111111110010;
    assign weights1[48][517] = 16'b1111111111101011;
    assign weights1[48][518] = 16'b1111111111100011;
    assign weights1[48][519] = 16'b1111111111101110;
    assign weights1[48][520] = 16'b0000000000000000;
    assign weights1[48][521] = 16'b0000000000000001;
    assign weights1[48][522] = 16'b0000000000000011;
    assign weights1[48][523] = 16'b0000000000101000;
    assign weights1[48][524] = 16'b0000000000010011;
    assign weights1[48][525] = 16'b0000000000100001;
    assign weights1[48][526] = 16'b0000000000011000;
    assign weights1[48][527] = 16'b0000000000100100;
    assign weights1[48][528] = 16'b0000000000100001;
    assign weights1[48][529] = 16'b0000000000110001;
    assign weights1[48][530] = 16'b0000000000010101;
    assign weights1[48][531] = 16'b0000000000000000;
    assign weights1[48][532] = 16'b0000000000011100;
    assign weights1[48][533] = 16'b0000000000010011;
    assign weights1[48][534] = 16'b0000000000000000;
    assign weights1[48][535] = 16'b0000000000001011;
    assign weights1[48][536] = 16'b0000000000000010;
    assign weights1[48][537] = 16'b0000000000000101;
    assign weights1[48][538] = 16'b1111111111101101;
    assign weights1[48][539] = 16'b1111111111100100;
    assign weights1[48][540] = 16'b1111111111110101;
    assign weights1[48][541] = 16'b1111111111100110;
    assign weights1[48][542] = 16'b1111111111111110;
    assign weights1[48][543] = 16'b1111111111111110;
    assign weights1[48][544] = 16'b1111111111111111;
    assign weights1[48][545] = 16'b0000000000001101;
    assign weights1[48][546] = 16'b0000000000010010;
    assign weights1[48][547] = 16'b0000000000010111;
    assign weights1[48][548] = 16'b0000000000011011;
    assign weights1[48][549] = 16'b0000000000100001;
    assign weights1[48][550] = 16'b0000000000011100;
    assign weights1[48][551] = 16'b1111111111110111;
    assign weights1[48][552] = 16'b0000000000110110;
    assign weights1[48][553] = 16'b0000000000100001;
    assign weights1[48][554] = 16'b0000000000011100;
    assign weights1[48][555] = 16'b0000000000100101;
    assign weights1[48][556] = 16'b0000000000100000;
    assign weights1[48][557] = 16'b0000000000001010;
    assign weights1[48][558] = 16'b0000000000000110;
    assign weights1[48][559] = 16'b1111111111111011;
    assign weights1[48][560] = 16'b0000000000101100;
    assign weights1[48][561] = 16'b0000000000011010;
    assign weights1[48][562] = 16'b0000000000011110;
    assign weights1[48][563] = 16'b0000000000101110;
    assign weights1[48][564] = 16'b0000000000011111;
    assign weights1[48][565] = 16'b0000000000011101;
    assign weights1[48][566] = 16'b0000000000001101;
    assign weights1[48][567] = 16'b0000000000001110;
    assign weights1[48][568] = 16'b0000000000011000;
    assign weights1[48][569] = 16'b0000000000011100;
    assign weights1[48][570] = 16'b0000000000010000;
    assign weights1[48][571] = 16'b0000000000010011;
    assign weights1[48][572] = 16'b0000000000101010;
    assign weights1[48][573] = 16'b0000000000100001;
    assign weights1[48][574] = 16'b0000000000111001;
    assign weights1[48][575] = 16'b0000000000110111;
    assign weights1[48][576] = 16'b0000000000101101;
    assign weights1[48][577] = 16'b0000000000101001;
    assign weights1[48][578] = 16'b0000000000100100;
    assign weights1[48][579] = 16'b0000000000110011;
    assign weights1[48][580] = 16'b0000000000011010;
    assign weights1[48][581] = 16'b0000000000011001;
    assign weights1[48][582] = 16'b0000000000010011;
    assign weights1[48][583] = 16'b0000000000010111;
    assign weights1[48][584] = 16'b0000000000010000;
    assign weights1[48][585] = 16'b1111111111110101;
    assign weights1[48][586] = 16'b1111111111101011;
    assign weights1[48][587] = 16'b1111111111011111;
    assign weights1[48][588] = 16'b0000000000101001;
    assign weights1[48][589] = 16'b0000000000101011;
    assign weights1[48][590] = 16'b0000000000011111;
    assign weights1[48][591] = 16'b0000000000110110;
    assign weights1[48][592] = 16'b0000000000100100;
    assign weights1[48][593] = 16'b0000000000011011;
    assign weights1[48][594] = 16'b0000000000011000;
    assign weights1[48][595] = 16'b0000000000110011;
    assign weights1[48][596] = 16'b0000000000011101;
    assign weights1[48][597] = 16'b0000000000110010;
    assign weights1[48][598] = 16'b0000000000110000;
    assign weights1[48][599] = 16'b0000000000100111;
    assign weights1[48][600] = 16'b0000000000110000;
    assign weights1[48][601] = 16'b0000000000111101;
    assign weights1[48][602] = 16'b0000000000010100;
    assign weights1[48][603] = 16'b0000000000100010;
    assign weights1[48][604] = 16'b0000000000100110;
    assign weights1[48][605] = 16'b0000000000001011;
    assign weights1[48][606] = 16'b0000000000100011;
    assign weights1[48][607] = 16'b0000000000100001;
    assign weights1[48][608] = 16'b0000000000011000;
    assign weights1[48][609] = 16'b0000000000100000;
    assign weights1[48][610] = 16'b0000000000010100;
    assign weights1[48][611] = 16'b1111111111111000;
    assign weights1[48][612] = 16'b1111111111110000;
    assign weights1[48][613] = 16'b1111111111001000;
    assign weights1[48][614] = 16'b1111111111001010;
    assign weights1[48][615] = 16'b1111111111011110;
    assign weights1[48][616] = 16'b0000000000010110;
    assign weights1[48][617] = 16'b0000000000010100;
    assign weights1[48][618] = 16'b0000000000010100;
    assign weights1[48][619] = 16'b0000000000101110;
    assign weights1[48][620] = 16'b0000000000100000;
    assign weights1[48][621] = 16'b0000000000110101;
    assign weights1[48][622] = 16'b0000000000110111;
    assign weights1[48][623] = 16'b0000000000000010;
    assign weights1[48][624] = 16'b0000000000011010;
    assign weights1[48][625] = 16'b0000000000011111;
    assign weights1[48][626] = 16'b1111111111111001;
    assign weights1[48][627] = 16'b0000000000011100;
    assign weights1[48][628] = 16'b0000000000011100;
    assign weights1[48][629] = 16'b0000000000001000;
    assign weights1[48][630] = 16'b0000000000000011;
    assign weights1[48][631] = 16'b0000000000101110;
    assign weights1[48][632] = 16'b0000000000011011;
    assign weights1[48][633] = 16'b0000000000011100;
    assign weights1[48][634] = 16'b0000000000011101;
    assign weights1[48][635] = 16'b0000000000110111;
    assign weights1[48][636] = 16'b0000000000001110;
    assign weights1[48][637] = 16'b0000000000011010;
    assign weights1[48][638] = 16'b1111111111011001;
    assign weights1[48][639] = 16'b1111111111100101;
    assign weights1[48][640] = 16'b1111111111010001;
    assign weights1[48][641] = 16'b1111111111001001;
    assign weights1[48][642] = 16'b1111111111001000;
    assign weights1[48][643] = 16'b1111111111010010;
    assign weights1[48][644] = 16'b0000000000010010;
    assign weights1[48][645] = 16'b0000000000000101;
    assign weights1[48][646] = 16'b0000000000001111;
    assign weights1[48][647] = 16'b0000000000010011;
    assign weights1[48][648] = 16'b0000000000010100;
    assign weights1[48][649] = 16'b0000000000011110;
    assign weights1[48][650] = 16'b0000000000100010;
    assign weights1[48][651] = 16'b0000000000010111;
    assign weights1[48][652] = 16'b0000000000011011;
    assign weights1[48][653] = 16'b0000000000010001;
    assign weights1[48][654] = 16'b0000000000011000;
    assign weights1[48][655] = 16'b0000000000010111;
    assign weights1[48][656] = 16'b0000000000100001;
    assign weights1[48][657] = 16'b0000000000011011;
    assign weights1[48][658] = 16'b0000000000011001;
    assign weights1[48][659] = 16'b0000000000011011;
    assign weights1[48][660] = 16'b0000000000000110;
    assign weights1[48][661] = 16'b1111111111110011;
    assign weights1[48][662] = 16'b0000000000000010;
    assign weights1[48][663] = 16'b1111111111111001;
    assign weights1[48][664] = 16'b1111111111101001;
    assign weights1[48][665] = 16'b1111111111001000;
    assign weights1[48][666] = 16'b1111111110100110;
    assign weights1[48][667] = 16'b1111111110110110;
    assign weights1[48][668] = 16'b1111111110110111;
    assign weights1[48][669] = 16'b1111111111001011;
    assign weights1[48][670] = 16'b1111111111000111;
    assign weights1[48][671] = 16'b1111111111011000;
    assign weights1[48][672] = 16'b0000000000000000;
    assign weights1[48][673] = 16'b1111111111111101;
    assign weights1[48][674] = 16'b1111111111111000;
    assign weights1[48][675] = 16'b1111111111100000;
    assign weights1[48][676] = 16'b0000000000000000;
    assign weights1[48][677] = 16'b1111111111111000;
    assign weights1[48][678] = 16'b1111111111111111;
    assign weights1[48][679] = 16'b0000000000000001;
    assign weights1[48][680] = 16'b0000000000001000;
    assign weights1[48][681] = 16'b0000000000001001;
    assign weights1[48][682] = 16'b1111111111101111;
    assign weights1[48][683] = 16'b1111111111110100;
    assign weights1[48][684] = 16'b1111111111111111;
    assign weights1[48][685] = 16'b1111111111101000;
    assign weights1[48][686] = 16'b0000000000001000;
    assign weights1[48][687] = 16'b1111111111010111;
    assign weights1[48][688] = 16'b1111111111101100;
    assign weights1[48][689] = 16'b1111111111101000;
    assign weights1[48][690] = 16'b1111111111010110;
    assign weights1[48][691] = 16'b1111111110001100;
    assign weights1[48][692] = 16'b1111111101101100;
    assign weights1[48][693] = 16'b1111111101111100;
    assign weights1[48][694] = 16'b1111111101111110;
    assign weights1[48][695] = 16'b1111111110011001;
    assign weights1[48][696] = 16'b1111111110110100;
    assign weights1[48][697] = 16'b1111111111001110;
    assign weights1[48][698] = 16'b1111111111011001;
    assign weights1[48][699] = 16'b1111111111011000;
    assign weights1[48][700] = 16'b1111111111111110;
    assign weights1[48][701] = 16'b1111111111110101;
    assign weights1[48][702] = 16'b1111111111100001;
    assign weights1[48][703] = 16'b1111111111010011;
    assign weights1[48][704] = 16'b1111111111000110;
    assign weights1[48][705] = 16'b1111111111001111;
    assign weights1[48][706] = 16'b1111111111010001;
    assign weights1[48][707] = 16'b1111111111011001;
    assign weights1[48][708] = 16'b1111111111011000;
    assign weights1[48][709] = 16'b1111111111010111;
    assign weights1[48][710] = 16'b1111111111010110;
    assign weights1[48][711] = 16'b1111111110111001;
    assign weights1[48][712] = 16'b1111111110101001;
    assign weights1[48][713] = 16'b1111111110101001;
    assign weights1[48][714] = 16'b1111111101101011;
    assign weights1[48][715] = 16'b1111111101110101;
    assign weights1[48][716] = 16'b1111111101011001;
    assign weights1[48][717] = 16'b1111111101010001;
    assign weights1[48][718] = 16'b1111111101001100;
    assign weights1[48][719] = 16'b1111111101101011;
    assign weights1[48][720] = 16'b1111111101110011;
    assign weights1[48][721] = 16'b1111111110000101;
    assign weights1[48][722] = 16'b1111111110011010;
    assign weights1[48][723] = 16'b1111111110101010;
    assign weights1[48][724] = 16'b1111111110110001;
    assign weights1[48][725] = 16'b1111111111010001;
    assign weights1[48][726] = 16'b1111111111011101;
    assign weights1[48][727] = 16'b1111111111100110;
    assign weights1[48][728] = 16'b1111111111111001;
    assign weights1[48][729] = 16'b1111111111110110;
    assign weights1[48][730] = 16'b1111111111011011;
    assign weights1[48][731] = 16'b1111111111010110;
    assign weights1[48][732] = 16'b1111111111001010;
    assign weights1[48][733] = 16'b1111111110110010;
    assign weights1[48][734] = 16'b1111111110101011;
    assign weights1[48][735] = 16'b1111111110100000;
    assign weights1[48][736] = 16'b1111111110010011;
    assign weights1[48][737] = 16'b1111111110000101;
    assign weights1[48][738] = 16'b1111111110000001;
    assign weights1[48][739] = 16'b1111111101101010;
    assign weights1[48][740] = 16'b1111111101110101;
    assign weights1[48][741] = 16'b1111111101101000;
    assign weights1[48][742] = 16'b1111111101110001;
    assign weights1[48][743] = 16'b1111111101101001;
    assign weights1[48][744] = 16'b1111111101101110;
    assign weights1[48][745] = 16'b1111111101110010;
    assign weights1[48][746] = 16'b1111111101111011;
    assign weights1[48][747] = 16'b1111111110000111;
    assign weights1[48][748] = 16'b1111111110100000;
    assign weights1[48][749] = 16'b1111111110110000;
    assign weights1[48][750] = 16'b1111111111000110;
    assign weights1[48][751] = 16'b1111111111000010;
    assign weights1[48][752] = 16'b1111111111000111;
    assign weights1[48][753] = 16'b1111111111011101;
    assign weights1[48][754] = 16'b1111111111100110;
    assign weights1[48][755] = 16'b1111111111110101;
    assign weights1[48][756] = 16'b1111111111111100;
    assign weights1[48][757] = 16'b1111111111111100;
    assign weights1[48][758] = 16'b1111111111110000;
    assign weights1[48][759] = 16'b1111111111101000;
    assign weights1[48][760] = 16'b1111111111011001;
    assign weights1[48][761] = 16'b1111111111001100;
    assign weights1[48][762] = 16'b1111111111001011;
    assign weights1[48][763] = 16'b1111111110111100;
    assign weights1[48][764] = 16'b1111111110111001;
    assign weights1[48][765] = 16'b1111111110101010;
    assign weights1[48][766] = 16'b1111111110100110;
    assign weights1[48][767] = 16'b1111111110100000;
    assign weights1[48][768] = 16'b1111111110100100;
    assign weights1[48][769] = 16'b1111111110100001;
    assign weights1[48][770] = 16'b1111111110011101;
    assign weights1[48][771] = 16'b1111111110100100;
    assign weights1[48][772] = 16'b1111111110011100;
    assign weights1[48][773] = 16'b1111111110100111;
    assign weights1[48][774] = 16'b1111111110101110;
    assign weights1[48][775] = 16'b1111111110110110;
    assign weights1[48][776] = 16'b1111111111000100;
    assign weights1[48][777] = 16'b1111111111001111;
    assign weights1[48][778] = 16'b1111111111011110;
    assign weights1[48][779] = 16'b1111111111100010;
    assign weights1[48][780] = 16'b1111111111011010;
    assign weights1[48][781] = 16'b1111111111101101;
    assign weights1[48][782] = 16'b1111111111110000;
    assign weights1[48][783] = 16'b1111111111111101;
    assign weights1[49][0] = 16'b0000000000000000;
    assign weights1[49][1] = 16'b0000000000000001;
    assign weights1[49][2] = 16'b0000000000000000;
    assign weights1[49][3] = 16'b0000000000000000;
    assign weights1[49][4] = 16'b1111111111111111;
    assign weights1[49][5] = 16'b1111111111111110;
    assign weights1[49][6] = 16'b1111111111111101;
    assign weights1[49][7] = 16'b1111111111111010;
    assign weights1[49][8] = 16'b1111111111111011;
    assign weights1[49][9] = 16'b1111111111111111;
    assign weights1[49][10] = 16'b1111111111111101;
    assign weights1[49][11] = 16'b1111111111111110;
    assign weights1[49][12] = 16'b1111111111111011;
    assign weights1[49][13] = 16'b1111111111110101;
    assign weights1[49][14] = 16'b1111111111110001;
    assign weights1[49][15] = 16'b1111111111111101;
    assign weights1[49][16] = 16'b1111111111111001;
    assign weights1[49][17] = 16'b0000000000001011;
    assign weights1[49][18] = 16'b0000000000000011;
    assign weights1[49][19] = 16'b1111111111111000;
    assign weights1[49][20] = 16'b1111111111110110;
    assign weights1[49][21] = 16'b1111111111111111;
    assign weights1[49][22] = 16'b1111111111111010;
    assign weights1[49][23] = 16'b1111111111111101;
    assign weights1[49][24] = 16'b1111111111111111;
    assign weights1[49][25] = 16'b0000000000000011;
    assign weights1[49][26] = 16'b0000000000000010;
    assign weights1[49][27] = 16'b0000000000000000;
    assign weights1[49][28] = 16'b0000000000000000;
    assign weights1[49][29] = 16'b0000000000000001;
    assign weights1[49][30] = 16'b0000000000000100;
    assign weights1[49][31] = 16'b0000000000000110;
    assign weights1[49][32] = 16'b0000000000000010;
    assign weights1[49][33] = 16'b0000000000000111;
    assign weights1[49][34] = 16'b0000000000001010;
    assign weights1[49][35] = 16'b0000000000000110;
    assign weights1[49][36] = 16'b0000000000001001;
    assign weights1[49][37] = 16'b0000000000001100;
    assign weights1[49][38] = 16'b0000000000000000;
    assign weights1[49][39] = 16'b1111111111101001;
    assign weights1[49][40] = 16'b1111111111110101;
    assign weights1[49][41] = 16'b1111111111110111;
    assign weights1[49][42] = 16'b1111111111100111;
    assign weights1[49][43] = 16'b0000000000001101;
    assign weights1[49][44] = 16'b0000000000001110;
    assign weights1[49][45] = 16'b0000000000001011;
    assign weights1[49][46] = 16'b1111111111111111;
    assign weights1[49][47] = 16'b1111111111111000;
    assign weights1[49][48] = 16'b1111111111111001;
    assign weights1[49][49] = 16'b0000000000000001;
    assign weights1[49][50] = 16'b0000000000000000;
    assign weights1[49][51] = 16'b0000000000000100;
    assign weights1[49][52] = 16'b0000000000000010;
    assign weights1[49][53] = 16'b0000000000000011;
    assign weights1[49][54] = 16'b0000000000000001;
    assign weights1[49][55] = 16'b1111111111111111;
    assign weights1[49][56] = 16'b0000000000000000;
    assign weights1[49][57] = 16'b0000000000000010;
    assign weights1[49][58] = 16'b0000000000001010;
    assign weights1[49][59] = 16'b0000000000001100;
    assign weights1[49][60] = 16'b0000000000001110;
    assign weights1[49][61] = 16'b0000000000010001;
    assign weights1[49][62] = 16'b0000000000010001;
    assign weights1[49][63] = 16'b0000000000010101;
    assign weights1[49][64] = 16'b0000000000001000;
    assign weights1[49][65] = 16'b0000000000001011;
    assign weights1[49][66] = 16'b1111111111111110;
    assign weights1[49][67] = 16'b1111111111101110;
    assign weights1[49][68] = 16'b0000000000000010;
    assign weights1[49][69] = 16'b0000000000000000;
    assign weights1[49][70] = 16'b1111111111110100;
    assign weights1[49][71] = 16'b1111111111101110;
    assign weights1[49][72] = 16'b1111111111110001;
    assign weights1[49][73] = 16'b1111111111110000;
    assign weights1[49][74] = 16'b1111111111110110;
    assign weights1[49][75] = 16'b0000000000000001;
    assign weights1[49][76] = 16'b1111111111111101;
    assign weights1[49][77] = 16'b1111111111111101;
    assign weights1[49][78] = 16'b1111111111111101;
    assign weights1[49][79] = 16'b0000000000000011;
    assign weights1[49][80] = 16'b0000000000000010;
    assign weights1[49][81] = 16'b0000000000000101;
    assign weights1[49][82] = 16'b0000000000000101;
    assign weights1[49][83] = 16'b0000000000000100;
    assign weights1[49][84] = 16'b0000000000000001;
    assign weights1[49][85] = 16'b0000000000000100;
    assign weights1[49][86] = 16'b0000000000001110;
    assign weights1[49][87] = 16'b0000000000010100;
    assign weights1[49][88] = 16'b0000000000011100;
    assign weights1[49][89] = 16'b0000000000100001;
    assign weights1[49][90] = 16'b0000000000011001;
    assign weights1[49][91] = 16'b0000000000001010;
    assign weights1[49][92] = 16'b0000000000011001;
    assign weights1[49][93] = 16'b0000000000010110;
    assign weights1[49][94] = 16'b0000000000010000;
    assign weights1[49][95] = 16'b0000000000000000;
    assign weights1[49][96] = 16'b1111111111101111;
    assign weights1[49][97] = 16'b1111111111111111;
    assign weights1[49][98] = 16'b1111111111111101;
    assign weights1[49][99] = 16'b1111111111110100;
    assign weights1[49][100] = 16'b1111111111110100;
    assign weights1[49][101] = 16'b1111111111100111;
    assign weights1[49][102] = 16'b1111111111011000;
    assign weights1[49][103] = 16'b1111111111100101;
    assign weights1[49][104] = 16'b1111111111011010;
    assign weights1[49][105] = 16'b1111111111110101;
    assign weights1[49][106] = 16'b1111111111111011;
    assign weights1[49][107] = 16'b0000000000000000;
    assign weights1[49][108] = 16'b0000000000000100;
    assign weights1[49][109] = 16'b0000000000000011;
    assign weights1[49][110] = 16'b0000000000001000;
    assign weights1[49][111] = 16'b0000000000000011;
    assign weights1[49][112] = 16'b0000000000000110;
    assign weights1[49][113] = 16'b0000000000001000;
    assign weights1[49][114] = 16'b0000000000010011;
    assign weights1[49][115] = 16'b0000000000011110;
    assign weights1[49][116] = 16'b0000000000011011;
    assign weights1[49][117] = 16'b0000000000011000;
    assign weights1[49][118] = 16'b0000000000011101;
    assign weights1[49][119] = 16'b0000000000011000;
    assign weights1[49][120] = 16'b0000000000001000;
    assign weights1[49][121] = 16'b0000000000011001;
    assign weights1[49][122] = 16'b1111111111111101;
    assign weights1[49][123] = 16'b0000000000001011;
    assign weights1[49][124] = 16'b1111111111110101;
    assign weights1[49][125] = 16'b1111111111111111;
    assign weights1[49][126] = 16'b1111111111111111;
    assign weights1[49][127] = 16'b1111111111111000;
    assign weights1[49][128] = 16'b0000000000010010;
    assign weights1[49][129] = 16'b0000000000000101;
    assign weights1[49][130] = 16'b0000000000010001;
    assign weights1[49][131] = 16'b1111111111111001;
    assign weights1[49][132] = 16'b1111111111110001;
    assign weights1[49][133] = 16'b1111111111101111;
    assign weights1[49][134] = 16'b1111111111111001;
    assign weights1[49][135] = 16'b0000000000000001;
    assign weights1[49][136] = 16'b0000000000001010;
    assign weights1[49][137] = 16'b0000000000000100;
    assign weights1[49][138] = 16'b0000000000001011;
    assign weights1[49][139] = 16'b0000000000001101;
    assign weights1[49][140] = 16'b0000000000000111;
    assign weights1[49][141] = 16'b0000000000010001;
    assign weights1[49][142] = 16'b0000000000010001;
    assign weights1[49][143] = 16'b0000000000011010;
    assign weights1[49][144] = 16'b0000000000010011;
    assign weights1[49][145] = 16'b0000000000001001;
    assign weights1[49][146] = 16'b0000000000001110;
    assign weights1[49][147] = 16'b0000000000010100;
    assign weights1[49][148] = 16'b0000000000000011;
    assign weights1[49][149] = 16'b0000000000010000;
    assign weights1[49][150] = 16'b1111111111111110;
    assign weights1[49][151] = 16'b0000000000001001;
    assign weights1[49][152] = 16'b1111111111101100;
    assign weights1[49][153] = 16'b0000000000001011;
    assign weights1[49][154] = 16'b1111111111100101;
    assign weights1[49][155] = 16'b1111111111110111;
    assign weights1[49][156] = 16'b1111111111110010;
    assign weights1[49][157] = 16'b1111111111110101;
    assign weights1[49][158] = 16'b1111111111111010;
    assign weights1[49][159] = 16'b1111111111111110;
    assign weights1[49][160] = 16'b1111111111110110;
    assign weights1[49][161] = 16'b0000000000000010;
    assign weights1[49][162] = 16'b0000000000001001;
    assign weights1[49][163] = 16'b0000000000000111;
    assign weights1[49][164] = 16'b0000000000001010;
    assign weights1[49][165] = 16'b0000000000000001;
    assign weights1[49][166] = 16'b0000000000001101;
    assign weights1[49][167] = 16'b0000000000000100;
    assign weights1[49][168] = 16'b0000000000001001;
    assign weights1[49][169] = 16'b0000000000001111;
    assign weights1[49][170] = 16'b0000000000010011;
    assign weights1[49][171] = 16'b0000000000010100;
    assign weights1[49][172] = 16'b0000000000001010;
    assign weights1[49][173] = 16'b0000000000010010;
    assign weights1[49][174] = 16'b1111111111111110;
    assign weights1[49][175] = 16'b0000000000010100;
    assign weights1[49][176] = 16'b1111111111111001;
    assign weights1[49][177] = 16'b1111111111111001;
    assign weights1[49][178] = 16'b0000000000001000;
    assign weights1[49][179] = 16'b1111111111111010;
    assign weights1[49][180] = 16'b1111111111110101;
    assign weights1[49][181] = 16'b1111111111110001;
    assign weights1[49][182] = 16'b0000000000000000;
    assign weights1[49][183] = 16'b1111111111110110;
    assign weights1[49][184] = 16'b1111111111111010;
    assign weights1[49][185] = 16'b0000000000000101;
    assign weights1[49][186] = 16'b0000000000001101;
    assign weights1[49][187] = 16'b1111111111101010;
    assign weights1[49][188] = 16'b0000000000011100;
    assign weights1[49][189] = 16'b0000000000011101;
    assign weights1[49][190] = 16'b0000000000000110;
    assign weights1[49][191] = 16'b0000000000000110;
    assign weights1[49][192] = 16'b0000000000001001;
    assign weights1[49][193] = 16'b0000000000001110;
    assign weights1[49][194] = 16'b0000000000001101;
    assign weights1[49][195] = 16'b1111111111111101;
    assign weights1[49][196] = 16'b0000000000001010;
    assign weights1[49][197] = 16'b0000000000010001;
    assign weights1[49][198] = 16'b0000000000001000;
    assign weights1[49][199] = 16'b0000000000001000;
    assign weights1[49][200] = 16'b0000000000000011;
    assign weights1[49][201] = 16'b0000000000000000;
    assign weights1[49][202] = 16'b1111111111111110;
    assign weights1[49][203] = 16'b1111111111111111;
    assign weights1[49][204] = 16'b0000000000000101;
    assign weights1[49][205] = 16'b0000000000000100;
    assign weights1[49][206] = 16'b1111111111110101;
    assign weights1[49][207] = 16'b1111111111111001;
    assign weights1[49][208] = 16'b1111111111101010;
    assign weights1[49][209] = 16'b0000000000010000;
    assign weights1[49][210] = 16'b1111111111111011;
    assign weights1[49][211] = 16'b1111111111110101;
    assign weights1[49][212] = 16'b0000000000001111;
    assign weights1[49][213] = 16'b0000000000000101;
    assign weights1[49][214] = 16'b0000000000000010;
    assign weights1[49][215] = 16'b0000000000001011;
    assign weights1[49][216] = 16'b0000000000011010;
    assign weights1[49][217] = 16'b0000000000000010;
    assign weights1[49][218] = 16'b0000000000001010;
    assign weights1[49][219] = 16'b1111111111111010;
    assign weights1[49][220] = 16'b1111111111110100;
    assign weights1[49][221] = 16'b1111111111101111;
    assign weights1[49][222] = 16'b0000000000001100;
    assign weights1[49][223] = 16'b1111111111110101;
    assign weights1[49][224] = 16'b0000000000001000;
    assign weights1[49][225] = 16'b0000000000000111;
    assign weights1[49][226] = 16'b0000000000000101;
    assign weights1[49][227] = 16'b0000000000001001;
    assign weights1[49][228] = 16'b0000000000000001;
    assign weights1[49][229] = 16'b0000000000001100;
    assign weights1[49][230] = 16'b1111111111111110;
    assign weights1[49][231] = 16'b1111111111111010;
    assign weights1[49][232] = 16'b1111111111101111;
    assign weights1[49][233] = 16'b1111111111100010;
    assign weights1[49][234] = 16'b1111111111010101;
    assign weights1[49][235] = 16'b1111111111101111;
    assign weights1[49][236] = 16'b1111111111111001;
    assign weights1[49][237] = 16'b1111111111111000;
    assign weights1[49][238] = 16'b1111111111110010;
    assign weights1[49][239] = 16'b0000000000100000;
    assign weights1[49][240] = 16'b1111111111110010;
    assign weights1[49][241] = 16'b0000000000001111;
    assign weights1[49][242] = 16'b1111111111110111;
    assign weights1[49][243] = 16'b0000000000000100;
    assign weights1[49][244] = 16'b1111111111111001;
    assign weights1[49][245] = 16'b1111111111111110;
    assign weights1[49][246] = 16'b0000000000011011;
    assign weights1[49][247] = 16'b1111111111111101;
    assign weights1[49][248] = 16'b1111111111010110;
    assign weights1[49][249] = 16'b0000000000001000;
    assign weights1[49][250] = 16'b1111111111111000;
    assign weights1[49][251] = 16'b1111111111110001;
    assign weights1[49][252] = 16'b0000000000000011;
    assign weights1[49][253] = 16'b0000000000000100;
    assign weights1[49][254] = 16'b0000000000000011;
    assign weights1[49][255] = 16'b0000000000000001;
    assign weights1[49][256] = 16'b1111111111110111;
    assign weights1[49][257] = 16'b1111111111110100;
    assign weights1[49][258] = 16'b1111111111110001;
    assign weights1[49][259] = 16'b1111111111100011;
    assign weights1[49][260] = 16'b1111111111001001;
    assign weights1[49][261] = 16'b1111111111000111;
    assign weights1[49][262] = 16'b1111111111000000;
    assign weights1[49][263] = 16'b1111111111100111;
    assign weights1[49][264] = 16'b1111111111101000;
    assign weights1[49][265] = 16'b1111111111101010;
    assign weights1[49][266] = 16'b0000000000000001;
    assign weights1[49][267] = 16'b0000000000000101;
    assign weights1[49][268] = 16'b0000000000001011;
    assign weights1[49][269] = 16'b0000000000000111;
    assign weights1[49][270] = 16'b0000000000000111;
    assign weights1[49][271] = 16'b0000000000000010;
    assign weights1[49][272] = 16'b1111111111111100;
    assign weights1[49][273] = 16'b0000000000000101;
    assign weights1[49][274] = 16'b1111111111111011;
    assign weights1[49][275] = 16'b1111111111100001;
    assign weights1[49][276] = 16'b0000000000001001;
    assign weights1[49][277] = 16'b1111111111111011;
    assign weights1[49][278] = 16'b1111111111111001;
    assign weights1[49][279] = 16'b1111111111111101;
    assign weights1[49][280] = 16'b0000000000000100;
    assign weights1[49][281] = 16'b1111111111111110;
    assign weights1[49][282] = 16'b0000000000000010;
    assign weights1[49][283] = 16'b0000000000000001;
    assign weights1[49][284] = 16'b1111111111111111;
    assign weights1[49][285] = 16'b1111111111110001;
    assign weights1[49][286] = 16'b1111111111101001;
    assign weights1[49][287] = 16'b1111111111001000;
    assign weights1[49][288] = 16'b1111111110110101;
    assign weights1[49][289] = 16'b1111111111001011;
    assign weights1[49][290] = 16'b1111111111000001;
    assign weights1[49][291] = 16'b1111111111101011;
    assign weights1[49][292] = 16'b1111111111100110;
    assign weights1[49][293] = 16'b1111111111101111;
    assign weights1[49][294] = 16'b0000000000000111;
    assign weights1[49][295] = 16'b0000000000001001;
    assign weights1[49][296] = 16'b1111111111110101;
    assign weights1[49][297] = 16'b1111111111111001;
    assign weights1[49][298] = 16'b0000000000000011;
    assign weights1[49][299] = 16'b0000000000000110;
    assign weights1[49][300] = 16'b0000000000010000;
    assign weights1[49][301] = 16'b0000000000001100;
    assign weights1[49][302] = 16'b1111111111111101;
    assign weights1[49][303] = 16'b0000000000000100;
    assign weights1[49][304] = 16'b1111111111111011;
    assign weights1[49][305] = 16'b0000000000000101;
    assign weights1[49][306] = 16'b0000000000001100;
    assign weights1[49][307] = 16'b0000000000001001;
    assign weights1[49][308] = 16'b0000000000000101;
    assign weights1[49][309] = 16'b1111111111111111;
    assign weights1[49][310] = 16'b0000000000000011;
    assign weights1[49][311] = 16'b1111111111111101;
    assign weights1[49][312] = 16'b1111111111110101;
    assign weights1[49][313] = 16'b1111111111101011;
    assign weights1[49][314] = 16'b1111111111011011;
    assign weights1[49][315] = 16'b1111111111010001;
    assign weights1[49][316] = 16'b1111111111000101;
    assign weights1[49][317] = 16'b1111111111001111;
    assign weights1[49][318] = 16'b1111111111100001;
    assign weights1[49][319] = 16'b0000000000000001;
    assign weights1[49][320] = 16'b0000000000001000;
    assign weights1[49][321] = 16'b0000000000000101;
    assign weights1[49][322] = 16'b0000000000000101;
    assign weights1[49][323] = 16'b0000000000000101;
    assign weights1[49][324] = 16'b0000000000000111;
    assign weights1[49][325] = 16'b1111111111101100;
    assign weights1[49][326] = 16'b0000000000000101;
    assign weights1[49][327] = 16'b1111111111110101;
    assign weights1[49][328] = 16'b1111111111110111;
    assign weights1[49][329] = 16'b0000000000001101;
    assign weights1[49][330] = 16'b0000000000001100;
    assign weights1[49][331] = 16'b0000000000011011;
    assign weights1[49][332] = 16'b0000000000000110;
    assign weights1[49][333] = 16'b0000000000001001;
    assign weights1[49][334] = 16'b0000000000011001;
    assign weights1[49][335] = 16'b0000000000001000;
    assign weights1[49][336] = 16'b0000000000000000;
    assign weights1[49][337] = 16'b1111111111111100;
    assign weights1[49][338] = 16'b0000000000000000;
    assign weights1[49][339] = 16'b1111111111110001;
    assign weights1[49][340] = 16'b1111111111011111;
    assign weights1[49][341] = 16'b1111111111010101;
    assign weights1[49][342] = 16'b1111111111001000;
    assign weights1[49][343] = 16'b1111111110110110;
    assign weights1[49][344] = 16'b1111111111000001;
    assign weights1[49][345] = 16'b1111111111010100;
    assign weights1[49][346] = 16'b1111111111110100;
    assign weights1[49][347] = 16'b1111111111111011;
    assign weights1[49][348] = 16'b0000000000000101;
    assign weights1[49][349] = 16'b1111111111111011;
    assign weights1[49][350] = 16'b0000000000001101;
    assign weights1[49][351] = 16'b0000000000001111;
    assign weights1[49][352] = 16'b1111111111110110;
    assign weights1[49][353] = 16'b1111111111101100;
    assign weights1[49][354] = 16'b0000000000001000;
    assign weights1[49][355] = 16'b0000000000000110;
    assign weights1[49][356] = 16'b0000000000010000;
    assign weights1[49][357] = 16'b0000000000100010;
    assign weights1[49][358] = 16'b0000000000001000;
    assign weights1[49][359] = 16'b0000000000010000;
    assign weights1[49][360] = 16'b0000000000000010;
    assign weights1[49][361] = 16'b1111111111111010;
    assign weights1[49][362] = 16'b0000000000000011;
    assign weights1[49][363] = 16'b0000000000001101;
    assign weights1[49][364] = 16'b0000000000000000;
    assign weights1[49][365] = 16'b1111111111111101;
    assign weights1[49][366] = 16'b1111111111110000;
    assign weights1[49][367] = 16'b1111111111100100;
    assign weights1[49][368] = 16'b1111111111010010;
    assign weights1[49][369] = 16'b1111111111001001;
    assign weights1[49][370] = 16'b1111111111000000;
    assign weights1[49][371] = 16'b1111111111010100;
    assign weights1[49][372] = 16'b1111111111000011;
    assign weights1[49][373] = 16'b1111111111000100;
    assign weights1[49][374] = 16'b0000000000001000;
    assign weights1[49][375] = 16'b0000000000000011;
    assign weights1[49][376] = 16'b0000000000011000;
    assign weights1[49][377] = 16'b0000000000011001;
    assign weights1[49][378] = 16'b0000000000001111;
    assign weights1[49][379] = 16'b1111111111101000;
    assign weights1[49][380] = 16'b1111111111010110;
    assign weights1[49][381] = 16'b1111111111010100;
    assign weights1[49][382] = 16'b1111111111110001;
    assign weights1[49][383] = 16'b0000000000000010;
    assign weights1[49][384] = 16'b0000000000001111;
    assign weights1[49][385] = 16'b1111111111111110;
    assign weights1[49][386] = 16'b1111111111110010;
    assign weights1[49][387] = 16'b0000000000000110;
    assign weights1[49][388] = 16'b0000000000010101;
    assign weights1[49][389] = 16'b0000000000000001;
    assign weights1[49][390] = 16'b0000000000000100;
    assign weights1[49][391] = 16'b0000000000001001;
    assign weights1[49][392] = 16'b1111111111111100;
    assign weights1[49][393] = 16'b0000000000000001;
    assign weights1[49][394] = 16'b1111111111101001;
    assign weights1[49][395] = 16'b1111111111011101;
    assign weights1[49][396] = 16'b1111111111001111;
    assign weights1[49][397] = 16'b1111111111000101;
    assign weights1[49][398] = 16'b1111111111000101;
    assign weights1[49][399] = 16'b1111111111010011;
    assign weights1[49][400] = 16'b1111111111010001;
    assign weights1[49][401] = 16'b1111111111101111;
    assign weights1[49][402] = 16'b0000000000001110;
    assign weights1[49][403] = 16'b0000000000100001;
    assign weights1[49][404] = 16'b0000000000011011;
    assign weights1[49][405] = 16'b0000000000010111;
    assign weights1[49][406] = 16'b0000000000000111;
    assign weights1[49][407] = 16'b1111111111101100;
    assign weights1[49][408] = 16'b1111111110111001;
    assign weights1[49][409] = 16'b1111111110100101;
    assign weights1[49][410] = 16'b1111111111000100;
    assign weights1[49][411] = 16'b0000000000010010;
    assign weights1[49][412] = 16'b1111111111101110;
    assign weights1[49][413] = 16'b0000000000000010;
    assign weights1[49][414] = 16'b0000000000000101;
    assign weights1[49][415] = 16'b0000000000000011;
    assign weights1[49][416] = 16'b1111111111111001;
    assign weights1[49][417] = 16'b0000000000000101;
    assign weights1[49][418] = 16'b0000000000000011;
    assign weights1[49][419] = 16'b1111111111111101;
    assign weights1[49][420] = 16'b1111111111111000;
    assign weights1[49][421] = 16'b1111111111111010;
    assign weights1[49][422] = 16'b1111111111100101;
    assign weights1[49][423] = 16'b1111111111100010;
    assign weights1[49][424] = 16'b1111111111011010;
    assign weights1[49][425] = 16'b1111111111010100;
    assign weights1[49][426] = 16'b1111111111001100;
    assign weights1[49][427] = 16'b1111111111100000;
    assign weights1[49][428] = 16'b1111111111101110;
    assign weights1[49][429] = 16'b1111111111101011;
    assign weights1[49][430] = 16'b0000000000011011;
    assign weights1[49][431] = 16'b0000000000001111;
    assign weights1[49][432] = 16'b0000000000010111;
    assign weights1[49][433] = 16'b0000000000010101;
    assign weights1[49][434] = 16'b0000000000000110;
    assign weights1[49][435] = 16'b0000000000010001;
    assign weights1[49][436] = 16'b1111111110110000;
    assign weights1[49][437] = 16'b1111111101111111;
    assign weights1[49][438] = 16'b1111111111000101;
    assign weights1[49][439] = 16'b1111111111110010;
    assign weights1[49][440] = 16'b1111111111111010;
    assign weights1[49][441] = 16'b1111111111111111;
    assign weights1[49][442] = 16'b1111111111110110;
    assign weights1[49][443] = 16'b1111111111111100;
    assign weights1[49][444] = 16'b0000000000000010;
    assign weights1[49][445] = 16'b0000000000001101;
    assign weights1[49][446] = 16'b1111111111111110;
    assign weights1[49][447] = 16'b0000000000001010;
    assign weights1[49][448] = 16'b1111111111111010;
    assign weights1[49][449] = 16'b1111111111110011;
    assign weights1[49][450] = 16'b1111111111101110;
    assign weights1[49][451] = 16'b1111111111101011;
    assign weights1[49][452] = 16'b1111111111100000;
    assign weights1[49][453] = 16'b1111111111100111;
    assign weights1[49][454] = 16'b1111111111100000;
    assign weights1[49][455] = 16'b1111111111101111;
    assign weights1[49][456] = 16'b1111111111100011;
    assign weights1[49][457] = 16'b0000000000001010;
    assign weights1[49][458] = 16'b0000000000010100;
    assign weights1[49][459] = 16'b0000000000010000;
    assign weights1[49][460] = 16'b0000000000111101;
    assign weights1[49][461] = 16'b0000000000101010;
    assign weights1[49][462] = 16'b1111111111111111;
    assign weights1[49][463] = 16'b1111111111100101;
    assign weights1[49][464] = 16'b1111111101110100;
    assign weights1[49][465] = 16'b1111111101111101;
    assign weights1[49][466] = 16'b1111111111110110;
    assign weights1[49][467] = 16'b1111111111101100;
    assign weights1[49][468] = 16'b1111111111100100;
    assign weights1[49][469] = 16'b1111111111101100;
    assign weights1[49][470] = 16'b1111111111101111;
    assign weights1[49][471] = 16'b1111111111100111;
    assign weights1[49][472] = 16'b0000000000000001;
    assign weights1[49][473] = 16'b1111111111110001;
    assign weights1[49][474] = 16'b1111111111110110;
    assign weights1[49][475] = 16'b0000000000001001;
    assign weights1[49][476] = 16'b1111111111110110;
    assign weights1[49][477] = 16'b1111111111110001;
    assign weights1[49][478] = 16'b1111111111110011;
    assign weights1[49][479] = 16'b1111111111110101;
    assign weights1[49][480] = 16'b1111111111101101;
    assign weights1[49][481] = 16'b1111111111100000;
    assign weights1[49][482] = 16'b1111111111111111;
    assign weights1[49][483] = 16'b1111111111110011;
    assign weights1[49][484] = 16'b1111111111110100;
    assign weights1[49][485] = 16'b1111111111111000;
    assign weights1[49][486] = 16'b0000000000010111;
    assign weights1[49][487] = 16'b0000000000011011;
    assign weights1[49][488] = 16'b0000000000101001;
    assign weights1[49][489] = 16'b1111111111101111;
    assign weights1[49][490] = 16'b1111111111110111;
    assign weights1[49][491] = 16'b1111111110111001;
    assign weights1[49][492] = 16'b1111111101000110;
    assign weights1[49][493] = 16'b1111111110101100;
    assign weights1[49][494] = 16'b1111111111100010;
    assign weights1[49][495] = 16'b1111111111110010;
    assign weights1[49][496] = 16'b1111111111100111;
    assign weights1[49][497] = 16'b1111111111101000;
    assign weights1[49][498] = 16'b1111111111110011;
    assign weights1[49][499] = 16'b1111111111110011;
    assign weights1[49][500] = 16'b1111111111111100;
    assign weights1[49][501] = 16'b1111111111110100;
    assign weights1[49][502] = 16'b1111111111111000;
    assign weights1[49][503] = 16'b0000000000000000;
    assign weights1[49][504] = 16'b1111111111110001;
    assign weights1[49][505] = 16'b1111111111111110;
    assign weights1[49][506] = 16'b1111111111111011;
    assign weights1[49][507] = 16'b1111111111111001;
    assign weights1[49][508] = 16'b0000000000000110;
    assign weights1[49][509] = 16'b1111111111111011;
    assign weights1[49][510] = 16'b0000000000000111;
    assign weights1[49][511] = 16'b1111111111111011;
    assign weights1[49][512] = 16'b1111111111111011;
    assign weights1[49][513] = 16'b1111111111111111;
    assign weights1[49][514] = 16'b0000000000011100;
    assign weights1[49][515] = 16'b0000000000000101;
    assign weights1[49][516] = 16'b0000000000000110;
    assign weights1[49][517] = 16'b1111111111110010;
    assign weights1[49][518] = 16'b1111111111110101;
    assign weights1[49][519] = 16'b1111111101111010;
    assign weights1[49][520] = 16'b1111111101100111;
    assign weights1[49][521] = 16'b1111111111100011;
    assign weights1[49][522] = 16'b1111111111111010;
    assign weights1[49][523] = 16'b1111111111100011;
    assign weights1[49][524] = 16'b1111111111111010;
    assign weights1[49][525] = 16'b1111111111110100;
    assign weights1[49][526] = 16'b1111111111111000;
    assign weights1[49][527] = 16'b1111111111111100;
    assign weights1[49][528] = 16'b1111111111111001;
    assign weights1[49][529] = 16'b1111111111110111;
    assign weights1[49][530] = 16'b1111111111110101;
    assign weights1[49][531] = 16'b0000000000000010;
    assign weights1[49][532] = 16'b1111111111111010;
    assign weights1[49][533] = 16'b1111111111111101;
    assign weights1[49][534] = 16'b0000000000001000;
    assign weights1[49][535] = 16'b0000000000001000;
    assign weights1[49][536] = 16'b0000000000000000;
    assign weights1[49][537] = 16'b0000000000010010;
    assign weights1[49][538] = 16'b0000000000001100;
    assign weights1[49][539] = 16'b1111111111110101;
    assign weights1[49][540] = 16'b1111111111110101;
    assign weights1[49][541] = 16'b0000000000001101;
    assign weights1[49][542] = 16'b1111111111111010;
    assign weights1[49][543] = 16'b1111111111111101;
    assign weights1[49][544] = 16'b1111111111111100;
    assign weights1[49][545] = 16'b1111111111100001;
    assign weights1[49][546] = 16'b1111111111000010;
    assign weights1[49][547] = 16'b1111111101000000;
    assign weights1[49][548] = 16'b1111111110101011;
    assign weights1[49][549] = 16'b1111111111100111;
    assign weights1[49][550] = 16'b1111111111110101;
    assign weights1[49][551] = 16'b1111111111110001;
    assign weights1[49][552] = 16'b1111111111111010;
    assign weights1[49][553] = 16'b1111111111111010;
    assign weights1[49][554] = 16'b0000000000000000;
    assign weights1[49][555] = 16'b1111111111110011;
    assign weights1[49][556] = 16'b1111111111101110;
    assign weights1[49][557] = 16'b0000000000000011;
    assign weights1[49][558] = 16'b1111111111111011;
    assign weights1[49][559] = 16'b1111111111111100;
    assign weights1[49][560] = 16'b1111111111111111;
    assign weights1[49][561] = 16'b0000000000000111;
    assign weights1[49][562] = 16'b0000000000010011;
    assign weights1[49][563] = 16'b0000000000001011;
    assign weights1[49][564] = 16'b0000000000000111;
    assign weights1[49][565] = 16'b0000000000000101;
    assign weights1[49][566] = 16'b0000000000000010;
    assign weights1[49][567] = 16'b1111111111111010;
    assign weights1[49][568] = 16'b1111111111111000;
    assign weights1[49][569] = 16'b1111111111110111;
    assign weights1[49][570] = 16'b1111111111111100;
    assign weights1[49][571] = 16'b0000000000001111;
    assign weights1[49][572] = 16'b1111111111101010;
    assign weights1[49][573] = 16'b1111111111100001;
    assign weights1[49][574] = 16'b1111111110101011;
    assign weights1[49][575] = 16'b1111111110100000;
    assign weights1[49][576] = 16'b1111111111110000;
    assign weights1[49][577] = 16'b0000000000000110;
    assign weights1[49][578] = 16'b0000000000000001;
    assign weights1[49][579] = 16'b0000000000001110;
    assign weights1[49][580] = 16'b0000000000000010;
    assign weights1[49][581] = 16'b1111111111110011;
    assign weights1[49][582] = 16'b0000000000000101;
    assign weights1[49][583] = 16'b1111111111111000;
    assign weights1[49][584] = 16'b1111111111110111;
    assign weights1[49][585] = 16'b1111111111111101;
    assign weights1[49][586] = 16'b1111111111111010;
    assign weights1[49][587] = 16'b0000000000000101;
    assign weights1[49][588] = 16'b0000000000000100;
    assign weights1[49][589] = 16'b0000000000000001;
    assign weights1[49][590] = 16'b0000000000010011;
    assign weights1[49][591] = 16'b0000000000010010;
    assign weights1[49][592] = 16'b0000000000010000;
    assign weights1[49][593] = 16'b1111111111100011;
    assign weights1[49][594] = 16'b1111111111110101;
    assign weights1[49][595] = 16'b1111111111110101;
    assign weights1[49][596] = 16'b0000000000011001;
    assign weights1[49][597] = 16'b1111111111111100;
    assign weights1[49][598] = 16'b1111111111111001;
    assign weights1[49][599] = 16'b1111111111101111;
    assign weights1[49][600] = 16'b1111111111111101;
    assign weights1[49][601] = 16'b1111111111011100;
    assign weights1[49][602] = 16'b1111111111101001;
    assign weights1[49][603] = 16'b1111111111101111;
    assign weights1[49][604] = 16'b0000000000000010;
    assign weights1[49][605] = 16'b0000000000000011;
    assign weights1[49][606] = 16'b1111111111111101;
    assign weights1[49][607] = 16'b0000000000000110;
    assign weights1[49][608] = 16'b0000000000001101;
    assign weights1[49][609] = 16'b0000000000001010;
    assign weights1[49][610] = 16'b0000000000000110;
    assign weights1[49][611] = 16'b1111111111110101;
    assign weights1[49][612] = 16'b0000000000000000;
    assign weights1[49][613] = 16'b1111111111111111;
    assign weights1[49][614] = 16'b0000000000000001;
    assign weights1[49][615] = 16'b0000000000001000;
    assign weights1[49][616] = 16'b0000000000000111;
    assign weights1[49][617] = 16'b0000000000000110;
    assign weights1[49][618] = 16'b0000000000010001;
    assign weights1[49][619] = 16'b0000000000000010;
    assign weights1[49][620] = 16'b0000000000000110;
    assign weights1[49][621] = 16'b1111111111110100;
    assign weights1[49][622] = 16'b0000000000000111;
    assign weights1[49][623] = 16'b1111111111110010;
    assign weights1[49][624] = 16'b0000000000001110;
    assign weights1[49][625] = 16'b1111111111111001;
    assign weights1[49][626] = 16'b1111111111111111;
    assign weights1[49][627] = 16'b1111111111110100;
    assign weights1[49][628] = 16'b0000000000000100;
    assign weights1[49][629] = 16'b0000000000001101;
    assign weights1[49][630] = 16'b0000000000010011;
    assign weights1[49][631] = 16'b1111111111110010;
    assign weights1[49][632] = 16'b0000000000000001;
    assign weights1[49][633] = 16'b1111111111111101;
    assign weights1[49][634] = 16'b1111111111111000;
    assign weights1[49][635] = 16'b0000000000001000;
    assign weights1[49][636] = 16'b0000000000010001;
    assign weights1[49][637] = 16'b1111111111111100;
    assign weights1[49][638] = 16'b1111111111111001;
    assign weights1[49][639] = 16'b0000000000000011;
    assign weights1[49][640] = 16'b0000000000000100;
    assign weights1[49][641] = 16'b0000000000001000;
    assign weights1[49][642] = 16'b0000000000001010;
    assign weights1[49][643] = 16'b0000000000001011;
    assign weights1[49][644] = 16'b0000000000000011;
    assign weights1[49][645] = 16'b0000000000001110;
    assign weights1[49][646] = 16'b0000000000000011;
    assign weights1[49][647] = 16'b0000000000000001;
    assign weights1[49][648] = 16'b0000000000010010;
    assign weights1[49][649] = 16'b0000000000010110;
    assign weights1[49][650] = 16'b0000000000000001;
    assign weights1[49][651] = 16'b0000000000010010;
    assign weights1[49][652] = 16'b1111111111111001;
    assign weights1[49][653] = 16'b0000000000000000;
    assign weights1[49][654] = 16'b1111111111100100;
    assign weights1[49][655] = 16'b0000000000000010;
    assign weights1[49][656] = 16'b1111111111110000;
    assign weights1[49][657] = 16'b0000000000011110;
    assign weights1[49][658] = 16'b0000000000011000;
    assign weights1[49][659] = 16'b0000000000011110;
    assign weights1[49][660] = 16'b1111111111111111;
    assign weights1[49][661] = 16'b0000000000001100;
    assign weights1[49][662] = 16'b0000000000001000;
    assign weights1[49][663] = 16'b1111111111111000;
    assign weights1[49][664] = 16'b0000000000010100;
    assign weights1[49][665] = 16'b0000000000001000;
    assign weights1[49][666] = 16'b0000000000000110;
    assign weights1[49][667] = 16'b0000000000010010;
    assign weights1[49][668] = 16'b0000000000000100;
    assign weights1[49][669] = 16'b0000000000010010;
    assign weights1[49][670] = 16'b0000000000001111;
    assign weights1[49][671] = 16'b0000000000000110;
    assign weights1[49][672] = 16'b0000000000000010;
    assign weights1[49][673] = 16'b0000000000000111;
    assign weights1[49][674] = 16'b0000000000000100;
    assign weights1[49][675] = 16'b1111111111111010;
    assign weights1[49][676] = 16'b0000000000001001;
    assign weights1[49][677] = 16'b0000000000000101;
    assign weights1[49][678] = 16'b1111111111111111;
    assign weights1[49][679] = 16'b0000000000011010;
    assign weights1[49][680] = 16'b0000000000001100;
    assign weights1[49][681] = 16'b1111111111111111;
    assign weights1[49][682] = 16'b0000000000000110;
    assign weights1[49][683] = 16'b1111111111111010;
    assign weights1[49][684] = 16'b0000000000001110;
    assign weights1[49][685] = 16'b0000000000011000;
    assign weights1[49][686] = 16'b0000000000101101;
    assign weights1[49][687] = 16'b0000000000011111;
    assign weights1[49][688] = 16'b0000000000100001;
    assign weights1[49][689] = 16'b0000000000100010;
    assign weights1[49][690] = 16'b0000000000001110;
    assign weights1[49][691] = 16'b0000000000001011;
    assign weights1[49][692] = 16'b0000000000000000;
    assign weights1[49][693] = 16'b1111111111111001;
    assign weights1[49][694] = 16'b0000000000001011;
    assign weights1[49][695] = 16'b0000000000001111;
    assign weights1[49][696] = 16'b0000000000001110;
    assign weights1[49][697] = 16'b0000000000001110;
    assign weights1[49][698] = 16'b0000000000000011;
    assign weights1[49][699] = 16'b0000000000000000;
    assign weights1[49][700] = 16'b0000000000000110;
    assign weights1[49][701] = 16'b0000000000001011;
    assign weights1[49][702] = 16'b0000000000000111;
    assign weights1[49][703] = 16'b0000000000000100;
    assign weights1[49][704] = 16'b0000000000010101;
    assign weights1[49][705] = 16'b1111111111111110;
    assign weights1[49][706] = 16'b0000000000000100;
    assign weights1[49][707] = 16'b0000000000001011;
    assign weights1[49][708] = 16'b1111111111111100;
    assign weights1[49][709] = 16'b1111111111110111;
    assign weights1[49][710] = 16'b0000000000100010;
    assign weights1[49][711] = 16'b0000000000010111;
    assign weights1[49][712] = 16'b0000000000011101;
    assign weights1[49][713] = 16'b0000000000101101;
    assign weights1[49][714] = 16'b0000000000100010;
    assign weights1[49][715] = 16'b0000000000101101;
    assign weights1[49][716] = 16'b0000000000110000;
    assign weights1[49][717] = 16'b0000000000101100;
    assign weights1[49][718] = 16'b0000000000100101;
    assign weights1[49][719] = 16'b0000000000010100;
    assign weights1[49][720] = 16'b0000000000011000;
    assign weights1[49][721] = 16'b0000000000000101;
    assign weights1[49][722] = 16'b0000000000010100;
    assign weights1[49][723] = 16'b0000000000000001;
    assign weights1[49][724] = 16'b0000000000001110;
    assign weights1[49][725] = 16'b0000000000000110;
    assign weights1[49][726] = 16'b0000000000000001;
    assign weights1[49][727] = 16'b1111111111111110;
    assign weights1[49][728] = 16'b0000000000000101;
    assign weights1[49][729] = 16'b0000000000001011;
    assign weights1[49][730] = 16'b0000000000001011;
    assign weights1[49][731] = 16'b0000000000001000;
    assign weights1[49][732] = 16'b0000000000001100;
    assign weights1[49][733] = 16'b0000000000000110;
    assign weights1[49][734] = 16'b0000000000000111;
    assign weights1[49][735] = 16'b0000000000001011;
    assign weights1[49][736] = 16'b1111111111111110;
    assign weights1[49][737] = 16'b1111111111111000;
    assign weights1[49][738] = 16'b1111111111111110;
    assign weights1[49][739] = 16'b0000000000010001;
    assign weights1[49][740] = 16'b0000000000010001;
    assign weights1[49][741] = 16'b0000000000011000;
    assign weights1[49][742] = 16'b0000000000010010;
    assign weights1[49][743] = 16'b0000000000010111;
    assign weights1[49][744] = 16'b0000000000101000;
    assign weights1[49][745] = 16'b0000000000011010;
    assign weights1[49][746] = 16'b0000000000011100;
    assign weights1[49][747] = 16'b0000000000001110;
    assign weights1[49][748] = 16'b0000000000010110;
    assign weights1[49][749] = 16'b0000000000000101;
    assign weights1[49][750] = 16'b0000000000010110;
    assign weights1[49][751] = 16'b0000000000000001;
    assign weights1[49][752] = 16'b0000000000000010;
    assign weights1[49][753] = 16'b1111111111111001;
    assign weights1[49][754] = 16'b1111111111111101;
    assign weights1[49][755] = 16'b1111111111111101;
    assign weights1[49][756] = 16'b0000000000000000;
    assign weights1[49][757] = 16'b0000000000000110;
    assign weights1[49][758] = 16'b0000000000001000;
    assign weights1[49][759] = 16'b0000000000001011;
    assign weights1[49][760] = 16'b0000000000000101;
    assign weights1[49][761] = 16'b0000000000000101;
    assign weights1[49][762] = 16'b1111111111111111;
    assign weights1[49][763] = 16'b1111111111111001;
    assign weights1[49][764] = 16'b0000000000000000;
    assign weights1[49][765] = 16'b1111111111111101;
    assign weights1[49][766] = 16'b0000000000000010;
    assign weights1[49][767] = 16'b0000000000010101;
    assign weights1[49][768] = 16'b0000000000100001;
    assign weights1[49][769] = 16'b0000000000011101;
    assign weights1[49][770] = 16'b0000000000100000;
    assign weights1[49][771] = 16'b0000000000010000;
    assign weights1[49][772] = 16'b0000000000010110;
    assign weights1[49][773] = 16'b0000000000011111;
    assign weights1[49][774] = 16'b0000000000001111;
    assign weights1[49][775] = 16'b0000000000001110;
    assign weights1[49][776] = 16'b0000000000011001;
    assign weights1[49][777] = 16'b0000000000001010;
    assign weights1[49][778] = 16'b0000000000001001;
    assign weights1[49][779] = 16'b1111111111110010;
    assign weights1[49][780] = 16'b1111111111111000;
    assign weights1[49][781] = 16'b1111111111110101;
    assign weights1[49][782] = 16'b1111111111111010;
    assign weights1[49][783] = 16'b1111111111111110;
    assign weights1[50][0] = 16'b0000000000000001;
    assign weights1[50][1] = 16'b0000000000000001;
    assign weights1[50][2] = 16'b0000000000000001;
    assign weights1[50][3] = 16'b1111111111111111;
    assign weights1[50][4] = 16'b1111111111111010;
    assign weights1[50][5] = 16'b1111111111101010;
    assign weights1[50][6] = 16'b1111111111100100;
    assign weights1[50][7] = 16'b1111111111101011;
    assign weights1[50][8] = 16'b1111111111100010;
    assign weights1[50][9] = 16'b1111111111011110;
    assign weights1[50][10] = 16'b1111111111011010;
    assign weights1[50][11] = 16'b1111111111101110;
    assign weights1[50][12] = 16'b1111111111110001;
    assign weights1[50][13] = 16'b1111111111100111;
    assign weights1[50][14] = 16'b0000000000000001;
    assign weights1[50][15] = 16'b1111111111111110;
    assign weights1[50][16] = 16'b0000000000000001;
    assign weights1[50][17] = 16'b0000000000010000;
    assign weights1[50][18] = 16'b0000000000010101;
    assign weights1[50][19] = 16'b0000000000100100;
    assign weights1[50][20] = 16'b0000000000100100;
    assign weights1[50][21] = 16'b0000000000100101;
    assign weights1[50][22] = 16'b0000000000001110;
    assign weights1[50][23] = 16'b0000000000100000;
    assign weights1[50][24] = 16'b0000000000011000;
    assign weights1[50][25] = 16'b0000000000011001;
    assign weights1[50][26] = 16'b0000000000001101;
    assign weights1[50][27] = 16'b0000000000000100;
    assign weights1[50][28] = 16'b0000000000000001;
    assign weights1[50][29] = 16'b0000000000000001;
    assign weights1[50][30] = 16'b0000000000000001;
    assign weights1[50][31] = 16'b1111111111111110;
    assign weights1[50][32] = 16'b1111111111110010;
    assign weights1[50][33] = 16'b1111111111101011;
    assign weights1[50][34] = 16'b1111111111100110;
    assign weights1[50][35] = 16'b1111111111101010;
    assign weights1[50][36] = 16'b1111111111100000;
    assign weights1[50][37] = 16'b1111111111011100;
    assign weights1[50][38] = 16'b1111111111100110;
    assign weights1[50][39] = 16'b1111111111111001;
    assign weights1[50][40] = 16'b1111111111111100;
    assign weights1[50][41] = 16'b1111111111110001;
    assign weights1[50][42] = 16'b0000000000000110;
    assign weights1[50][43] = 16'b1111111111111101;
    assign weights1[50][44] = 16'b1111111111111111;
    assign weights1[50][45] = 16'b0000000000001111;
    assign weights1[50][46] = 16'b0000000000011011;
    assign weights1[50][47] = 16'b0000000000011101;
    assign weights1[50][48] = 16'b0000000000011001;
    assign weights1[50][49] = 16'b0000000000100111;
    assign weights1[50][50] = 16'b0000000000100101;
    assign weights1[50][51] = 16'b0000000000100010;
    assign weights1[50][52] = 16'b0000000000101111;
    assign weights1[50][53] = 16'b0000000000100101;
    assign weights1[50][54] = 16'b0000000000011110;
    assign weights1[50][55] = 16'b0000000000001001;
    assign weights1[50][56] = 16'b1111111111111111;
    assign weights1[50][57] = 16'b0000000000000000;
    assign weights1[50][58] = 16'b1111111111111110;
    assign weights1[50][59] = 16'b1111111111111010;
    assign weights1[50][60] = 16'b1111111111101000;
    assign weights1[50][61] = 16'b1111111111110100;
    assign weights1[50][62] = 16'b1111111111110010;
    assign weights1[50][63] = 16'b1111111111110110;
    assign weights1[50][64] = 16'b1111111111100010;
    assign weights1[50][65] = 16'b0000000000001101;
    assign weights1[50][66] = 16'b0000000000001101;
    assign weights1[50][67] = 16'b0000000000001010;
    assign weights1[50][68] = 16'b0000000000000000;
    assign weights1[50][69] = 16'b0000000000001101;
    assign weights1[50][70] = 16'b0000000000010000;
    assign weights1[50][71] = 16'b0000000000011100;
    assign weights1[50][72] = 16'b0000000000010000;
    assign weights1[50][73] = 16'b0000000000011001;
    assign weights1[50][74] = 16'b0000000000011101;
    assign weights1[50][75] = 16'b0000000000011001;
    assign weights1[50][76] = 16'b0000000000011000;
    assign weights1[50][77] = 16'b0000000000100100;
    assign weights1[50][78] = 16'b0000000000101111;
    assign weights1[50][79] = 16'b0000000000010111;
    assign weights1[50][80] = 16'b0000000000100110;
    assign weights1[50][81] = 16'b0000000000100001;
    assign weights1[50][82] = 16'b0000000000011101;
    assign weights1[50][83] = 16'b0000000000010101;
    assign weights1[50][84] = 16'b1111111111111101;
    assign weights1[50][85] = 16'b1111111111111010;
    assign weights1[50][86] = 16'b1111111111110111;
    assign weights1[50][87] = 16'b1111111111101110;
    assign weights1[50][88] = 16'b1111111111101010;
    assign weights1[50][89] = 16'b1111111111110000;
    assign weights1[50][90] = 16'b1111111111101110;
    assign weights1[50][91] = 16'b1111111111110110;
    assign weights1[50][92] = 16'b1111111111111010;
    assign weights1[50][93] = 16'b0000000000000010;
    assign weights1[50][94] = 16'b0000000000010010;
    assign weights1[50][95] = 16'b0000000000000101;
    assign weights1[50][96] = 16'b0000000000001110;
    assign weights1[50][97] = 16'b0000000000011100;
    assign weights1[50][98] = 16'b1111111111110111;
    assign weights1[50][99] = 16'b0000000000011110;
    assign weights1[50][100] = 16'b0000000000011101;
    assign weights1[50][101] = 16'b0000000000001010;
    assign weights1[50][102] = 16'b0000000000011011;
    assign weights1[50][103] = 16'b0000000000010101;
    assign weights1[50][104] = 16'b0000000000100101;
    assign weights1[50][105] = 16'b0000000000011100;
    assign weights1[50][106] = 16'b0000000000100111;
    assign weights1[50][107] = 16'b0000000000100110;
    assign weights1[50][108] = 16'b0000000000101110;
    assign weights1[50][109] = 16'b0000000000011010;
    assign weights1[50][110] = 16'b0000000000011010;
    assign weights1[50][111] = 16'b0000000000001011;
    assign weights1[50][112] = 16'b1111111111111011;
    assign weights1[50][113] = 16'b1111111111110001;
    assign weights1[50][114] = 16'b1111111111110101;
    assign weights1[50][115] = 16'b1111111111110011;
    assign weights1[50][116] = 16'b1111111111100000;
    assign weights1[50][117] = 16'b0000000000000101;
    assign weights1[50][118] = 16'b0000000000000010;
    assign weights1[50][119] = 16'b0000000000001000;
    assign weights1[50][120] = 16'b1111111111110100;
    assign weights1[50][121] = 16'b0000000000000110;
    assign weights1[50][122] = 16'b0000000000100000;
    assign weights1[50][123] = 16'b0000000000010010;
    assign weights1[50][124] = 16'b0000000000001000;
    assign weights1[50][125] = 16'b0000000000001101;
    assign weights1[50][126] = 16'b0000000000100001;
    assign weights1[50][127] = 16'b0000000000101001;
    assign weights1[50][128] = 16'b0000000000001111;
    assign weights1[50][129] = 16'b0000000000010001;
    assign weights1[50][130] = 16'b0000000000010110;
    assign weights1[50][131] = 16'b0000000000010001;
    assign weights1[50][132] = 16'b0000000000110001;
    assign weights1[50][133] = 16'b0000000001000101;
    assign weights1[50][134] = 16'b0000000001001010;
    assign weights1[50][135] = 16'b0000000000111010;
    assign weights1[50][136] = 16'b0000000000110111;
    assign weights1[50][137] = 16'b0000000000010010;
    assign weights1[50][138] = 16'b1111111111111011;
    assign weights1[50][139] = 16'b1111111111110100;
    assign weights1[50][140] = 16'b1111111111111101;
    assign weights1[50][141] = 16'b1111111111101101;
    assign weights1[50][142] = 16'b1111111111101001;
    assign weights1[50][143] = 16'b1111111111101001;
    assign weights1[50][144] = 16'b1111111111110100;
    assign weights1[50][145] = 16'b1111111111111011;
    assign weights1[50][146] = 16'b1111111111111111;
    assign weights1[50][147] = 16'b1111111111111001;
    assign weights1[50][148] = 16'b0000000000000001;
    assign weights1[50][149] = 16'b0000000000000011;
    assign weights1[50][150] = 16'b0000000000000001;
    assign weights1[50][151] = 16'b0000000000001110;
    assign weights1[50][152] = 16'b0000000000001001;
    assign weights1[50][153] = 16'b0000000000011100;
    assign weights1[50][154] = 16'b0000000000001000;
    assign weights1[50][155] = 16'b0000000000010101;
    assign weights1[50][156] = 16'b0000000000010000;
    assign weights1[50][157] = 16'b0000000000111100;
    assign weights1[50][158] = 16'b0000000000101101;
    assign weights1[50][159] = 16'b0000000000110011;
    assign weights1[50][160] = 16'b0000000001011010;
    assign weights1[50][161] = 16'b0000000000111100;
    assign weights1[50][162] = 16'b0000000000101001;
    assign weights1[50][163] = 16'b0000000000010110;
    assign weights1[50][164] = 16'b0000000000001110;
    assign weights1[50][165] = 16'b1111111111100110;
    assign weights1[50][166] = 16'b1111111111010000;
    assign weights1[50][167] = 16'b1111111111011111;
    assign weights1[50][168] = 16'b1111111111111011;
    assign weights1[50][169] = 16'b1111111111110001;
    assign weights1[50][170] = 16'b0000000000000001;
    assign weights1[50][171] = 16'b1111111111101111;
    assign weights1[50][172] = 16'b1111111111111000;
    assign weights1[50][173] = 16'b1111111111111001;
    assign weights1[50][174] = 16'b0000000000000010;
    assign weights1[50][175] = 16'b1111111111111011;
    assign weights1[50][176] = 16'b0000000000001110;
    assign weights1[50][177] = 16'b0000000000011000;
    assign weights1[50][178] = 16'b0000000000001011;
    assign weights1[50][179] = 16'b0000000000001111;
    assign weights1[50][180] = 16'b0000000000010000;
    assign weights1[50][181] = 16'b0000000000000010;
    assign weights1[50][182] = 16'b0000000000011111;
    assign weights1[50][183] = 16'b0000000000100000;
    assign weights1[50][184] = 16'b0000000000111011;
    assign weights1[50][185] = 16'b0000000000100100;
    assign weights1[50][186] = 16'b0000000000110110;
    assign weights1[50][187] = 16'b0000000000111000;
    assign weights1[50][188] = 16'b1111111111110110;
    assign weights1[50][189] = 16'b1111111111100001;
    assign weights1[50][190] = 16'b1111111111001010;
    assign weights1[50][191] = 16'b1111111110011001;
    assign weights1[50][192] = 16'b1111111110100001;
    assign weights1[50][193] = 16'b1111111110011101;
    assign weights1[50][194] = 16'b1111111110101110;
    assign weights1[50][195] = 16'b1111111111000000;
    assign weights1[50][196] = 16'b1111111111111001;
    assign weights1[50][197] = 16'b1111111111110101;
    assign weights1[50][198] = 16'b1111111111110100;
    assign weights1[50][199] = 16'b1111111111111000;
    assign weights1[50][200] = 16'b0000000000000010;
    assign weights1[50][201] = 16'b0000000000000110;
    assign weights1[50][202] = 16'b0000000000001111;
    assign weights1[50][203] = 16'b0000000000000010;
    assign weights1[50][204] = 16'b0000000000000001;
    assign weights1[50][205] = 16'b0000000000000010;
    assign weights1[50][206] = 16'b0000000000010001;
    assign weights1[50][207] = 16'b0000000000001010;
    assign weights1[50][208] = 16'b0000000000010101;
    assign weights1[50][209] = 16'b1111111111110111;
    assign weights1[50][210] = 16'b0000000000000010;
    assign weights1[50][211] = 16'b1111111111111001;
    assign weights1[50][212] = 16'b1111111111100110;
    assign weights1[50][213] = 16'b1111111110111110;
    assign weights1[50][214] = 16'b1111111110001001;
    assign weights1[50][215] = 16'b1111111101011010;
    assign weights1[50][216] = 16'b1111111101001111;
    assign weights1[50][217] = 16'b1111111101001011;
    assign weights1[50][218] = 16'b1111111101000010;
    assign weights1[50][219] = 16'b1111111101100011;
    assign weights1[50][220] = 16'b1111111101111010;
    assign weights1[50][221] = 16'b1111111110001000;
    assign weights1[50][222] = 16'b1111111110010111;
    assign weights1[50][223] = 16'b1111111110011110;
    assign weights1[50][224] = 16'b1111111111110100;
    assign weights1[50][225] = 16'b1111111111110010;
    assign weights1[50][226] = 16'b1111111111111010;
    assign weights1[50][227] = 16'b1111111111111100;
    assign weights1[50][228] = 16'b1111111111111100;
    assign weights1[50][229] = 16'b0000000000000001;
    assign weights1[50][230] = 16'b0000000000000100;
    assign weights1[50][231] = 16'b1111111111111100;
    assign weights1[50][232] = 16'b0000000000001101;
    assign weights1[50][233] = 16'b0000000000000001;
    assign weights1[50][234] = 16'b0000000000000100;
    assign weights1[50][235] = 16'b1111111111101110;
    assign weights1[50][236] = 16'b1111111111101110;
    assign weights1[50][237] = 16'b1111111111001100;
    assign weights1[50][238] = 16'b1111111110010111;
    assign weights1[50][239] = 16'b1111111101100111;
    assign weights1[50][240] = 16'b1111111100110011;
    assign weights1[50][241] = 16'b1111111011110010;
    assign weights1[50][242] = 16'b1111111011101110;
    assign weights1[50][243] = 16'b1111111011111101;
    assign weights1[50][244] = 16'b1111111100101011;
    assign weights1[50][245] = 16'b1111111100110011;
    assign weights1[50][246] = 16'b1111111101010101;
    assign weights1[50][247] = 16'b1111111101100011;
    assign weights1[50][248] = 16'b1111111101101100;
    assign weights1[50][249] = 16'b1111111110000000;
    assign weights1[50][250] = 16'b1111111110000010;
    assign weights1[50][251] = 16'b1111111110001101;
    assign weights1[50][252] = 16'b1111111111101111;
    assign weights1[50][253] = 16'b0000000000000100;
    assign weights1[50][254] = 16'b0000000000001100;
    assign weights1[50][255] = 16'b1111111111111111;
    assign weights1[50][256] = 16'b0000000000001111;
    assign weights1[50][257] = 16'b0000000000001000;
    assign weights1[50][258] = 16'b0000000000001010;
    assign weights1[50][259] = 16'b1111111111111110;
    assign weights1[50][260] = 16'b0000000000000011;
    assign weights1[50][261] = 16'b1111111111111011;
    assign weights1[50][262] = 16'b1111111111111010;
    assign weights1[50][263] = 16'b1111111111110001;
    assign weights1[50][264] = 16'b1111111111110001;
    assign weights1[50][265] = 16'b1111111111010110;
    assign weights1[50][266] = 16'b1111111111011111;
    assign weights1[50][267] = 16'b1111111111101000;
    assign weights1[50][268] = 16'b1111111111100100;
    assign weights1[50][269] = 16'b1111111111011011;
    assign weights1[50][270] = 16'b1111111111000010;
    assign weights1[50][271] = 16'b1111111110101001;
    assign weights1[50][272] = 16'b1111111110000010;
    assign weights1[50][273] = 16'b1111111101010101;
    assign weights1[50][274] = 16'b1111111101011100;
    assign weights1[50][275] = 16'b1111111101100011;
    assign weights1[50][276] = 16'b1111111101110100;
    assign weights1[50][277] = 16'b1111111110000001;
    assign weights1[50][278] = 16'b1111111110100101;
    assign weights1[50][279] = 16'b1111111110100110;
    assign weights1[50][280] = 16'b1111111111110000;
    assign weights1[50][281] = 16'b1111111111111110;
    assign weights1[50][282] = 16'b0000000000000011;
    assign weights1[50][283] = 16'b0000000000001101;
    assign weights1[50][284] = 16'b1111111111111101;
    assign weights1[50][285] = 16'b0000000000000001;
    assign weights1[50][286] = 16'b1111111111111100;
    assign weights1[50][287] = 16'b0000000000000000;
    assign weights1[50][288] = 16'b0000000000000001;
    assign weights1[50][289] = 16'b0000000000000001;
    assign weights1[50][290] = 16'b1111111111111011;
    assign weights1[50][291] = 16'b1111111111110001;
    assign weights1[50][292] = 16'b1111111111111110;
    assign weights1[50][293] = 16'b1111111111110011;
    assign weights1[50][294] = 16'b0000000000000010;
    assign weights1[50][295] = 16'b0000000000000000;
    assign weights1[50][296] = 16'b1111111111111001;
    assign weights1[50][297] = 16'b0000000000001000;
    assign weights1[50][298] = 16'b1111111111110010;
    assign weights1[50][299] = 16'b1111111111111100;
    assign weights1[50][300] = 16'b1111111111100111;
    assign weights1[50][301] = 16'b1111111111101111;
    assign weights1[50][302] = 16'b1111111111011101;
    assign weights1[50][303] = 16'b1111111111011100;
    assign weights1[50][304] = 16'b1111111111001011;
    assign weights1[50][305] = 16'b1111111111101011;
    assign weights1[50][306] = 16'b1111111111010100;
    assign weights1[50][307] = 16'b1111111111001001;
    assign weights1[50][308] = 16'b1111111111110101;
    assign weights1[50][309] = 16'b1111111111111100;
    assign weights1[50][310] = 16'b0000000000001000;
    assign weights1[50][311] = 16'b0000000000001001;
    assign weights1[50][312] = 16'b0000000000000011;
    assign weights1[50][313] = 16'b0000000000001001;
    assign weights1[50][314] = 16'b0000000000000000;
    assign weights1[50][315] = 16'b0000000000000011;
    assign weights1[50][316] = 16'b1111111111111010;
    assign weights1[50][317] = 16'b0000000000000110;
    assign weights1[50][318] = 16'b1111111111111000;
    assign weights1[50][319] = 16'b0000000000000101;
    assign weights1[50][320] = 16'b0000000000000000;
    assign weights1[50][321] = 16'b0000000000000001;
    assign weights1[50][322] = 16'b1111111111111010;
    assign weights1[50][323] = 16'b1111111111110001;
    assign weights1[50][324] = 16'b0000000000010001;
    assign weights1[50][325] = 16'b0000000000001010;
    assign weights1[50][326] = 16'b0000000000010001;
    assign weights1[50][327] = 16'b0000000000011001;
    assign weights1[50][328] = 16'b0000000000100011;
    assign weights1[50][329] = 16'b0000000000000110;
    assign weights1[50][330] = 16'b0000000000010100;
    assign weights1[50][331] = 16'b0000000000001111;
    assign weights1[50][332] = 16'b0000000000100010;
    assign weights1[50][333] = 16'b0000000000010001;
    assign weights1[50][334] = 16'b0000000000001001;
    assign weights1[50][335] = 16'b0000000000000111;
    assign weights1[50][336] = 16'b1111111111111010;
    assign weights1[50][337] = 16'b0000000000000011;
    assign weights1[50][338] = 16'b1111111111111100;
    assign weights1[50][339] = 16'b0000000000001000;
    assign weights1[50][340] = 16'b0000000000001000;
    assign weights1[50][341] = 16'b0000000000001010;
    assign weights1[50][342] = 16'b0000000000010001;
    assign weights1[50][343] = 16'b0000000000000100;
    assign weights1[50][344] = 16'b1111111111110111;
    assign weights1[50][345] = 16'b1111111111110110;
    assign weights1[50][346] = 16'b1111111111111010;
    assign weights1[50][347] = 16'b0000000000001110;
    assign weights1[50][348] = 16'b1111111111101001;
    assign weights1[50][349] = 16'b1111111111111110;
    assign weights1[50][350] = 16'b1111111111111000;
    assign weights1[50][351] = 16'b1111111111101101;
    assign weights1[50][352] = 16'b0000000000000000;
    assign weights1[50][353] = 16'b1111111111110110;
    assign weights1[50][354] = 16'b0000000000010010;
    assign weights1[50][355] = 16'b0000000000010010;
    assign weights1[50][356] = 16'b0000000000011011;
    assign weights1[50][357] = 16'b0000000000110000;
    assign weights1[50][358] = 16'b0000000000010111;
    assign weights1[50][359] = 16'b0000000000010100;
    assign weights1[50][360] = 16'b0000000000100001;
    assign weights1[50][361] = 16'b0000000000001101;
    assign weights1[50][362] = 16'b0000000000110101;
    assign weights1[50][363] = 16'b0000000000110110;
    assign weights1[50][364] = 16'b1111111111111111;
    assign weights1[50][365] = 16'b1111111111111100;
    assign weights1[50][366] = 16'b0000000000000111;
    assign weights1[50][367] = 16'b1111111111111100;
    assign weights1[50][368] = 16'b0000000000000011;
    assign weights1[50][369] = 16'b1111111111111010;
    assign weights1[50][370] = 16'b1111111111111111;
    assign weights1[50][371] = 16'b0000000000000010;
    assign weights1[50][372] = 16'b0000000000000100;
    assign weights1[50][373] = 16'b1111111111111110;
    assign weights1[50][374] = 16'b0000000000000101;
    assign weights1[50][375] = 16'b1111111111111101;
    assign weights1[50][376] = 16'b1111111111110111;
    assign weights1[50][377] = 16'b0000000000000011;
    assign weights1[50][378] = 16'b0000000000000000;
    assign weights1[50][379] = 16'b0000000000001010;
    assign weights1[50][380] = 16'b0000000000001001;
    assign weights1[50][381] = 16'b0000000000010110;
    assign weights1[50][382] = 16'b0000000000001101;
    assign weights1[50][383] = 16'b0000000000011100;
    assign weights1[50][384] = 16'b0000000000010111;
    assign weights1[50][385] = 16'b0000000000010001;
    assign weights1[50][386] = 16'b0000000000010111;
    assign weights1[50][387] = 16'b0000000000010101;
    assign weights1[50][388] = 16'b0000000000101110;
    assign weights1[50][389] = 16'b0000000000001000;
    assign weights1[50][390] = 16'b0000000000001100;
    assign weights1[50][391] = 16'b0000000000110010;
    assign weights1[50][392] = 16'b1111111111110111;
    assign weights1[50][393] = 16'b0000000000000100;
    assign weights1[50][394] = 16'b0000000000000111;
    assign weights1[50][395] = 16'b0000000000001000;
    assign weights1[50][396] = 16'b1111111111111110;
    assign weights1[50][397] = 16'b0000000000010011;
    assign weights1[50][398] = 16'b1111111111110000;
    assign weights1[50][399] = 16'b0000000000001101;
    assign weights1[50][400] = 16'b1111111111110011;
    assign weights1[50][401] = 16'b1111111111111101;
    assign weights1[50][402] = 16'b1111111111111111;
    assign weights1[50][403] = 16'b1111111111111100;
    assign weights1[50][404] = 16'b1111111111111011;
    assign weights1[50][405] = 16'b1111111111111011;
    assign weights1[50][406] = 16'b0000000000000110;
    assign weights1[50][407] = 16'b0000000000000010;
    assign weights1[50][408] = 16'b1111111111110111;
    assign weights1[50][409] = 16'b0000000000001000;
    assign weights1[50][410] = 16'b0000000000010011;
    assign weights1[50][411] = 16'b0000000000000001;
    assign weights1[50][412] = 16'b0000000000001111;
    assign weights1[50][413] = 16'b0000000000000000;
    assign weights1[50][414] = 16'b0000000000000010;
    assign weights1[50][415] = 16'b1111111111110101;
    assign weights1[50][416] = 16'b0000000000001111;
    assign weights1[50][417] = 16'b0000000000000010;
    assign weights1[50][418] = 16'b0000000000101001;
    assign weights1[50][419] = 16'b0000000000100001;
    assign weights1[50][420] = 16'b0000000000000000;
    assign weights1[50][421] = 16'b1111111111111010;
    assign weights1[50][422] = 16'b0000000000001011;
    assign weights1[50][423] = 16'b1111111111110111;
    assign weights1[50][424] = 16'b0000000000000100;
    assign weights1[50][425] = 16'b0000000000010001;
    assign weights1[50][426] = 16'b0000000000000110;
    assign weights1[50][427] = 16'b0000000000001010;
    assign weights1[50][428] = 16'b0000000000000010;
    assign weights1[50][429] = 16'b1111111111111110;
    assign weights1[50][430] = 16'b1111111111111001;
    assign weights1[50][431] = 16'b1111111111100111;
    assign weights1[50][432] = 16'b1111111111110000;
    assign weights1[50][433] = 16'b1111111111110111;
    assign weights1[50][434] = 16'b1111111111111111;
    assign weights1[50][435] = 16'b0000000000000000;
    assign weights1[50][436] = 16'b0000000000000101;
    assign weights1[50][437] = 16'b1111111111111001;
    assign weights1[50][438] = 16'b0000000000000001;
    assign weights1[50][439] = 16'b1111111111110001;
    assign weights1[50][440] = 16'b1111111111110111;
    assign weights1[50][441] = 16'b1111111111110111;
    assign weights1[50][442] = 16'b0000000000000101;
    assign weights1[50][443] = 16'b1111111111011010;
    assign weights1[50][444] = 16'b1111111111111001;
    assign weights1[50][445] = 16'b0000000000000011;
    assign weights1[50][446] = 16'b0000000000001110;
    assign weights1[50][447] = 16'b0000000000001100;
    assign weights1[50][448] = 16'b1111111111110001;
    assign weights1[50][449] = 16'b1111111111111101;
    assign weights1[50][450] = 16'b0000000000001010;
    assign weights1[50][451] = 16'b0000000000001001;
    assign weights1[50][452] = 16'b1111111111111110;
    assign weights1[50][453] = 16'b1111111111110101;
    assign weights1[50][454] = 16'b0000000000000100;
    assign weights1[50][455] = 16'b1111111111111110;
    assign weights1[50][456] = 16'b0000000000000011;
    assign weights1[50][457] = 16'b1111111111111110;
    assign weights1[50][458] = 16'b1111111111111110;
    assign weights1[50][459] = 16'b1111111111111011;
    assign weights1[50][460] = 16'b0000000000001011;
    assign weights1[50][461] = 16'b1111111111111101;
    assign weights1[50][462] = 16'b1111111111111100;
    assign weights1[50][463] = 16'b1111111111111001;
    assign weights1[50][464] = 16'b1111111111110000;
    assign weights1[50][465] = 16'b0000000000001110;
    assign weights1[50][466] = 16'b1111111111111101;
    assign weights1[50][467] = 16'b1111111111111001;
    assign weights1[50][468] = 16'b1111111111110001;
    assign weights1[50][469] = 16'b1111111111111010;
    assign weights1[50][470] = 16'b0000000000000000;
    assign weights1[50][471] = 16'b1111111111100101;
    assign weights1[50][472] = 16'b1111111111101111;
    assign weights1[50][473] = 16'b1111111111110001;
    assign weights1[50][474] = 16'b1111111111101001;
    assign weights1[50][475] = 16'b0000000000011010;
    assign weights1[50][476] = 16'b1111111111111010;
    assign weights1[50][477] = 16'b0000000000000001;
    assign weights1[50][478] = 16'b1111111111110111;
    assign weights1[50][479] = 16'b1111111111110101;
    assign weights1[50][480] = 16'b1111111111101111;
    assign weights1[50][481] = 16'b1111111111111101;
    assign weights1[50][482] = 16'b0000000000001010;
    assign weights1[50][483] = 16'b0000000000000101;
    assign weights1[50][484] = 16'b0000000000000001;
    assign weights1[50][485] = 16'b0000000000001010;
    assign weights1[50][486] = 16'b0000000000000001;
    assign weights1[50][487] = 16'b0000000000000010;
    assign weights1[50][488] = 16'b1111111111110110;
    assign weights1[50][489] = 16'b1111111111111000;
    assign weights1[50][490] = 16'b0000000000000110;
    assign weights1[50][491] = 16'b1111111111110101;
    assign weights1[50][492] = 16'b1111111111101110;
    assign weights1[50][493] = 16'b1111111111110011;
    assign weights1[50][494] = 16'b1111111111101111;
    assign weights1[50][495] = 16'b0000000000001100;
    assign weights1[50][496] = 16'b0000000000000010;
    assign weights1[50][497] = 16'b0000000000010001;
    assign weights1[50][498] = 16'b1111111111110011;
    assign weights1[50][499] = 16'b0000000000000010;
    assign weights1[50][500] = 16'b0000000000000101;
    assign weights1[50][501] = 16'b1111111111100111;
    assign weights1[50][502] = 16'b0000000000000001;
    assign weights1[50][503] = 16'b0000000000001000;
    assign weights1[50][504] = 16'b0000000000001000;
    assign weights1[50][505] = 16'b0000000000001010;
    assign weights1[50][506] = 16'b0000000000000110;
    assign weights1[50][507] = 16'b0000000000000011;
    assign weights1[50][508] = 16'b0000000000001011;
    assign weights1[50][509] = 16'b0000000000001010;
    assign weights1[50][510] = 16'b1111111111111010;
    assign weights1[50][511] = 16'b1111111111110110;
    assign weights1[50][512] = 16'b0000000000000100;
    assign weights1[50][513] = 16'b1111111111110110;
    assign weights1[50][514] = 16'b1111111111111010;
    assign weights1[50][515] = 16'b1111111111111111;
    assign weights1[50][516] = 16'b1111111111111000;
    assign weights1[50][517] = 16'b1111111111111100;
    assign weights1[50][518] = 16'b1111111111111000;
    assign weights1[50][519] = 16'b1111111111111100;
    assign weights1[50][520] = 16'b1111111111110111;
    assign weights1[50][521] = 16'b1111111111110100;
    assign weights1[50][522] = 16'b0000000000001101;
    assign weights1[50][523] = 16'b0000000000000011;
    assign weights1[50][524] = 16'b1111111111111010;
    assign weights1[50][525] = 16'b0000000000000101;
    assign weights1[50][526] = 16'b1111111111111100;
    assign weights1[50][527] = 16'b1111111111111111;
    assign weights1[50][528] = 16'b1111111111111101;
    assign weights1[50][529] = 16'b1111111111111001;
    assign weights1[50][530] = 16'b1111111111111111;
    assign weights1[50][531] = 16'b1111111111111111;
    assign weights1[50][532] = 16'b1111111111110110;
    assign weights1[50][533] = 16'b0000000000001101;
    assign weights1[50][534] = 16'b1111111111111100;
    assign weights1[50][535] = 16'b1111111111111111;
    assign weights1[50][536] = 16'b1111111111110011;
    assign weights1[50][537] = 16'b1111111111111101;
    assign weights1[50][538] = 16'b1111111111111110;
    assign weights1[50][539] = 16'b0000000000000010;
    assign weights1[50][540] = 16'b1111111111111000;
    assign weights1[50][541] = 16'b1111111111111111;
    assign weights1[50][542] = 16'b0000000000000000;
    assign weights1[50][543] = 16'b0000000000000101;
    assign weights1[50][544] = 16'b0000000000001101;
    assign weights1[50][545] = 16'b0000000000000010;
    assign weights1[50][546] = 16'b0000000000000100;
    assign weights1[50][547] = 16'b0000000000000011;
    assign weights1[50][548] = 16'b1111111111111001;
    assign weights1[50][549] = 16'b0000000000000111;
    assign weights1[50][550] = 16'b1111111111101111;
    assign weights1[50][551] = 16'b1111111111110100;
    assign weights1[50][552] = 16'b0000000000000011;
    assign weights1[50][553] = 16'b1111111111101011;
    assign weights1[50][554] = 16'b0000000000000000;
    assign weights1[50][555] = 16'b1111111111110010;
    assign weights1[50][556] = 16'b0000000000001111;
    assign weights1[50][557] = 16'b1111111111111100;
    assign weights1[50][558] = 16'b1111111111111110;
    assign weights1[50][559] = 16'b0000000000000101;
    assign weights1[50][560] = 16'b1111111111110101;
    assign weights1[50][561] = 16'b1111111111101100;
    assign weights1[50][562] = 16'b0000000000000100;
    assign weights1[50][563] = 16'b0000000000000011;
    assign weights1[50][564] = 16'b1111111111110101;
    assign weights1[50][565] = 16'b1111111111111110;
    assign weights1[50][566] = 16'b1111111111111011;
    assign weights1[50][567] = 16'b0000000000000001;
    assign weights1[50][568] = 16'b0000000000001000;
    assign weights1[50][569] = 16'b0000000000010011;
    assign weights1[50][570] = 16'b1111111111101101;
    assign weights1[50][571] = 16'b0000000000000011;
    assign weights1[50][572] = 16'b0000000000001100;
    assign weights1[50][573] = 16'b1111111111110110;
    assign weights1[50][574] = 16'b0000000000000110;
    assign weights1[50][575] = 16'b0000000000000101;
    assign weights1[50][576] = 16'b0000000000000110;
    assign weights1[50][577] = 16'b1111111111111111;
    assign weights1[50][578] = 16'b1111111111111111;
    assign weights1[50][579] = 16'b0000000000001010;
    assign weights1[50][580] = 16'b1111111111110110;
    assign weights1[50][581] = 16'b1111111111111110;
    assign weights1[50][582] = 16'b0000000000011100;
    assign weights1[50][583] = 16'b0000000000011100;
    assign weights1[50][584] = 16'b1111111111110001;
    assign weights1[50][585] = 16'b0000000000000010;
    assign weights1[50][586] = 16'b1111111111110111;
    assign weights1[50][587] = 16'b1111111111110110;
    assign weights1[50][588] = 16'b1111111111111010;
    assign weights1[50][589] = 16'b1111111111111111;
    assign weights1[50][590] = 16'b0000000000000110;
    assign weights1[50][591] = 16'b0000000000001000;
    assign weights1[50][592] = 16'b1111111111111011;
    assign weights1[50][593] = 16'b0000000000000111;
    assign weights1[50][594] = 16'b0000000000010000;
    assign weights1[50][595] = 16'b1111111111101010;
    assign weights1[50][596] = 16'b1111111111111010;
    assign weights1[50][597] = 16'b0000000000000000;
    assign weights1[50][598] = 16'b1111111111111001;
    assign weights1[50][599] = 16'b0000000000000001;
    assign weights1[50][600] = 16'b0000000000000000;
    assign weights1[50][601] = 16'b0000000000000111;
    assign weights1[50][602] = 16'b0000000000000001;
    assign weights1[50][603] = 16'b1111111111111100;
    assign weights1[50][604] = 16'b1111111111111001;
    assign weights1[50][605] = 16'b0000000000000010;
    assign weights1[50][606] = 16'b1111111111111100;
    assign weights1[50][607] = 16'b1111111111111100;
    assign weights1[50][608] = 16'b0000000000010111;
    assign weights1[50][609] = 16'b1111111111111000;
    assign weights1[50][610] = 16'b1111111111110001;
    assign weights1[50][611] = 16'b1111111111110101;
    assign weights1[50][612] = 16'b1111111111101110;
    assign weights1[50][613] = 16'b0000000000001010;
    assign weights1[50][614] = 16'b1111111111100001;
    assign weights1[50][615] = 16'b1111111111110011;
    assign weights1[50][616] = 16'b1111111111111000;
    assign weights1[50][617] = 16'b0000000000000101;
    assign weights1[50][618] = 16'b0000000000000001;
    assign weights1[50][619] = 16'b1111111111111001;
    assign weights1[50][620] = 16'b1111111111111111;
    assign weights1[50][621] = 16'b1111111111111010;
    assign weights1[50][622] = 16'b1111111111111010;
    assign weights1[50][623] = 16'b1111111111110111;
    assign weights1[50][624] = 16'b0000000000001100;
    assign weights1[50][625] = 16'b1111111111111010;
    assign weights1[50][626] = 16'b1111111111111101;
    assign weights1[50][627] = 16'b1111111111111010;
    assign weights1[50][628] = 16'b1111111111110110;
    assign weights1[50][629] = 16'b1111111111110100;
    assign weights1[50][630] = 16'b1111111111111001;
    assign weights1[50][631] = 16'b0000000000000100;
    assign weights1[50][632] = 16'b0000000000000100;
    assign weights1[50][633] = 16'b0000000000000101;
    assign weights1[50][634] = 16'b1111111111111011;
    assign weights1[50][635] = 16'b0000000000010001;
    assign weights1[50][636] = 16'b1111111111110101;
    assign weights1[50][637] = 16'b1111111111111101;
    assign weights1[50][638] = 16'b1111111111111100;
    assign weights1[50][639] = 16'b1111111111111111;
    assign weights1[50][640] = 16'b1111111111111111;
    assign weights1[50][641] = 16'b0000000000000101;
    assign weights1[50][642] = 16'b1111111111110010;
    assign weights1[50][643] = 16'b0000000000000100;
    assign weights1[50][644] = 16'b0000000000000011;
    assign weights1[50][645] = 16'b1111111111111110;
    assign weights1[50][646] = 16'b1111111111111111;
    assign weights1[50][647] = 16'b0000000000001101;
    assign weights1[50][648] = 16'b0000000000000011;
    assign weights1[50][649] = 16'b0000000000000000;
    assign weights1[50][650] = 16'b0000000000000001;
    assign weights1[50][651] = 16'b1111111111111101;
    assign weights1[50][652] = 16'b1111111111110011;
    assign weights1[50][653] = 16'b0000000000000110;
    assign weights1[50][654] = 16'b0000000000000001;
    assign weights1[50][655] = 16'b0000000000011101;
    assign weights1[50][656] = 16'b0000000000001100;
    assign weights1[50][657] = 16'b1111111111111001;
    assign weights1[50][658] = 16'b1111111111111101;
    assign weights1[50][659] = 16'b0000000000000001;
    assign weights1[50][660] = 16'b1111111111101100;
    assign weights1[50][661] = 16'b1111111111110000;
    assign weights1[50][662] = 16'b1111111111101011;
    assign weights1[50][663] = 16'b0000000000000011;
    assign weights1[50][664] = 16'b0000000000001001;
    assign weights1[50][665] = 16'b1111111111110001;
    assign weights1[50][666] = 16'b1111111111101101;
    assign weights1[50][667] = 16'b0000000000000010;
    assign weights1[50][668] = 16'b1111111111101000;
    assign weights1[50][669] = 16'b1111111111111011;
    assign weights1[50][670] = 16'b1111111111110100;
    assign weights1[50][671] = 16'b1111111111110111;
    assign weights1[50][672] = 16'b1111111111111111;
    assign weights1[50][673] = 16'b0000000000000111;
    assign weights1[50][674] = 16'b0000000000001010;
    assign weights1[50][675] = 16'b0000000000001001;
    assign weights1[50][676] = 16'b1111111111110111;
    assign weights1[50][677] = 16'b0000000000000010;
    assign weights1[50][678] = 16'b1111111111110011;
    assign weights1[50][679] = 16'b1111111111110111;
    assign weights1[50][680] = 16'b0000000000001000;
    assign weights1[50][681] = 16'b1111111111101100;
    assign weights1[50][682] = 16'b1111111111111011;
    assign weights1[50][683] = 16'b1111111111110110;
    assign weights1[50][684] = 16'b0000000000001010;
    assign weights1[50][685] = 16'b1111111111110110;
    assign weights1[50][686] = 16'b1111111111111101;
    assign weights1[50][687] = 16'b0000000000000100;
    assign weights1[50][688] = 16'b0000000000000110;
    assign weights1[50][689] = 16'b0000000000001001;
    assign weights1[50][690] = 16'b1111111111101000;
    assign weights1[50][691] = 16'b0000000000010011;
    assign weights1[50][692] = 16'b1111111111110010;
    assign weights1[50][693] = 16'b1111111111110101;
    assign weights1[50][694] = 16'b1111111111110000;
    assign weights1[50][695] = 16'b1111111111110111;
    assign weights1[50][696] = 16'b1111111111100101;
    assign weights1[50][697] = 16'b1111111111101100;
    assign weights1[50][698] = 16'b1111111111110011;
    assign weights1[50][699] = 16'b1111111111111011;
    assign weights1[50][700] = 16'b1111111111111011;
    assign weights1[50][701] = 16'b0000000000000011;
    assign weights1[50][702] = 16'b1111111111110101;
    assign weights1[50][703] = 16'b0000000000001011;
    assign weights1[50][704] = 16'b1111111111111001;
    assign weights1[50][705] = 16'b0000000000010101;
    assign weights1[50][706] = 16'b1111111111111000;
    assign weights1[50][707] = 16'b1111111111111111;
    assign weights1[50][708] = 16'b1111111111111011;
    assign weights1[50][709] = 16'b1111111111101101;
    assign weights1[50][710] = 16'b1111111111111000;
    assign weights1[50][711] = 16'b1111111111110011;
    assign weights1[50][712] = 16'b1111111111101100;
    assign weights1[50][713] = 16'b1111111111110011;
    assign weights1[50][714] = 16'b1111111111110000;
    assign weights1[50][715] = 16'b0000000000000000;
    assign weights1[50][716] = 16'b0000000000000000;
    assign weights1[50][717] = 16'b0000000000000001;
    assign weights1[50][718] = 16'b0000000000000111;
    assign weights1[50][719] = 16'b1111111111111110;
    assign weights1[50][720] = 16'b0000000000000010;
    assign weights1[50][721] = 16'b1111111111110000;
    assign weights1[50][722] = 16'b1111111111101100;
    assign weights1[50][723] = 16'b1111111111110110;
    assign weights1[50][724] = 16'b1111111111101110;
    assign weights1[50][725] = 16'b1111111111110101;
    assign weights1[50][726] = 16'b1111111111110101;
    assign weights1[50][727] = 16'b1111111111111100;
    assign weights1[50][728] = 16'b1111111111111101;
    assign weights1[50][729] = 16'b1111111111111101;
    assign weights1[50][730] = 16'b1111111111111110;
    assign weights1[50][731] = 16'b1111111111111111;
    assign weights1[50][732] = 16'b1111111111111101;
    assign weights1[50][733] = 16'b0000000000000100;
    assign weights1[50][734] = 16'b1111111111111111;
    assign weights1[50][735] = 16'b1111111111111010;
    assign weights1[50][736] = 16'b0000000000001110;
    assign weights1[50][737] = 16'b0000000000000111;
    assign weights1[50][738] = 16'b0000000000000101;
    assign weights1[50][739] = 16'b1111111111111101;
    assign weights1[50][740] = 16'b0000000000000111;
    assign weights1[50][741] = 16'b0000000000001111;
    assign weights1[50][742] = 16'b1111111111101111;
    assign weights1[50][743] = 16'b1111111111111100;
    assign weights1[50][744] = 16'b1111111111101111;
    assign weights1[50][745] = 16'b1111111111101100;
    assign weights1[50][746] = 16'b1111111111111001;
    assign weights1[50][747] = 16'b1111111111101001;
    assign weights1[50][748] = 16'b1111111111110100;
    assign weights1[50][749] = 16'b1111111111101001;
    assign weights1[50][750] = 16'b1111111111101010;
    assign weights1[50][751] = 16'b1111111111110100;
    assign weights1[50][752] = 16'b1111111111111011;
    assign weights1[50][753] = 16'b1111111111111111;
    assign weights1[50][754] = 16'b1111111111111110;
    assign weights1[50][755] = 16'b0000000000000001;
    assign weights1[50][756] = 16'b1111111111111110;
    assign weights1[50][757] = 16'b1111111111111101;
    assign weights1[50][758] = 16'b0000000000000111;
    assign weights1[50][759] = 16'b0000000000001001;
    assign weights1[50][760] = 16'b0000000000000001;
    assign weights1[50][761] = 16'b0000000000001011;
    assign weights1[50][762] = 16'b1111111111111110;
    assign weights1[50][763] = 16'b0000000000000001;
    assign weights1[50][764] = 16'b0000000000000011;
    assign weights1[50][765] = 16'b0000000000000001;
    assign weights1[50][766] = 16'b1111111111101010;
    assign weights1[50][767] = 16'b1111111111011101;
    assign weights1[50][768] = 16'b1111111111100000;
    assign weights1[50][769] = 16'b1111111111011101;
    assign weights1[50][770] = 16'b1111111111011010;
    assign weights1[50][771] = 16'b1111111111011101;
    assign weights1[50][772] = 16'b1111111111100010;
    assign weights1[50][773] = 16'b1111111111011110;
    assign weights1[50][774] = 16'b1111111111011111;
    assign weights1[50][775] = 16'b1111111111100010;
    assign weights1[50][776] = 16'b1111111111101110;
    assign weights1[50][777] = 16'b1111111111101011;
    assign weights1[50][778] = 16'b1111111111110111;
    assign weights1[50][779] = 16'b1111111111111010;
    assign weights1[50][780] = 16'b0000000000000000;
    assign weights1[50][781] = 16'b0000000000000001;
    assign weights1[50][782] = 16'b0000000000000001;
    assign weights1[50][783] = 16'b0000000000000100;
    assign weights1[51][0] = 16'b0000000000000000;
    assign weights1[51][1] = 16'b0000000000000001;
    assign weights1[51][2] = 16'b0000000000000001;
    assign weights1[51][3] = 16'b1111111111111110;
    assign weights1[51][4] = 16'b0000000000000001;
    assign weights1[51][5] = 16'b1111111111110111;
    assign weights1[51][6] = 16'b1111111111110111;
    assign weights1[51][7] = 16'b1111111111110100;
    assign weights1[51][8] = 16'b1111111111101110;
    assign weights1[51][9] = 16'b1111111111110100;
    assign weights1[51][10] = 16'b1111111111110010;
    assign weights1[51][11] = 16'b1111111111111000;
    assign weights1[51][12] = 16'b1111111111111011;
    assign weights1[51][13] = 16'b1111111111111011;
    assign weights1[51][14] = 16'b1111111111110111;
    assign weights1[51][15] = 16'b1111111111110001;
    assign weights1[51][16] = 16'b1111111111111011;
    assign weights1[51][17] = 16'b1111111111110100;
    assign weights1[51][18] = 16'b1111111111111011;
    assign weights1[51][19] = 16'b1111111111111000;
    assign weights1[51][20] = 16'b1111111111111001;
    assign weights1[51][21] = 16'b1111111111111110;
    assign weights1[51][22] = 16'b1111111111111010;
    assign weights1[51][23] = 16'b0000000000000000;
    assign weights1[51][24] = 16'b0000000000000100;
    assign weights1[51][25] = 16'b0000000000000100;
    assign weights1[51][26] = 16'b0000000000000011;
    assign weights1[51][27] = 16'b0000000000000010;
    assign weights1[51][28] = 16'b0000000000000000;
    assign weights1[51][29] = 16'b0000000000000001;
    assign weights1[51][30] = 16'b1111111111111100;
    assign weights1[51][31] = 16'b1111111111111101;
    assign weights1[51][32] = 16'b1111111111110101;
    assign weights1[51][33] = 16'b1111111111111010;
    assign weights1[51][34] = 16'b1111111111110101;
    assign weights1[51][35] = 16'b1111111111110100;
    assign weights1[51][36] = 16'b1111111111110001;
    assign weights1[51][37] = 16'b1111111111101110;
    assign weights1[51][38] = 16'b1111111111111001;
    assign weights1[51][39] = 16'b1111111111111100;
    assign weights1[51][40] = 16'b1111111111111101;
    assign weights1[51][41] = 16'b1111111111111010;
    assign weights1[51][42] = 16'b1111111111110111;
    assign weights1[51][43] = 16'b1111111111101110;
    assign weights1[51][44] = 16'b1111111111110011;
    assign weights1[51][45] = 16'b1111111111111011;
    assign weights1[51][46] = 16'b1111111111111010;
    assign weights1[51][47] = 16'b1111111111110110;
    assign weights1[51][48] = 16'b1111111111110100;
    assign weights1[51][49] = 16'b1111111111101111;
    assign weights1[51][50] = 16'b1111111111110010;
    assign weights1[51][51] = 16'b1111111111111001;
    assign weights1[51][52] = 16'b1111111111111111;
    assign weights1[51][53] = 16'b1111111111111111;
    assign weights1[51][54] = 16'b0000000000000011;
    assign weights1[51][55] = 16'b0000000000000010;
    assign weights1[51][56] = 16'b0000000000000000;
    assign weights1[51][57] = 16'b1111111111111101;
    assign weights1[51][58] = 16'b1111111111111001;
    assign weights1[51][59] = 16'b1111111111111001;
    assign weights1[51][60] = 16'b0000000000000001;
    assign weights1[51][61] = 16'b1111111111111101;
    assign weights1[51][62] = 16'b1111111111110110;
    assign weights1[51][63] = 16'b1111111111111000;
    assign weights1[51][64] = 16'b1111111111111110;
    assign weights1[51][65] = 16'b0000000000000011;
    assign weights1[51][66] = 16'b1111111111110111;
    assign weights1[51][67] = 16'b1111111111110111;
    assign weights1[51][68] = 16'b1111111111111101;
    assign weights1[51][69] = 16'b1111111111110100;
    assign weights1[51][70] = 16'b1111111111101110;
    assign weights1[51][71] = 16'b1111111111101100;
    assign weights1[51][72] = 16'b1111111111101001;
    assign weights1[51][73] = 16'b1111111111110000;
    assign weights1[51][74] = 16'b1111111111110100;
    assign weights1[51][75] = 16'b1111111111110100;
    assign weights1[51][76] = 16'b1111111111101110;
    assign weights1[51][77] = 16'b1111111111101101;
    assign weights1[51][78] = 16'b1111111111110000;
    assign weights1[51][79] = 16'b1111111111110111;
    assign weights1[51][80] = 16'b1111111111110100;
    assign weights1[51][81] = 16'b1111111111111001;
    assign weights1[51][82] = 16'b1111111111111111;
    assign weights1[51][83] = 16'b0000000000000010;
    assign weights1[51][84] = 16'b1111111111111101;
    assign weights1[51][85] = 16'b1111111111110110;
    assign weights1[51][86] = 16'b1111111111110011;
    assign weights1[51][87] = 16'b1111111111110111;
    assign weights1[51][88] = 16'b1111111111111110;
    assign weights1[51][89] = 16'b0000000000000010;
    assign weights1[51][90] = 16'b0000000000000000;
    assign weights1[51][91] = 16'b1111111111111010;
    assign weights1[51][92] = 16'b0000000000000100;
    assign weights1[51][93] = 16'b0000000000000100;
    assign weights1[51][94] = 16'b1111111111110110;
    assign weights1[51][95] = 16'b1111111111111010;
    assign weights1[51][96] = 16'b0000000000000001;
    assign weights1[51][97] = 16'b0000000000000111;
    assign weights1[51][98] = 16'b0000000000000000;
    assign weights1[51][99] = 16'b1111111111110011;
    assign weights1[51][100] = 16'b1111111111110001;
    assign weights1[51][101] = 16'b1111111111100011;
    assign weights1[51][102] = 16'b1111111111101101;
    assign weights1[51][103] = 16'b1111111111111001;
    assign weights1[51][104] = 16'b0000000000000010;
    assign weights1[51][105] = 16'b1111111111110000;
    assign weights1[51][106] = 16'b1111111111111011;
    assign weights1[51][107] = 16'b1111111111111001;
    assign weights1[51][108] = 16'b1111111111110101;
    assign weights1[51][109] = 16'b1111111111111011;
    assign weights1[51][110] = 16'b0000000000000100;
    assign weights1[51][111] = 16'b1111111111111111;
    assign weights1[51][112] = 16'b1111111111111010;
    assign weights1[51][113] = 16'b1111111111110011;
    assign weights1[51][114] = 16'b1111111111110000;
    assign weights1[51][115] = 16'b1111111111110000;
    assign weights1[51][116] = 16'b0000000000000000;
    assign weights1[51][117] = 16'b0000000000000111;
    assign weights1[51][118] = 16'b0000000000000100;
    assign weights1[51][119] = 16'b0000000000000110;
    assign weights1[51][120] = 16'b0000000000001101;
    assign weights1[51][121] = 16'b0000000000000110;
    assign weights1[51][122] = 16'b1111111111111010;
    assign weights1[51][123] = 16'b1111111111110100;
    assign weights1[51][124] = 16'b1111111111111001;
    assign weights1[51][125] = 16'b1111111111111000;
    assign weights1[51][126] = 16'b1111111111110101;
    assign weights1[51][127] = 16'b1111111111101111;
    assign weights1[51][128] = 16'b0000000000000001;
    assign weights1[51][129] = 16'b1111111111111011;
    assign weights1[51][130] = 16'b1111111111111011;
    assign weights1[51][131] = 16'b1111111111111111;
    assign weights1[51][132] = 16'b0000000000000000;
    assign weights1[51][133] = 16'b1111111111111101;
    assign weights1[51][134] = 16'b0000000000000011;
    assign weights1[51][135] = 16'b0000000000000101;
    assign weights1[51][136] = 16'b1111111111111110;
    assign weights1[51][137] = 16'b1111111111111100;
    assign weights1[51][138] = 16'b1111111111111110;
    assign weights1[51][139] = 16'b0000000000000001;
    assign weights1[51][140] = 16'b1111111111111001;
    assign weights1[51][141] = 16'b1111111111110100;
    assign weights1[51][142] = 16'b1111111111101111;
    assign weights1[51][143] = 16'b1111111111110010;
    assign weights1[51][144] = 16'b1111111111111101;
    assign weights1[51][145] = 16'b1111111111111110;
    assign weights1[51][146] = 16'b0000000000010010;
    assign weights1[51][147] = 16'b0000000000010011;
    assign weights1[51][148] = 16'b0000000000010100;
    assign weights1[51][149] = 16'b1111111111111110;
    assign weights1[51][150] = 16'b1111111111110101;
    assign weights1[51][151] = 16'b1111111111110111;
    assign weights1[51][152] = 16'b1111111111110111;
    assign weights1[51][153] = 16'b1111111111111011;
    assign weights1[51][154] = 16'b0000000000000000;
    assign weights1[51][155] = 16'b0000000000001001;
    assign weights1[51][156] = 16'b0000000000000000;
    assign weights1[51][157] = 16'b0000000000000101;
    assign weights1[51][158] = 16'b0000000000001000;
    assign weights1[51][159] = 16'b0000000000001011;
    assign weights1[51][160] = 16'b0000000000001001;
    assign weights1[51][161] = 16'b1111111111111110;
    assign weights1[51][162] = 16'b1111111111111010;
    assign weights1[51][163] = 16'b0000000000000000;
    assign weights1[51][164] = 16'b0000000000001000;
    assign weights1[51][165] = 16'b0000000000000001;
    assign weights1[51][166] = 16'b0000000000000111;
    assign weights1[51][167] = 16'b0000000000000010;
    assign weights1[51][168] = 16'b1111111111111001;
    assign weights1[51][169] = 16'b1111111111111010;
    assign weights1[51][170] = 16'b1111111111110111;
    assign weights1[51][171] = 16'b1111111111110111;
    assign weights1[51][172] = 16'b1111111111111100;
    assign weights1[51][173] = 16'b0000000000010001;
    assign weights1[51][174] = 16'b0000000000011010;
    assign weights1[51][175] = 16'b0000000000011010;
    assign weights1[51][176] = 16'b0000000000010011;
    assign weights1[51][177] = 16'b0000000000000100;
    assign weights1[51][178] = 16'b1111111111110101;
    assign weights1[51][179] = 16'b0000000000000000;
    assign weights1[51][180] = 16'b0000000000000011;
    assign weights1[51][181] = 16'b0000000000000010;
    assign weights1[51][182] = 16'b1111111111110111;
    assign weights1[51][183] = 16'b1111111111111110;
    assign weights1[51][184] = 16'b0000000000000111;
    assign weights1[51][185] = 16'b0000000000000111;
    assign weights1[51][186] = 16'b0000000000010000;
    assign weights1[51][187] = 16'b0000000000010010;
    assign weights1[51][188] = 16'b0000000000010110;
    assign weights1[51][189] = 16'b0000000000010110;
    assign weights1[51][190] = 16'b0000000000011000;
    assign weights1[51][191] = 16'b0000000000001100;
    assign weights1[51][192] = 16'b0000000000001001;
    assign weights1[51][193] = 16'b0000000000001011;
    assign weights1[51][194] = 16'b0000000000001100;
    assign weights1[51][195] = 16'b0000000000000001;
    assign weights1[51][196] = 16'b1111111111111100;
    assign weights1[51][197] = 16'b1111111111111101;
    assign weights1[51][198] = 16'b1111111111111000;
    assign weights1[51][199] = 16'b1111111111111111;
    assign weights1[51][200] = 16'b0000000000001010;
    assign weights1[51][201] = 16'b0000000000001100;
    assign weights1[51][202] = 16'b0000000000011110;
    assign weights1[51][203] = 16'b0000000000100111;
    assign weights1[51][204] = 16'b0000000000010010;
    assign weights1[51][205] = 16'b0000000000001110;
    assign weights1[51][206] = 16'b0000000000001011;
    assign weights1[51][207] = 16'b0000000000001010;
    assign weights1[51][208] = 16'b0000000000000110;
    assign weights1[51][209] = 16'b0000000000001001;
    assign weights1[51][210] = 16'b0000000000000110;
    assign weights1[51][211] = 16'b0000000000001001;
    assign weights1[51][212] = 16'b0000000000001100;
    assign weights1[51][213] = 16'b0000000000001001;
    assign weights1[51][214] = 16'b0000000000001111;
    assign weights1[51][215] = 16'b0000000000011001;
    assign weights1[51][216] = 16'b0000000000010111;
    assign weights1[51][217] = 16'b0000000000010100;
    assign weights1[51][218] = 16'b0000000000011000;
    assign weights1[51][219] = 16'b0000000000011010;
    assign weights1[51][220] = 16'b0000000000010011;
    assign weights1[51][221] = 16'b0000000000010010;
    assign weights1[51][222] = 16'b0000000000001111;
    assign weights1[51][223] = 16'b0000000000001100;
    assign weights1[51][224] = 16'b1111111111111000;
    assign weights1[51][225] = 16'b1111111111111001;
    assign weights1[51][226] = 16'b1111111111111100;
    assign weights1[51][227] = 16'b0000000000000101;
    assign weights1[51][228] = 16'b0000000000000011;
    assign weights1[51][229] = 16'b0000000000010100;
    assign weights1[51][230] = 16'b0000000000011100;
    assign weights1[51][231] = 16'b0000000000011000;
    assign weights1[51][232] = 16'b0000000000011001;
    assign weights1[51][233] = 16'b0000000000100010;
    assign weights1[51][234] = 16'b0000000000001011;
    assign weights1[51][235] = 16'b1111111111110110;
    assign weights1[51][236] = 16'b0000000000000001;
    assign weights1[51][237] = 16'b0000000000011000;
    assign weights1[51][238] = 16'b0000000000010001;
    assign weights1[51][239] = 16'b0000000000001100;
    assign weights1[51][240] = 16'b0000000000001100;
    assign weights1[51][241] = 16'b0000000000001010;
    assign weights1[51][242] = 16'b0000000000011000;
    assign weights1[51][243] = 16'b0000000000010100;
    assign weights1[51][244] = 16'b0000000000010011;
    assign weights1[51][245] = 16'b0000000000010010;
    assign weights1[51][246] = 16'b0000000000011001;
    assign weights1[51][247] = 16'b0000000000010101;
    assign weights1[51][248] = 16'b0000000000011110;
    assign weights1[51][249] = 16'b0000000000010001;
    assign weights1[51][250] = 16'b0000000000001111;
    assign weights1[51][251] = 16'b0000000000011001;
    assign weights1[51][252] = 16'b1111111111111001;
    assign weights1[51][253] = 16'b1111111111111010;
    assign weights1[51][254] = 16'b0000000000000010;
    assign weights1[51][255] = 16'b0000000000010001;
    assign weights1[51][256] = 16'b0000000000000100;
    assign weights1[51][257] = 16'b0000000000010111;
    assign weights1[51][258] = 16'b0000000000100110;
    assign weights1[51][259] = 16'b0000000000100110;
    assign weights1[51][260] = 16'b0000000000010100;
    assign weights1[51][261] = 16'b0000000000001100;
    assign weights1[51][262] = 16'b0000000000000010;
    assign weights1[51][263] = 16'b0000000000000001;
    assign weights1[51][264] = 16'b0000000000001001;
    assign weights1[51][265] = 16'b0000000000001101;
    assign weights1[51][266] = 16'b0000000000001111;
    assign weights1[51][267] = 16'b0000000000001001;
    assign weights1[51][268] = 16'b0000000000000101;
    assign weights1[51][269] = 16'b0000000000001011;
    assign weights1[51][270] = 16'b0000000000010001;
    assign weights1[51][271] = 16'b0000000000011001;
    assign weights1[51][272] = 16'b0000000000011000;
    assign weights1[51][273] = 16'b0000000000011001;
    assign weights1[51][274] = 16'b0000000000011011;
    assign weights1[51][275] = 16'b0000000000010110;
    assign weights1[51][276] = 16'b0000000000011001;
    assign weights1[51][277] = 16'b0000000000001010;
    assign weights1[51][278] = 16'b0000000000001100;
    assign weights1[51][279] = 16'b0000000000010110;
    assign weights1[51][280] = 16'b1111111111111110;
    assign weights1[51][281] = 16'b0000000000000101;
    assign weights1[51][282] = 16'b0000000000001101;
    assign weights1[51][283] = 16'b0000000000000101;
    assign weights1[51][284] = 16'b0000000000000110;
    assign weights1[51][285] = 16'b0000000000011101;
    assign weights1[51][286] = 16'b0000000000100100;
    assign weights1[51][287] = 16'b0000000000011011;
    assign weights1[51][288] = 16'b0000000000010110;
    assign weights1[51][289] = 16'b0000000000000100;
    assign weights1[51][290] = 16'b1111111111110110;
    assign weights1[51][291] = 16'b0000000000000101;
    assign weights1[51][292] = 16'b0000000000001011;
    assign weights1[51][293] = 16'b0000000000010111;
    assign weights1[51][294] = 16'b0000000000010010;
    assign weights1[51][295] = 16'b1111111111111111;
    assign weights1[51][296] = 16'b0000000000000001;
    assign weights1[51][297] = 16'b0000000000001011;
    assign weights1[51][298] = 16'b0000000000000111;
    assign weights1[51][299] = 16'b0000000000011000;
    assign weights1[51][300] = 16'b0000000000011011;
    assign weights1[51][301] = 16'b0000000000011001;
    assign weights1[51][302] = 16'b0000000000010100;
    assign weights1[51][303] = 16'b0000000000010001;
    assign weights1[51][304] = 16'b0000000000010111;
    assign weights1[51][305] = 16'b0000000000000100;
    assign weights1[51][306] = 16'b0000000000010100;
    assign weights1[51][307] = 16'b0000000000001111;
    assign weights1[51][308] = 16'b1111111111111111;
    assign weights1[51][309] = 16'b0000000000000001;
    assign weights1[51][310] = 16'b0000000000000010;
    assign weights1[51][311] = 16'b0000000000000101;
    assign weights1[51][312] = 16'b0000000000001011;
    assign weights1[51][313] = 16'b0000000000001011;
    assign weights1[51][314] = 16'b0000000000010011;
    assign weights1[51][315] = 16'b0000000000100101;
    assign weights1[51][316] = 16'b0000000000011010;
    assign weights1[51][317] = 16'b0000000000000101;
    assign weights1[51][318] = 16'b1111111111111110;
    assign weights1[51][319] = 16'b0000000000000000;
    assign weights1[51][320] = 16'b0000000000000111;
    assign weights1[51][321] = 16'b0000000000000011;
    assign weights1[51][322] = 16'b1111111111111100;
    assign weights1[51][323] = 16'b1111111111111010;
    assign weights1[51][324] = 16'b1111111111111001;
    assign weights1[51][325] = 16'b1111111111111011;
    assign weights1[51][326] = 16'b1111111111110000;
    assign weights1[51][327] = 16'b1111111111111101;
    assign weights1[51][328] = 16'b0000000000001010;
    assign weights1[51][329] = 16'b0000000000011001;
    assign weights1[51][330] = 16'b0000000000011010;
    assign weights1[51][331] = 16'b0000000000011011;
    assign weights1[51][332] = 16'b0000000000001101;
    assign weights1[51][333] = 16'b0000000000000100;
    assign weights1[51][334] = 16'b0000000000001010;
    assign weights1[51][335] = 16'b0000000000001101;
    assign weights1[51][336] = 16'b1111111111111110;
    assign weights1[51][337] = 16'b0000000000000110;
    assign weights1[51][338] = 16'b0000000000001011;
    assign weights1[51][339] = 16'b0000000000001111;
    assign weights1[51][340] = 16'b0000000000001011;
    assign weights1[51][341] = 16'b0000000000001011;
    assign weights1[51][342] = 16'b0000000000011111;
    assign weights1[51][343] = 16'b0000000000011010;
    assign weights1[51][344] = 16'b0000000000001111;
    assign weights1[51][345] = 16'b1111111111110101;
    assign weights1[51][346] = 16'b1111111111110011;
    assign weights1[51][347] = 16'b0000000000000000;
    assign weights1[51][348] = 16'b0000000000000010;
    assign weights1[51][349] = 16'b0000000000001101;
    assign weights1[51][350] = 16'b1111111111111100;
    assign weights1[51][351] = 16'b1111111111110000;
    assign weights1[51][352] = 16'b1111111111100111;
    assign weights1[51][353] = 16'b1111111111101010;
    assign weights1[51][354] = 16'b1111111111101110;
    assign weights1[51][355] = 16'b1111111111110010;
    assign weights1[51][356] = 16'b0000000000001100;
    assign weights1[51][357] = 16'b0000000000010001;
    assign weights1[51][358] = 16'b0000000000100000;
    assign weights1[51][359] = 16'b0000000000100101;
    assign weights1[51][360] = 16'b0000000000011111;
    assign weights1[51][361] = 16'b0000000000001101;
    assign weights1[51][362] = 16'b0000000000001100;
    assign weights1[51][363] = 16'b0000000000001010;
    assign weights1[51][364] = 16'b0000000000000010;
    assign weights1[51][365] = 16'b0000000000000011;
    assign weights1[51][366] = 16'b0000000000000110;
    assign weights1[51][367] = 16'b0000000000010100;
    assign weights1[51][368] = 16'b0000000000011001;
    assign weights1[51][369] = 16'b0000000000010111;
    assign weights1[51][370] = 16'b0000000000100100;
    assign weights1[51][371] = 16'b0000000000010011;
    assign weights1[51][372] = 16'b0000000000001110;
    assign weights1[51][373] = 16'b0000000000000001;
    assign weights1[51][374] = 16'b1111111111110000;
    assign weights1[51][375] = 16'b1111111111110110;
    assign weights1[51][376] = 16'b0000000000000000;
    assign weights1[51][377] = 16'b0000000000000001;
    assign weights1[51][378] = 16'b1111111111101010;
    assign weights1[51][379] = 16'b1111111111101010;
    assign weights1[51][380] = 16'b1111111111101000;
    assign weights1[51][381] = 16'b1111111111011111;
    assign weights1[51][382] = 16'b1111111111011101;
    assign weights1[51][383] = 16'b1111111111101111;
    assign weights1[51][384] = 16'b1111111111111101;
    assign weights1[51][385] = 16'b0000000000010100;
    assign weights1[51][386] = 16'b0000000000010101;
    assign weights1[51][387] = 16'b0000000000100000;
    assign weights1[51][388] = 16'b0000000000011011;
    assign weights1[51][389] = 16'b0000000000011010;
    assign weights1[51][390] = 16'b0000000000001010;
    assign weights1[51][391] = 16'b0000000000001101;
    assign weights1[51][392] = 16'b1111111111111111;
    assign weights1[51][393] = 16'b0000000000000011;
    assign weights1[51][394] = 16'b1111111111111011;
    assign weights1[51][395] = 16'b0000000000001100;
    assign weights1[51][396] = 16'b0000000000010011;
    assign weights1[51][397] = 16'b0000000000011101;
    assign weights1[51][398] = 16'b0000000000011010;
    assign weights1[51][399] = 16'b0000000000010100;
    assign weights1[51][400] = 16'b0000000000000100;
    assign weights1[51][401] = 16'b0000000000000010;
    assign weights1[51][402] = 16'b1111111111110000;
    assign weights1[51][403] = 16'b1111111111100101;
    assign weights1[51][404] = 16'b1111111111110000;
    assign weights1[51][405] = 16'b1111111111101101;
    assign weights1[51][406] = 16'b1111111111101111;
    assign weights1[51][407] = 16'b1111111111101100;
    assign weights1[51][408] = 16'b1111111111101011;
    assign weights1[51][409] = 16'b1111111111101111;
    assign weights1[51][410] = 16'b1111111111101100;
    assign weights1[51][411] = 16'b1111111111101010;
    assign weights1[51][412] = 16'b1111111111101011;
    assign weights1[51][413] = 16'b0000000000000100;
    assign weights1[51][414] = 16'b0000000000100011;
    assign weights1[51][415] = 16'b0000000000100010;
    assign weights1[51][416] = 16'b0000000000100001;
    assign weights1[51][417] = 16'b0000000000010011;
    assign weights1[51][418] = 16'b0000000000010110;
    assign weights1[51][419] = 16'b0000000000010001;
    assign weights1[51][420] = 16'b1111111111111001;
    assign weights1[51][421] = 16'b1111111111111001;
    assign weights1[51][422] = 16'b0000000000000110;
    assign weights1[51][423] = 16'b0000000000000100;
    assign weights1[51][424] = 16'b0000000000001010;
    assign weights1[51][425] = 16'b0000000000011100;
    assign weights1[51][426] = 16'b0000000000011111;
    assign weights1[51][427] = 16'b0000000000011000;
    assign weights1[51][428] = 16'b0000000000000111;
    assign weights1[51][429] = 16'b1111111111101110;
    assign weights1[51][430] = 16'b1111111111101111;
    assign weights1[51][431] = 16'b1111111111101001;
    assign weights1[51][432] = 16'b1111111111101101;
    assign weights1[51][433] = 16'b1111111111110010;
    assign weights1[51][434] = 16'b1111111111110011;
    assign weights1[51][435] = 16'b1111111111110001;
    assign weights1[51][436] = 16'b1111111111110011;
    assign weights1[51][437] = 16'b1111111111100001;
    assign weights1[51][438] = 16'b1111111111101001;
    assign weights1[51][439] = 16'b1111111111100111;
    assign weights1[51][440] = 16'b1111111111100101;
    assign weights1[51][441] = 16'b0000000000000000;
    assign weights1[51][442] = 16'b0000000000001110;
    assign weights1[51][443] = 16'b0000000000011001;
    assign weights1[51][444] = 16'b0000000000011010;
    assign weights1[51][445] = 16'b0000000000011001;
    assign weights1[51][446] = 16'b0000000000001110;
    assign weights1[51][447] = 16'b0000000000001101;
    assign weights1[51][448] = 16'b1111111111110110;
    assign weights1[51][449] = 16'b1111111111110111;
    assign weights1[51][450] = 16'b1111111111111111;
    assign weights1[51][451] = 16'b1111111111110011;
    assign weights1[51][452] = 16'b1111111111111111;
    assign weights1[51][453] = 16'b0000000000010000;
    assign weights1[51][454] = 16'b0000000000010001;
    assign weights1[51][455] = 16'b0000000000001110;
    assign weights1[51][456] = 16'b1111111111111110;
    assign weights1[51][457] = 16'b1111111111110001;
    assign weights1[51][458] = 16'b1111111111101111;
    assign weights1[51][459] = 16'b1111111111110100;
    assign weights1[51][460] = 16'b1111111111110111;
    assign weights1[51][461] = 16'b1111111111111100;
    assign weights1[51][462] = 16'b1111111111111101;
    assign weights1[51][463] = 16'b0000000000000000;
    assign weights1[51][464] = 16'b1111111111101111;
    assign weights1[51][465] = 16'b1111111111101011;
    assign weights1[51][466] = 16'b1111111111101000;
    assign weights1[51][467] = 16'b1111111111010111;
    assign weights1[51][468] = 16'b1111111111101100;
    assign weights1[51][469] = 16'b1111111111111110;
    assign weights1[51][470] = 16'b0000000000001000;
    assign weights1[51][471] = 16'b0000000000010011;
    assign weights1[51][472] = 16'b0000000000011001;
    assign weights1[51][473] = 16'b0000000000001010;
    assign weights1[51][474] = 16'b0000000000000110;
    assign weights1[51][475] = 16'b0000000000001011;
    assign weights1[51][476] = 16'b1111111111111100;
    assign weights1[51][477] = 16'b1111111111110100;
    assign weights1[51][478] = 16'b1111111111110111;
    assign weights1[51][479] = 16'b1111111111110010;
    assign weights1[51][480] = 16'b1111111111111011;
    assign weights1[51][481] = 16'b0000000000000111;
    assign weights1[51][482] = 16'b0000000000001010;
    assign weights1[51][483] = 16'b0000000000010001;
    assign weights1[51][484] = 16'b0000000000001000;
    assign weights1[51][485] = 16'b0000000000001000;
    assign weights1[51][486] = 16'b0000000000000000;
    assign weights1[51][487] = 16'b0000000000000000;
    assign weights1[51][488] = 16'b1111111111101111;
    assign weights1[51][489] = 16'b1111111111110101;
    assign weights1[51][490] = 16'b0000000000000100;
    assign weights1[51][491] = 16'b0000000000001100;
    assign weights1[51][492] = 16'b1111111111111010;
    assign weights1[51][493] = 16'b1111111111100001;
    assign weights1[51][494] = 16'b1111111111100101;
    assign weights1[51][495] = 16'b1111111111100001;
    assign weights1[51][496] = 16'b1111111111101011;
    assign weights1[51][497] = 16'b1111111111110111;
    assign weights1[51][498] = 16'b0000000000010001;
    assign weights1[51][499] = 16'b0000000000010011;
    assign weights1[51][500] = 16'b0000000000100001;
    assign weights1[51][501] = 16'b1111111111111110;
    assign weights1[51][502] = 16'b0000000000000010;
    assign weights1[51][503] = 16'b0000000000001000;
    assign weights1[51][504] = 16'b1111111111110101;
    assign weights1[51][505] = 16'b1111111111110100;
    assign weights1[51][506] = 16'b1111111111111011;
    assign weights1[51][507] = 16'b1111111111110000;
    assign weights1[51][508] = 16'b1111111111110000;
    assign weights1[51][509] = 16'b1111111111111100;
    assign weights1[51][510] = 16'b0000000000001100;
    assign weights1[51][511] = 16'b0000000000001010;
    assign weights1[51][512] = 16'b0000000000001110;
    assign weights1[51][513] = 16'b0000000000001101;
    assign weights1[51][514] = 16'b0000000000000011;
    assign weights1[51][515] = 16'b1111111111111011;
    assign weights1[51][516] = 16'b0000000000000001;
    assign weights1[51][517] = 16'b0000000000001000;
    assign weights1[51][518] = 16'b0000000000001011;
    assign weights1[51][519] = 16'b0000000000000001;
    assign weights1[51][520] = 16'b0000000000000100;
    assign weights1[51][521] = 16'b1111111111100111;
    assign weights1[51][522] = 16'b1111111111011000;
    assign weights1[51][523] = 16'b1111111111010111;
    assign weights1[51][524] = 16'b1111111111101000;
    assign weights1[51][525] = 16'b1111111111111001;
    assign weights1[51][526] = 16'b0000000000001011;
    assign weights1[51][527] = 16'b0000000000011000;
    assign weights1[51][528] = 16'b0000000000010101;
    assign weights1[51][529] = 16'b0000000000000101;
    assign weights1[51][530] = 16'b0000000000001001;
    assign weights1[51][531] = 16'b0000000000000011;
    assign weights1[51][532] = 16'b1111111111110100;
    assign weights1[51][533] = 16'b1111111111101100;
    assign weights1[51][534] = 16'b1111111111110011;
    assign weights1[51][535] = 16'b1111111111101111;
    assign weights1[51][536] = 16'b1111111111101101;
    assign weights1[51][537] = 16'b0000000000000001;
    assign weights1[51][538] = 16'b0000000000001110;
    assign weights1[51][539] = 16'b0000000000011001;
    assign weights1[51][540] = 16'b0000000000010111;
    assign weights1[51][541] = 16'b0000000000001001;
    assign weights1[51][542] = 16'b1111111111111100;
    assign weights1[51][543] = 16'b1111111111111000;
    assign weights1[51][544] = 16'b1111111111111000;
    assign weights1[51][545] = 16'b0000000000001010;
    assign weights1[51][546] = 16'b0000000000010010;
    assign weights1[51][547] = 16'b0000000000010010;
    assign weights1[51][548] = 16'b0000000000001011;
    assign weights1[51][549] = 16'b1111111111101000;
    assign weights1[51][550] = 16'b1111111111011001;
    assign weights1[51][551] = 16'b1111111111100100;
    assign weights1[51][552] = 16'b1111111111110100;
    assign weights1[51][553] = 16'b1111111111110101;
    assign weights1[51][554] = 16'b0000000000000110;
    assign weights1[51][555] = 16'b0000000000001110;
    assign weights1[51][556] = 16'b0000000000010001;
    assign weights1[51][557] = 16'b0000000000000110;
    assign weights1[51][558] = 16'b0000000000000010;
    assign weights1[51][559] = 16'b1111111111110110;
    assign weights1[51][560] = 16'b1111111111110100;
    assign weights1[51][561] = 16'b1111111111110001;
    assign weights1[51][562] = 16'b1111111111110110;
    assign weights1[51][563] = 16'b1111111111101111;
    assign weights1[51][564] = 16'b1111111111110001;
    assign weights1[51][565] = 16'b0000000000000001;
    assign weights1[51][566] = 16'b0000000000001001;
    assign weights1[51][567] = 16'b0000000000010100;
    assign weights1[51][568] = 16'b0000000000001100;
    assign weights1[51][569] = 16'b0000000000001010;
    assign weights1[51][570] = 16'b1111111111111100;
    assign weights1[51][571] = 16'b1111111111110111;
    assign weights1[51][572] = 16'b1111111111111001;
    assign weights1[51][573] = 16'b0000000000001001;
    assign weights1[51][574] = 16'b0000000000001000;
    assign weights1[51][575] = 16'b0000000000010010;
    assign weights1[51][576] = 16'b1111111111111011;
    assign weights1[51][577] = 16'b1111111111011011;
    assign weights1[51][578] = 16'b1111111111101000;
    assign weights1[51][579] = 16'b1111111111100111;
    assign weights1[51][580] = 16'b1111111111110100;
    assign weights1[51][581] = 16'b1111111111110111;
    assign weights1[51][582] = 16'b0000000000000000;
    assign weights1[51][583] = 16'b0000000000001101;
    assign weights1[51][584] = 16'b0000000000010001;
    assign weights1[51][585] = 16'b0000000000000110;
    assign weights1[51][586] = 16'b1111111111111101;
    assign weights1[51][587] = 16'b1111111111111010;
    assign weights1[51][588] = 16'b1111111111110101;
    assign weights1[51][589] = 16'b1111111111111000;
    assign weights1[51][590] = 16'b1111111111110110;
    assign weights1[51][591] = 16'b1111111111111101;
    assign weights1[51][592] = 16'b1111111111110111;
    assign weights1[51][593] = 16'b1111111111110001;
    assign weights1[51][594] = 16'b1111111111110001;
    assign weights1[51][595] = 16'b0000000000001000;
    assign weights1[51][596] = 16'b0000000000001110;
    assign weights1[51][597] = 16'b0000000000011001;
    assign weights1[51][598] = 16'b0000000000000010;
    assign weights1[51][599] = 16'b1111111111110101;
    assign weights1[51][600] = 16'b0000000000000110;
    assign weights1[51][601] = 16'b0000000000000101;
    assign weights1[51][602] = 16'b0000000000000000;
    assign weights1[51][603] = 16'b0000000000001010;
    assign weights1[51][604] = 16'b1111111111100111;
    assign weights1[51][605] = 16'b1111111111010100;
    assign weights1[51][606] = 16'b1111111111011011;
    assign weights1[51][607] = 16'b1111111111110110;
    assign weights1[51][608] = 16'b0000000000000001;
    assign weights1[51][609] = 16'b1111111111111011;
    assign weights1[51][610] = 16'b1111111111111000;
    assign weights1[51][611] = 16'b0000000000000100;
    assign weights1[51][612] = 16'b0000000000001000;
    assign weights1[51][613] = 16'b1111111111111111;
    assign weights1[51][614] = 16'b1111111111110101;
    assign weights1[51][615] = 16'b1111111111110111;
    assign weights1[51][616] = 16'b0000000000000010;
    assign weights1[51][617] = 16'b1111111111111001;
    assign weights1[51][618] = 16'b1111111111110110;
    assign weights1[51][619] = 16'b1111111111101111;
    assign weights1[51][620] = 16'b1111111111100111;
    assign weights1[51][621] = 16'b1111111111101111;
    assign weights1[51][622] = 16'b1111111111111100;
    assign weights1[51][623] = 16'b0000000000001000;
    assign weights1[51][624] = 16'b0000000000001110;
    assign weights1[51][625] = 16'b0000000000010011;
    assign weights1[51][626] = 16'b0000000000010111;
    assign weights1[51][627] = 16'b0000000000001001;
    assign weights1[51][628] = 16'b0000000000000011;
    assign weights1[51][629] = 16'b0000000000000111;
    assign weights1[51][630] = 16'b0000000000000000;
    assign weights1[51][631] = 16'b1111111111110001;
    assign weights1[51][632] = 16'b1111111111101111;
    assign weights1[51][633] = 16'b1111111111100110;
    assign weights1[51][634] = 16'b1111111111101111;
    assign weights1[51][635] = 16'b1111111111111100;
    assign weights1[51][636] = 16'b1111111111111001;
    assign weights1[51][637] = 16'b1111111111110100;
    assign weights1[51][638] = 16'b1111111111111000;
    assign weights1[51][639] = 16'b1111111111110111;
    assign weights1[51][640] = 16'b1111111111111000;
    assign weights1[51][641] = 16'b1111111111111011;
    assign weights1[51][642] = 16'b1111111111110100;
    assign weights1[51][643] = 16'b1111111111111001;
    assign weights1[51][644] = 16'b0000000000000001;
    assign weights1[51][645] = 16'b1111111111111011;
    assign weights1[51][646] = 16'b1111111111110100;
    assign weights1[51][647] = 16'b1111111111111000;
    assign weights1[51][648] = 16'b1111111111101110;
    assign weights1[51][649] = 16'b1111111111101111;
    assign weights1[51][650] = 16'b1111111111101100;
    assign weights1[51][651] = 16'b1111111111101110;
    assign weights1[51][652] = 16'b1111111111110001;
    assign weights1[51][653] = 16'b0000000000000010;
    assign weights1[51][654] = 16'b0000000000001011;
    assign weights1[51][655] = 16'b0000000000010100;
    assign weights1[51][656] = 16'b0000000000001100;
    assign weights1[51][657] = 16'b1111111111111111;
    assign weights1[51][658] = 16'b1111111111110010;
    assign weights1[51][659] = 16'b1111111111110010;
    assign weights1[51][660] = 16'b1111111111111000;
    assign weights1[51][661] = 16'b1111111111110010;
    assign weights1[51][662] = 16'b1111111111110000;
    assign weights1[51][663] = 16'b0000000000000011;
    assign weights1[51][664] = 16'b1111111111111001;
    assign weights1[51][665] = 16'b1111111111110101;
    assign weights1[51][666] = 16'b1111111111101100;
    assign weights1[51][667] = 16'b1111111111101000;
    assign weights1[51][668] = 16'b1111111111101101;
    assign weights1[51][669] = 16'b1111111111110100;
    assign weights1[51][670] = 16'b1111111111110111;
    assign weights1[51][671] = 16'b1111111111111011;
    assign weights1[51][672] = 16'b1111111111111100;
    assign weights1[51][673] = 16'b0000000000000001;
    assign weights1[51][674] = 16'b1111111111110111;
    assign weights1[51][675] = 16'b1111111111111100;
    assign weights1[51][676] = 16'b1111111111110110;
    assign weights1[51][677] = 16'b1111111111110010;
    assign weights1[51][678] = 16'b1111111111100110;
    assign weights1[51][679] = 16'b1111111111011001;
    assign weights1[51][680] = 16'b1111111111100110;
    assign weights1[51][681] = 16'b1111111111101011;
    assign weights1[51][682] = 16'b1111111111111110;
    assign weights1[51][683] = 16'b0000000000000111;
    assign weights1[51][684] = 16'b0000000000000100;
    assign weights1[51][685] = 16'b1111111111111010;
    assign weights1[51][686] = 16'b1111111111110111;
    assign weights1[51][687] = 16'b1111111111110110;
    assign weights1[51][688] = 16'b1111111111111011;
    assign weights1[51][689] = 16'b1111111111101100;
    assign weights1[51][690] = 16'b1111111111110010;
    assign weights1[51][691] = 16'b1111111111111101;
    assign weights1[51][692] = 16'b1111111111110011;
    assign weights1[51][693] = 16'b1111111111100011;
    assign weights1[51][694] = 16'b1111111111101001;
    assign weights1[51][695] = 16'b1111111111101011;
    assign weights1[51][696] = 16'b1111111111110010;
    assign weights1[51][697] = 16'b1111111111101011;
    assign weights1[51][698] = 16'b1111111111111111;
    assign weights1[51][699] = 16'b1111111111111011;
    assign weights1[51][700] = 16'b1111111111111110;
    assign weights1[51][701] = 16'b1111111111111110;
    assign weights1[51][702] = 16'b1111111111111110;
    assign weights1[51][703] = 16'b1111111111111011;
    assign weights1[51][704] = 16'b1111111111111001;
    assign weights1[51][705] = 16'b1111111111110100;
    assign weights1[51][706] = 16'b1111111111110000;
    assign weights1[51][707] = 16'b1111111111111000;
    assign weights1[51][708] = 16'b1111111111110001;
    assign weights1[51][709] = 16'b1111111111101000;
    assign weights1[51][710] = 16'b1111111111101001;
    assign weights1[51][711] = 16'b1111111111101010;
    assign weights1[51][712] = 16'b1111111111101001;
    assign weights1[51][713] = 16'b1111111111100111;
    assign weights1[51][714] = 16'b1111111111110011;
    assign weights1[51][715] = 16'b1111111111111011;
    assign weights1[51][716] = 16'b1111111111111101;
    assign weights1[51][717] = 16'b1111111111110110;
    assign weights1[51][718] = 16'b1111111111110101;
    assign weights1[51][719] = 16'b1111111111110110;
    assign weights1[51][720] = 16'b1111111111101000;
    assign weights1[51][721] = 16'b1111111111101101;
    assign weights1[51][722] = 16'b1111111111101101;
    assign weights1[51][723] = 16'b1111111111110000;
    assign weights1[51][724] = 16'b1111111111100101;
    assign weights1[51][725] = 16'b1111111111110000;
    assign weights1[51][726] = 16'b1111111111111011;
    assign weights1[51][727] = 16'b1111111111111100;
    assign weights1[51][728] = 16'b0000000000000000;
    assign weights1[51][729] = 16'b1111111111111011;
    assign weights1[51][730] = 16'b1111111111111000;
    assign weights1[51][731] = 16'b1111111111110111;
    assign weights1[51][732] = 16'b1111111111111011;
    assign weights1[51][733] = 16'b0000000000000011;
    assign weights1[51][734] = 16'b1111111111111111;
    assign weights1[51][735] = 16'b0000000000000010;
    assign weights1[51][736] = 16'b0000000000000100;
    assign weights1[51][737] = 16'b1111111111111100;
    assign weights1[51][738] = 16'b1111111111110001;
    assign weights1[51][739] = 16'b1111111111111100;
    assign weights1[51][740] = 16'b1111111111111000;
    assign weights1[51][741] = 16'b1111111111111010;
    assign weights1[51][742] = 16'b1111111111110111;
    assign weights1[51][743] = 16'b1111111111111111;
    assign weights1[51][744] = 16'b0000000000000011;
    assign weights1[51][745] = 16'b1111111111111100;
    assign weights1[51][746] = 16'b1111111111110100;
    assign weights1[51][747] = 16'b1111111111110011;
    assign weights1[51][748] = 16'b1111111111100111;
    assign weights1[51][749] = 16'b1111111111100111;
    assign weights1[51][750] = 16'b1111111111101110;
    assign weights1[51][751] = 16'b1111111111101101;
    assign weights1[51][752] = 16'b1111111111101110;
    assign weights1[51][753] = 16'b1111111111110100;
    assign weights1[51][754] = 16'b1111111111111001;
    assign weights1[51][755] = 16'b1111111111111101;
    assign weights1[51][756] = 16'b1111111111111110;
    assign weights1[51][757] = 16'b1111111111111010;
    assign weights1[51][758] = 16'b1111111111111001;
    assign weights1[51][759] = 16'b1111111111110101;
    assign weights1[51][760] = 16'b1111111111110000;
    assign weights1[51][761] = 16'b1111111111110110;
    assign weights1[51][762] = 16'b1111111111111010;
    assign weights1[51][763] = 16'b1111111111111111;
    assign weights1[51][764] = 16'b1111111111111000;
    assign weights1[51][765] = 16'b0000000000000000;
    assign weights1[51][766] = 16'b1111111111111011;
    assign weights1[51][767] = 16'b0000000000000111;
    assign weights1[51][768] = 16'b0000000000000000;
    assign weights1[51][769] = 16'b0000000000000010;
    assign weights1[51][770] = 16'b0000000000000010;
    assign weights1[51][771] = 16'b0000000000001111;
    assign weights1[51][772] = 16'b0000000000001001;
    assign weights1[51][773] = 16'b1111111111111011;
    assign weights1[51][774] = 16'b1111111111111000;
    assign weights1[51][775] = 16'b1111111111110010;
    assign weights1[51][776] = 16'b1111111111101000;
    assign weights1[51][777] = 16'b1111111111101010;
    assign weights1[51][778] = 16'b1111111111101101;
    assign weights1[51][779] = 16'b1111111111110000;
    assign weights1[51][780] = 16'b1111111111110101;
    assign weights1[51][781] = 16'b1111111111111100;
    assign weights1[51][782] = 16'b1111111111111101;
    assign weights1[51][783] = 16'b1111111111111110;
    assign weights1[52][0] = 16'b1111111111111111;
    assign weights1[52][1] = 16'b1111111111111111;
    assign weights1[52][2] = 16'b1111111111111111;
    assign weights1[52][3] = 16'b1111111111111111;
    assign weights1[52][4] = 16'b0000000000000001;
    assign weights1[52][5] = 16'b0000000000000011;
    assign weights1[52][6] = 16'b0000000000000010;
    assign weights1[52][7] = 16'b0000000000000100;
    assign weights1[52][8] = 16'b0000000000010011;
    assign weights1[52][9] = 16'b0000000000011010;
    assign weights1[52][10] = 16'b0000000000100101;
    assign weights1[52][11] = 16'b0000000000110101;
    assign weights1[52][12] = 16'b0000000000111000;
    assign weights1[52][13] = 16'b0000000001000100;
    assign weights1[52][14] = 16'b0000000001001111;
    assign weights1[52][15] = 16'b0000000001001001;
    assign weights1[52][16] = 16'b0000000000110010;
    assign weights1[52][17] = 16'b0000000000101100;
    assign weights1[52][18] = 16'b0000000000100010;
    assign weights1[52][19] = 16'b0000000000100111;
    assign weights1[52][20] = 16'b0000000000100001;
    assign weights1[52][21] = 16'b0000000000010111;
    assign weights1[52][22] = 16'b0000000000010000;
    assign weights1[52][23] = 16'b0000000000010010;
    assign weights1[52][24] = 16'b0000000000001100;
    assign weights1[52][25] = 16'b0000000000000111;
    assign weights1[52][26] = 16'b0000000000000101;
    assign weights1[52][27] = 16'b0000000000000001;
    assign weights1[52][28] = 16'b0000000000000000;
    assign weights1[52][29] = 16'b1111111111111111;
    assign weights1[52][30] = 16'b1111111111111111;
    assign weights1[52][31] = 16'b1111111111111111;
    assign weights1[52][32] = 16'b1111111111111111;
    assign weights1[52][33] = 16'b1111111111111001;
    assign weights1[52][34] = 16'b1111111111111011;
    assign weights1[52][35] = 16'b0000000000000111;
    assign weights1[52][36] = 16'b0000000000010111;
    assign weights1[52][37] = 16'b0000000000011000;
    assign weights1[52][38] = 16'b0000000000100010;
    assign weights1[52][39] = 16'b0000000000101010;
    assign weights1[52][40] = 16'b0000000001000011;
    assign weights1[52][41] = 16'b0000000001010000;
    assign weights1[52][42] = 16'b0000000001000110;
    assign weights1[52][43] = 16'b0000000000111011;
    assign weights1[52][44] = 16'b0000000000110010;
    assign weights1[52][45] = 16'b0000000000111111;
    assign weights1[52][46] = 16'b0000000000100010;
    assign weights1[52][47] = 16'b0000000000011011;
    assign weights1[52][48] = 16'b0000000000011100;
    assign weights1[52][49] = 16'b0000000000011110;
    assign weights1[52][50] = 16'b0000000000011010;
    assign weights1[52][51] = 16'b0000000000011011;
    assign weights1[52][52] = 16'b0000000000001111;
    assign weights1[52][53] = 16'b0000000000001110;
    assign weights1[52][54] = 16'b0000000000001010;
    assign weights1[52][55] = 16'b0000000000000100;
    assign weights1[52][56] = 16'b1111111111111111;
    assign weights1[52][57] = 16'b1111111111111111;
    assign weights1[52][58] = 16'b1111111111111110;
    assign weights1[52][59] = 16'b1111111111111011;
    assign weights1[52][60] = 16'b1111111111111011;
    assign weights1[52][61] = 16'b1111111111110101;
    assign weights1[52][62] = 16'b1111111111110101;
    assign weights1[52][63] = 16'b1111111111111111;
    assign weights1[52][64] = 16'b0000000000000011;
    assign weights1[52][65] = 16'b1111111111111110;
    assign weights1[52][66] = 16'b0000000000001001;
    assign weights1[52][67] = 16'b0000000000001110;
    assign weights1[52][68] = 16'b0000000000010110;
    assign weights1[52][69] = 16'b0000000000111010;
    assign weights1[52][70] = 16'b0000000000101111;
    assign weights1[52][71] = 16'b0000000000111011;
    assign weights1[52][72] = 16'b0000000000111111;
    assign weights1[52][73] = 16'b0000000000110101;
    assign weights1[52][74] = 16'b0000000000100010;
    assign weights1[52][75] = 16'b0000000000101000;
    assign weights1[52][76] = 16'b0000000000011110;
    assign weights1[52][77] = 16'b0000000000110011;
    assign weights1[52][78] = 16'b0000000000010011;
    assign weights1[52][79] = 16'b0000000000011011;
    assign weights1[52][80] = 16'b0000000000010001;
    assign weights1[52][81] = 16'b0000000000001000;
    assign weights1[52][82] = 16'b0000000000001000;
    assign weights1[52][83] = 16'b0000000000001001;
    assign weights1[52][84] = 16'b1111111111111101;
    assign weights1[52][85] = 16'b1111111111111101;
    assign weights1[52][86] = 16'b1111111111111100;
    assign weights1[52][87] = 16'b1111111111110101;
    assign weights1[52][88] = 16'b1111111111101111;
    assign weights1[52][89] = 16'b1111111111101100;
    assign weights1[52][90] = 16'b1111111111100001;
    assign weights1[52][91] = 16'b1111111111100101;
    assign weights1[52][92] = 16'b1111111111101110;
    assign weights1[52][93] = 16'b1111111111101000;
    assign weights1[52][94] = 16'b1111111111100010;
    assign weights1[52][95] = 16'b1111111111101010;
    assign weights1[52][96] = 16'b1111111111110000;
    assign weights1[52][97] = 16'b0000000000000101;
    assign weights1[52][98] = 16'b0000000000010100;
    assign weights1[52][99] = 16'b0000000000011011;
    assign weights1[52][100] = 16'b0000000000101011;
    assign weights1[52][101] = 16'b0000000000100101;
    assign weights1[52][102] = 16'b0000000000110101;
    assign weights1[52][103] = 16'b0000000000101000;
    assign weights1[52][104] = 16'b0000000000100101;
    assign weights1[52][105] = 16'b0000000000100111;
    assign weights1[52][106] = 16'b0000000000001110;
    assign weights1[52][107] = 16'b0000000000010111;
    assign weights1[52][108] = 16'b0000000000001000;
    assign weights1[52][109] = 16'b0000000000001001;
    assign weights1[52][110] = 16'b0000000000001100;
    assign weights1[52][111] = 16'b0000000000000110;
    assign weights1[52][112] = 16'b1111111111111011;
    assign weights1[52][113] = 16'b1111111111111101;
    assign weights1[52][114] = 16'b1111111111110000;
    assign weights1[52][115] = 16'b1111111111110001;
    assign weights1[52][116] = 16'b1111111111100011;
    assign weights1[52][117] = 16'b1111111111011101;
    assign weights1[52][118] = 16'b1111111111010001;
    assign weights1[52][119] = 16'b1111111111010000;
    assign weights1[52][120] = 16'b1111111111001110;
    assign weights1[52][121] = 16'b1111111110111011;
    assign weights1[52][122] = 16'b1111111110110011;
    assign weights1[52][123] = 16'b1111111110111101;
    assign weights1[52][124] = 16'b1111111111001001;
    assign weights1[52][125] = 16'b1111111111001111;
    assign weights1[52][126] = 16'b1111111111010110;
    assign weights1[52][127] = 16'b1111111111110001;
    assign weights1[52][128] = 16'b1111111111111001;
    assign weights1[52][129] = 16'b0000000000000111;
    assign weights1[52][130] = 16'b0000000000001111;
    assign weights1[52][131] = 16'b0000000000010100;
    assign weights1[52][132] = 16'b0000000000011010;
    assign weights1[52][133] = 16'b0000000000001011;
    assign weights1[52][134] = 16'b0000000000011011;
    assign weights1[52][135] = 16'b0000000000010110;
    assign weights1[52][136] = 16'b0000000000011010;
    assign weights1[52][137] = 16'b1111111111111001;
    assign weights1[52][138] = 16'b1111111111111111;
    assign weights1[52][139] = 16'b0000000000001000;
    assign weights1[52][140] = 16'b1111111111111100;
    assign weights1[52][141] = 16'b1111111111110001;
    assign weights1[52][142] = 16'b1111111111100001;
    assign weights1[52][143] = 16'b1111111111011000;
    assign weights1[52][144] = 16'b1111111111001100;
    assign weights1[52][145] = 16'b1111111111001100;
    assign weights1[52][146] = 16'b1111111110111000;
    assign weights1[52][147] = 16'b1111111110100111;
    assign weights1[52][148] = 16'b1111111110101010;
    assign weights1[52][149] = 16'b1111111110100100;
    assign weights1[52][150] = 16'b1111111110100101;
    assign weights1[52][151] = 16'b1111111110101000;
    assign weights1[52][152] = 16'b1111111110110000;
    assign weights1[52][153] = 16'b1111111110101110;
    assign weights1[52][154] = 16'b1111111110110111;
    assign weights1[52][155] = 16'b1111111110111011;
    assign weights1[52][156] = 16'b1111111111001111;
    assign weights1[52][157] = 16'b1111111111011010;
    assign weights1[52][158] = 16'b1111111111010111;
    assign weights1[52][159] = 16'b1111111111101010;
    assign weights1[52][160] = 16'b0000000000000011;
    assign weights1[52][161] = 16'b1111111111101100;
    assign weights1[52][162] = 16'b0000000000000011;
    assign weights1[52][163] = 16'b0000000000001111;
    assign weights1[52][164] = 16'b0000000000010010;
    assign weights1[52][165] = 16'b0000000000000111;
    assign weights1[52][166] = 16'b0000000000001100;
    assign weights1[52][167] = 16'b0000000000000111;
    assign weights1[52][168] = 16'b1111111111111000;
    assign weights1[52][169] = 16'b1111111111101110;
    assign weights1[52][170] = 16'b1111111111101001;
    assign weights1[52][171] = 16'b1111111111010110;
    assign weights1[52][172] = 16'b1111111111000101;
    assign weights1[52][173] = 16'b1111111110111110;
    assign weights1[52][174] = 16'b1111111110011011;
    assign weights1[52][175] = 16'b1111111110000110;
    assign weights1[52][176] = 16'b1111111110010010;
    assign weights1[52][177] = 16'b1111111110000011;
    assign weights1[52][178] = 16'b1111111110000110;
    assign weights1[52][179] = 16'b1111111110001010;
    assign weights1[52][180] = 16'b1111111110010111;
    assign weights1[52][181] = 16'b1111111110011011;
    assign weights1[52][182] = 16'b1111111110100000;
    assign weights1[52][183] = 16'b1111111110101000;
    assign weights1[52][184] = 16'b1111111110110011;
    assign weights1[52][185] = 16'b1111111110110111;
    assign weights1[52][186] = 16'b1111111111001101;
    assign weights1[52][187] = 16'b1111111111010111;
    assign weights1[52][188] = 16'b1111111111100010;
    assign weights1[52][189] = 16'b1111111111110110;
    assign weights1[52][190] = 16'b1111111111101000;
    assign weights1[52][191] = 16'b0000000000001000;
    assign weights1[52][192] = 16'b0000000000001011;
    assign weights1[52][193] = 16'b0000000000000001;
    assign weights1[52][194] = 16'b0000000000001000;
    assign weights1[52][195] = 16'b0000000000001010;
    assign weights1[52][196] = 16'b1111111111111000;
    assign weights1[52][197] = 16'b1111111111101111;
    assign weights1[52][198] = 16'b1111111111101101;
    assign weights1[52][199] = 16'b1111111111100001;
    assign weights1[52][200] = 16'b1111111111011100;
    assign weights1[52][201] = 16'b1111111111011111;
    assign weights1[52][202] = 16'b1111111111001001;
    assign weights1[52][203] = 16'b1111111110111110;
    assign weights1[52][204] = 16'b1111111111000100;
    assign weights1[52][205] = 16'b1111111110101111;
    assign weights1[52][206] = 16'b1111111110100110;
    assign weights1[52][207] = 16'b1111111110010011;
    assign weights1[52][208] = 16'b1111111110011000;
    assign weights1[52][209] = 16'b1111111110011100;
    assign weights1[52][210] = 16'b1111111110110110;
    assign weights1[52][211] = 16'b1111111110110111;
    assign weights1[52][212] = 16'b1111111110101010;
    assign weights1[52][213] = 16'b1111111110100111;
    assign weights1[52][214] = 16'b1111111111001100;
    assign weights1[52][215] = 16'b1111111111100000;
    assign weights1[52][216] = 16'b1111111111101100;
    assign weights1[52][217] = 16'b1111111111011000;
    assign weights1[52][218] = 16'b1111111111110100;
    assign weights1[52][219] = 16'b0000000000010010;
    assign weights1[52][220] = 16'b0000000000001100;
    assign weights1[52][221] = 16'b1111111111111111;
    assign weights1[52][222] = 16'b0000000000000110;
    assign weights1[52][223] = 16'b1111111111111110;
    assign weights1[52][224] = 16'b1111111111111011;
    assign weights1[52][225] = 16'b1111111111111000;
    assign weights1[52][226] = 16'b1111111111110110;
    assign weights1[52][227] = 16'b1111111111110111;
    assign weights1[52][228] = 16'b1111111111111111;
    assign weights1[52][229] = 16'b0000000000000001;
    assign weights1[52][230] = 16'b0000000000001011;
    assign weights1[52][231] = 16'b1111111111110000;
    assign weights1[52][232] = 16'b1111111111011101;
    assign weights1[52][233] = 16'b1111111111110010;
    assign weights1[52][234] = 16'b1111111110111111;
    assign weights1[52][235] = 16'b1111111111000111;
    assign weights1[52][236] = 16'b1111111110101101;
    assign weights1[52][237] = 16'b1111111111000011;
    assign weights1[52][238] = 16'b1111111111001110;
    assign weights1[52][239] = 16'b1111111111000001;
    assign weights1[52][240] = 16'b1111111111011011;
    assign weights1[52][241] = 16'b1111111111101001;
    assign weights1[52][242] = 16'b1111111111100111;
    assign weights1[52][243] = 16'b1111111111100000;
    assign weights1[52][244] = 16'b1111111111111101;
    assign weights1[52][245] = 16'b0000000000000011;
    assign weights1[52][246] = 16'b1111111111101110;
    assign weights1[52][247] = 16'b1111111111111100;
    assign weights1[52][248] = 16'b1111111111111100;
    assign weights1[52][249] = 16'b0000000000000111;
    assign weights1[52][250] = 16'b1111111111101001;
    assign weights1[52][251] = 16'b1111111111110110;
    assign weights1[52][252] = 16'b0000000000000110;
    assign weights1[52][253] = 16'b1111111111111011;
    assign weights1[52][254] = 16'b0000000000001010;
    assign weights1[52][255] = 16'b0000000000011001;
    assign weights1[52][256] = 16'b0000000000101011;
    assign weights1[52][257] = 16'b0000000000011100;
    assign weights1[52][258] = 16'b0000000000100000;
    assign weights1[52][259] = 16'b0000000000011000;
    assign weights1[52][260] = 16'b0000000000001000;
    assign weights1[52][261] = 16'b1111111111110111;
    assign weights1[52][262] = 16'b1111111111110111;
    assign weights1[52][263] = 16'b1111111111100101;
    assign weights1[52][264] = 16'b1111111111101111;
    assign weights1[52][265] = 16'b1111111111011111;
    assign weights1[52][266] = 16'b1111111111110011;
    assign weights1[52][267] = 16'b1111111111111010;
    assign weights1[52][268] = 16'b0000000000001111;
    assign weights1[52][269] = 16'b0000000000001001;
    assign weights1[52][270] = 16'b0000000000000010;
    assign weights1[52][271] = 16'b1111111111110000;
    assign weights1[52][272] = 16'b1111111111110101;
    assign weights1[52][273] = 16'b0000000000000100;
    assign weights1[52][274] = 16'b1111111111111011;
    assign weights1[52][275] = 16'b1111111111111000;
    assign weights1[52][276] = 16'b1111111111111100;
    assign weights1[52][277] = 16'b1111111111110000;
    assign weights1[52][278] = 16'b1111111111110110;
    assign weights1[52][279] = 16'b1111111111111110;
    assign weights1[52][280] = 16'b0000000000001111;
    assign weights1[52][281] = 16'b0000000000010001;
    assign weights1[52][282] = 16'b0000000000100110;
    assign weights1[52][283] = 16'b0000000000101100;
    assign weights1[52][284] = 16'b0000000000101000;
    assign weights1[52][285] = 16'b0000000000100101;
    assign weights1[52][286] = 16'b0000000000011110;
    assign weights1[52][287] = 16'b0000000000101110;
    assign weights1[52][288] = 16'b0000000000101010;
    assign weights1[52][289] = 16'b0000000000100100;
    assign weights1[52][290] = 16'b0000000000001111;
    assign weights1[52][291] = 16'b0000000000011001;
    assign weights1[52][292] = 16'b0000000000011011;
    assign weights1[52][293] = 16'b1111111111111000;
    assign weights1[52][294] = 16'b0000000000000000;
    assign weights1[52][295] = 16'b1111111111110010;
    assign weights1[52][296] = 16'b1111111111110110;
    assign weights1[52][297] = 16'b1111111111111100;
    assign weights1[52][298] = 16'b0000000000000001;
    assign weights1[52][299] = 16'b0000000000001100;
    assign weights1[52][300] = 16'b0000000000001100;
    assign weights1[52][301] = 16'b1111111111111110;
    assign weights1[52][302] = 16'b0000000000010101;
    assign weights1[52][303] = 16'b0000000000001011;
    assign weights1[52][304] = 16'b1111111111111011;
    assign weights1[52][305] = 16'b1111111111111100;
    assign weights1[52][306] = 16'b0000000000000101;
    assign weights1[52][307] = 16'b1111111111111000;
    assign weights1[52][308] = 16'b0000000000010101;
    assign weights1[52][309] = 16'b0000000000011110;
    assign weights1[52][310] = 16'b0000000000101010;
    assign weights1[52][311] = 16'b0000000000100000;
    assign weights1[52][312] = 16'b0000000000100001;
    assign weights1[52][313] = 16'b0000000000010111;
    assign weights1[52][314] = 16'b0000000000011101;
    assign weights1[52][315] = 16'b0000000000001011;
    assign weights1[52][316] = 16'b0000000000101010;
    assign weights1[52][317] = 16'b0000000000011100;
    assign weights1[52][318] = 16'b0000000000100100;
    assign weights1[52][319] = 16'b0000000000011101;
    assign weights1[52][320] = 16'b0000000000011101;
    assign weights1[52][321] = 16'b0000000000001111;
    assign weights1[52][322] = 16'b0000000000100011;
    assign weights1[52][323] = 16'b0000000000011001;
    assign weights1[52][324] = 16'b0000000000010011;
    assign weights1[52][325] = 16'b0000000000000010;
    assign weights1[52][326] = 16'b0000000000011010;
    assign weights1[52][327] = 16'b1111111111111101;
    assign weights1[52][328] = 16'b0000000000001001;
    assign weights1[52][329] = 16'b0000000000010000;
    assign weights1[52][330] = 16'b0000000000000001;
    assign weights1[52][331] = 16'b0000000000000001;
    assign weights1[52][332] = 16'b1111111111100101;
    assign weights1[52][333] = 16'b0000000000000111;
    assign weights1[52][334] = 16'b0000000000001010;
    assign weights1[52][335] = 16'b1111111111101111;
    assign weights1[52][336] = 16'b0000000000011010;
    assign weights1[52][337] = 16'b0000000000010111;
    assign weights1[52][338] = 16'b0000000000011100;
    assign weights1[52][339] = 16'b0000000000001111;
    assign weights1[52][340] = 16'b1111111111110011;
    assign weights1[52][341] = 16'b0000000000000110;
    assign weights1[52][342] = 16'b0000000000001001;
    assign weights1[52][343] = 16'b0000000000011110;
    assign weights1[52][344] = 16'b0000000000110011;
    assign weights1[52][345] = 16'b0000000000010010;
    assign weights1[52][346] = 16'b0000000000010100;
    assign weights1[52][347] = 16'b0000000000101101;
    assign weights1[52][348] = 16'b0000000000100110;
    assign weights1[52][349] = 16'b0000000000110011;
    assign weights1[52][350] = 16'b0000000000101111;
    assign weights1[52][351] = 16'b0000000000011011;
    assign weights1[52][352] = 16'b0000000000101000;
    assign weights1[52][353] = 16'b0000000000010110;
    assign weights1[52][354] = 16'b0000000000010111;
    assign weights1[52][355] = 16'b0000000000011000;
    assign weights1[52][356] = 16'b0000000000010001;
    assign weights1[52][357] = 16'b0000000000000011;
    assign weights1[52][358] = 16'b1111111111111100;
    assign weights1[52][359] = 16'b1111111111111101;
    assign weights1[52][360] = 16'b0000000000000110;
    assign weights1[52][361] = 16'b0000000000001000;
    assign weights1[52][362] = 16'b1111111111111101;
    assign weights1[52][363] = 16'b1111111111111100;
    assign weights1[52][364] = 16'b0000000000011001;
    assign weights1[52][365] = 16'b0000000000010111;
    assign weights1[52][366] = 16'b0000000000001000;
    assign weights1[52][367] = 16'b1111111111111000;
    assign weights1[52][368] = 16'b1111111111111110;
    assign weights1[52][369] = 16'b0000000000010100;
    assign weights1[52][370] = 16'b1111111111110111;
    assign weights1[52][371] = 16'b1111111111110110;
    assign weights1[52][372] = 16'b0000000000001010;
    assign weights1[52][373] = 16'b0000000000011010;
    assign weights1[52][374] = 16'b0000000000011111;
    assign weights1[52][375] = 16'b0000000000011111;
    assign weights1[52][376] = 16'b0000000000101110;
    assign weights1[52][377] = 16'b0000000000011111;
    assign weights1[52][378] = 16'b0000000000011000;
    assign weights1[52][379] = 16'b0000000000101100;
    assign weights1[52][380] = 16'b0000000000011001;
    assign weights1[52][381] = 16'b0000000000100100;
    assign weights1[52][382] = 16'b0000000000110000;
    assign weights1[52][383] = 16'b0000000000001010;
    assign weights1[52][384] = 16'b0000000000010000;
    assign weights1[52][385] = 16'b0000000000010110;
    assign weights1[52][386] = 16'b0000000000000101;
    assign weights1[52][387] = 16'b0000000000000011;
    assign weights1[52][388] = 16'b0000000000000100;
    assign weights1[52][389] = 16'b0000000000001100;
    assign weights1[52][390] = 16'b0000000000010000;
    assign weights1[52][391] = 16'b1111111111110010;
    assign weights1[52][392] = 16'b0000000000010011;
    assign weights1[52][393] = 16'b0000000000001100;
    assign weights1[52][394] = 16'b0000000000000001;
    assign weights1[52][395] = 16'b1111111111111111;
    assign weights1[52][396] = 16'b0000000000000001;
    assign weights1[52][397] = 16'b1111111111011111;
    assign weights1[52][398] = 16'b1111111111110001;
    assign weights1[52][399] = 16'b1111111111110010;
    assign weights1[52][400] = 16'b0000000000000011;
    assign weights1[52][401] = 16'b1111111111111001;
    assign weights1[52][402] = 16'b0000000000000000;
    assign weights1[52][403] = 16'b1111111111111111;
    assign weights1[52][404] = 16'b0000000000001011;
    assign weights1[52][405] = 16'b0000000000000010;
    assign weights1[52][406] = 16'b0000000000000111;
    assign weights1[52][407] = 16'b0000000000001100;
    assign weights1[52][408] = 16'b0000000000010000;
    assign weights1[52][409] = 16'b0000000000000010;
    assign weights1[52][410] = 16'b0000000000001011;
    assign weights1[52][411] = 16'b0000000000011011;
    assign weights1[52][412] = 16'b0000000000001110;
    assign weights1[52][413] = 16'b1111111111111000;
    assign weights1[52][414] = 16'b0000000000010011;
    assign weights1[52][415] = 16'b0000000000011001;
    assign weights1[52][416] = 16'b1111111111111100;
    assign weights1[52][417] = 16'b0000000000000111;
    assign weights1[52][418] = 16'b0000000000001000;
    assign weights1[52][419] = 16'b1111111111111111;
    assign weights1[52][420] = 16'b0000000000010110;
    assign weights1[52][421] = 16'b0000000000010011;
    assign weights1[52][422] = 16'b0000000000000000;
    assign weights1[52][423] = 16'b1111111111110011;
    assign weights1[52][424] = 16'b1111111111100011;
    assign weights1[52][425] = 16'b1111111111110000;
    assign weights1[52][426] = 16'b0000000000000101;
    assign weights1[52][427] = 16'b1111111111111000;
    assign weights1[52][428] = 16'b1111111111110111;
    assign weights1[52][429] = 16'b1111111111111110;
    assign weights1[52][430] = 16'b1111111111111110;
    assign weights1[52][431] = 16'b1111111111110000;
    assign weights1[52][432] = 16'b1111111111100000;
    assign weights1[52][433] = 16'b1111111111100111;
    assign weights1[52][434] = 16'b1111111111100111;
    assign weights1[52][435] = 16'b1111111111011001;
    assign weights1[52][436] = 16'b1111111111011011;
    assign weights1[52][437] = 16'b1111111111110011;
    assign weights1[52][438] = 16'b1111111111111000;
    assign weights1[52][439] = 16'b1111111111110110;
    assign weights1[52][440] = 16'b0000000000000110;
    assign weights1[52][441] = 16'b1111111111110111;
    assign weights1[52][442] = 16'b1111111111111111;
    assign weights1[52][443] = 16'b1111111111110111;
    assign weights1[52][444] = 16'b0000000000001011;
    assign weights1[52][445] = 16'b0000000000001010;
    assign weights1[52][446] = 16'b1111111111111110;
    assign weights1[52][447] = 16'b0000000000010001;
    assign weights1[52][448] = 16'b0000000000001010;
    assign weights1[52][449] = 16'b0000000000000111;
    assign weights1[52][450] = 16'b0000000000000100;
    assign weights1[52][451] = 16'b0000000000000001;
    assign weights1[52][452] = 16'b1111111111111110;
    assign weights1[52][453] = 16'b1111111111111010;
    assign weights1[52][454] = 16'b1111111111110100;
    assign weights1[52][455] = 16'b1111111111111111;
    assign weights1[52][456] = 16'b0000000000000111;
    assign weights1[52][457] = 16'b1111111111101100;
    assign weights1[52][458] = 16'b1111111111011110;
    assign weights1[52][459] = 16'b1111111111110111;
    assign weights1[52][460] = 16'b1111111111011001;
    assign weights1[52][461] = 16'b1111111111010111;
    assign weights1[52][462] = 16'b1111111111010011;
    assign weights1[52][463] = 16'b1111111111010000;
    assign weights1[52][464] = 16'b1111111111011010;
    assign weights1[52][465] = 16'b1111111111011110;
    assign weights1[52][466] = 16'b1111111111101000;
    assign weights1[52][467] = 16'b1111111111110111;
    assign weights1[52][468] = 16'b1111111111110100;
    assign weights1[52][469] = 16'b1111111111110010;
    assign weights1[52][470] = 16'b1111111111111001;
    assign weights1[52][471] = 16'b1111111111110000;
    assign weights1[52][472] = 16'b1111111111111001;
    assign weights1[52][473] = 16'b0000000000000001;
    assign weights1[52][474] = 16'b0000000000000011;
    assign weights1[52][475] = 16'b0000000000011000;
    assign weights1[52][476] = 16'b0000000000000100;
    assign weights1[52][477] = 16'b0000000000000110;
    assign weights1[52][478] = 16'b1111111111110100;
    assign weights1[52][479] = 16'b1111111111111010;
    assign weights1[52][480] = 16'b0000000000001101;
    assign weights1[52][481] = 16'b1111111111111001;
    assign weights1[52][482] = 16'b0000000000011001;
    assign weights1[52][483] = 16'b1111111111111010;
    assign weights1[52][484] = 16'b1111111111101010;
    assign weights1[52][485] = 16'b1111111111100100;
    assign weights1[52][486] = 16'b1111111111011110;
    assign weights1[52][487] = 16'b1111111111011100;
    assign weights1[52][488] = 16'b1111111111010101;
    assign weights1[52][489] = 16'b1111111111010101;
    assign weights1[52][490] = 16'b1111111111100000;
    assign weights1[52][491] = 16'b1111111111010111;
    assign weights1[52][492] = 16'b1111111111011000;
    assign weights1[52][493] = 16'b1111111111010111;
    assign weights1[52][494] = 16'b1111111111100000;
    assign weights1[52][495] = 16'b1111111111001011;
    assign weights1[52][496] = 16'b1111111111101010;
    assign weights1[52][497] = 16'b1111111111110010;
    assign weights1[52][498] = 16'b0000000000001000;
    assign weights1[52][499] = 16'b1111111111101101;
    assign weights1[52][500] = 16'b0000000000010010;
    assign weights1[52][501] = 16'b0000000000000001;
    assign weights1[52][502] = 16'b0000000000000010;
    assign weights1[52][503] = 16'b0000000000010111;
    assign weights1[52][504] = 16'b1111111111111110;
    assign weights1[52][505] = 16'b1111111111111001;
    assign weights1[52][506] = 16'b1111111111101110;
    assign weights1[52][507] = 16'b1111111111110011;
    assign weights1[52][508] = 16'b1111111111111010;
    assign weights1[52][509] = 16'b1111111111110101;
    assign weights1[52][510] = 16'b0000000000000000;
    assign weights1[52][511] = 16'b1111111111100001;
    assign weights1[52][512] = 16'b1111111111100110;
    assign weights1[52][513] = 16'b1111111111010111;
    assign weights1[52][514] = 16'b1111111111010011;
    assign weights1[52][515] = 16'b1111111111010111;
    assign weights1[52][516] = 16'b1111111111011011;
    assign weights1[52][517] = 16'b1111111111011011;
    assign weights1[52][518] = 16'b1111111111101011;
    assign weights1[52][519] = 16'b1111111111010011;
    assign weights1[52][520] = 16'b1111111111100010;
    assign weights1[52][521] = 16'b1111111111101011;
    assign weights1[52][522] = 16'b1111111111100100;
    assign weights1[52][523] = 16'b1111111111011100;
    assign weights1[52][524] = 16'b1111111111110010;
    assign weights1[52][525] = 16'b0000000000001000;
    assign weights1[52][526] = 16'b1111111111101101;
    assign weights1[52][527] = 16'b0000000000001000;
    assign weights1[52][528] = 16'b0000000000010010;
    assign weights1[52][529] = 16'b0000000000000100;
    assign weights1[52][530] = 16'b0000000000011001;
    assign weights1[52][531] = 16'b0000000000010000;
    assign weights1[52][532] = 16'b0000000000000001;
    assign weights1[52][533] = 16'b1111111111110111;
    assign weights1[52][534] = 16'b1111111111111010;
    assign weights1[52][535] = 16'b1111111111111000;
    assign weights1[52][536] = 16'b1111111111101010;
    assign weights1[52][537] = 16'b1111111111101111;
    assign weights1[52][538] = 16'b1111111111101000;
    assign weights1[52][539] = 16'b1111111111011000;
    assign weights1[52][540] = 16'b1111111111100000;
    assign weights1[52][541] = 16'b1111111111011101;
    assign weights1[52][542] = 16'b1111111111001101;
    assign weights1[52][543] = 16'b1111111111001101;
    assign weights1[52][544] = 16'b1111111111011100;
    assign weights1[52][545] = 16'b1111111111100101;
    assign weights1[52][546] = 16'b1111111111010111;
    assign weights1[52][547] = 16'b1111111111101000;
    assign weights1[52][548] = 16'b1111111111101111;
    assign weights1[52][549] = 16'b0000000000000000;
    assign weights1[52][550] = 16'b1111111111011101;
    assign weights1[52][551] = 16'b1111111111111100;
    assign weights1[52][552] = 16'b1111111111111111;
    assign weights1[52][553] = 16'b1111111111111111;
    assign weights1[52][554] = 16'b0000000000001000;
    assign weights1[52][555] = 16'b0000000000001111;
    assign weights1[52][556] = 16'b0000000000001000;
    assign weights1[52][557] = 16'b0000000000000110;
    assign weights1[52][558] = 16'b0000000000010101;
    assign weights1[52][559] = 16'b0000000000011100;
    assign weights1[52][560] = 16'b0000000000000110;
    assign weights1[52][561] = 16'b0000000000001001;
    assign weights1[52][562] = 16'b1111111111111100;
    assign weights1[52][563] = 16'b1111111111110100;
    assign weights1[52][564] = 16'b1111111111100011;
    assign weights1[52][565] = 16'b1111111111101100;
    assign weights1[52][566] = 16'b1111111111110011;
    assign weights1[52][567] = 16'b1111111111110010;
    assign weights1[52][568] = 16'b1111111111011111;
    assign weights1[52][569] = 16'b1111111111101010;
    assign weights1[52][570] = 16'b1111111111100111;
    assign weights1[52][571] = 16'b1111111111100011;
    assign weights1[52][572] = 16'b1111111111100011;
    assign weights1[52][573] = 16'b1111111111011110;
    assign weights1[52][574] = 16'b1111111111101001;
    assign weights1[52][575] = 16'b0000000000000000;
    assign weights1[52][576] = 16'b1111111111101010;
    assign weights1[52][577] = 16'b1111111111101010;
    assign weights1[52][578] = 16'b1111111111111100;
    assign weights1[52][579] = 16'b0000000000000011;
    assign weights1[52][580] = 16'b0000000000010011;
    assign weights1[52][581] = 16'b0000000000000000;
    assign weights1[52][582] = 16'b0000000000010010;
    assign weights1[52][583] = 16'b0000000000001010;
    assign weights1[52][584] = 16'b0000000000000111;
    assign weights1[52][585] = 16'b0000000000001000;
    assign weights1[52][586] = 16'b0000000000010101;
    assign weights1[52][587] = 16'b0000000000010000;
    assign weights1[52][588] = 16'b0000000000000111;
    assign weights1[52][589] = 16'b1111111111111110;
    assign weights1[52][590] = 16'b1111111111111001;
    assign weights1[52][591] = 16'b1111111111111000;
    assign weights1[52][592] = 16'b1111111111111100;
    assign weights1[52][593] = 16'b0000000000001011;
    assign weights1[52][594] = 16'b1111111111111010;
    assign weights1[52][595] = 16'b1111111111110011;
    assign weights1[52][596] = 16'b1111111111110111;
    assign weights1[52][597] = 16'b1111111111101110;
    assign weights1[52][598] = 16'b1111111111011110;
    assign weights1[52][599] = 16'b1111111111100110;
    assign weights1[52][600] = 16'b1111111111100011;
    assign weights1[52][601] = 16'b1111111111101010;
    assign weights1[52][602] = 16'b1111111111110110;
    assign weights1[52][603] = 16'b1111111111101000;
    assign weights1[52][604] = 16'b1111111111110010;
    assign weights1[52][605] = 16'b0000000000000101;
    assign weights1[52][606] = 16'b1111111111111100;
    assign weights1[52][607] = 16'b1111111111111111;
    assign weights1[52][608] = 16'b0000000000100010;
    assign weights1[52][609] = 16'b0000000000001000;
    assign weights1[52][610] = 16'b0000000000001101;
    assign weights1[52][611] = 16'b0000000000010110;
    assign weights1[52][612] = 16'b1111111111111100;
    assign weights1[52][613] = 16'b0000000000000111;
    assign weights1[52][614] = 16'b0000000000001101;
    assign weights1[52][615] = 16'b0000000000010010;
    assign weights1[52][616] = 16'b0000000000001000;
    assign weights1[52][617] = 16'b0000000000000000;
    assign weights1[52][618] = 16'b0000000000001010;
    assign weights1[52][619] = 16'b0000000000000011;
    assign weights1[52][620] = 16'b0000000000001010;
    assign weights1[52][621] = 16'b0000000000001111;
    assign weights1[52][622] = 16'b1111111111111010;
    assign weights1[52][623] = 16'b0000000000000110;
    assign weights1[52][624] = 16'b0000000000001011;
    assign weights1[52][625] = 16'b0000000000010100;
    assign weights1[52][626] = 16'b1111111111111001;
    assign weights1[52][627] = 16'b0000000000010101;
    assign weights1[52][628] = 16'b0000000000001010;
    assign weights1[52][629] = 16'b0000000000001001;
    assign weights1[52][630] = 16'b0000000000000010;
    assign weights1[52][631] = 16'b0000000000000111;
    assign weights1[52][632] = 16'b0000000000000101;
    assign weights1[52][633] = 16'b0000000000000000;
    assign weights1[52][634] = 16'b0000000000001000;
    assign weights1[52][635] = 16'b0000000000000101;
    assign weights1[52][636] = 16'b1111111111110111;
    assign weights1[52][637] = 16'b0000000000000011;
    assign weights1[52][638] = 16'b0000000000010000;
    assign weights1[52][639] = 16'b0000000000001011;
    assign weights1[52][640] = 16'b0000000000001011;
    assign weights1[52][641] = 16'b0000000000010101;
    assign weights1[52][642] = 16'b0000000000000100;
    assign weights1[52][643] = 16'b0000000000001001;
    assign weights1[52][644] = 16'b0000000000000101;
    assign weights1[52][645] = 16'b0000000000000101;
    assign weights1[52][646] = 16'b0000000000010000;
    assign weights1[52][647] = 16'b0000000000001000;
    assign weights1[52][648] = 16'b0000000000001001;
    assign weights1[52][649] = 16'b0000000000010100;
    assign weights1[52][650] = 16'b0000000000000101;
    assign weights1[52][651] = 16'b0000000000000111;
    assign weights1[52][652] = 16'b0000000000011000;
    assign weights1[52][653] = 16'b0000000000010011;
    assign weights1[52][654] = 16'b0000000000011011;
    assign weights1[52][655] = 16'b0000000000011100;
    assign weights1[52][656] = 16'b0000000000001010;
    assign weights1[52][657] = 16'b0000000000010111;
    assign weights1[52][658] = 16'b0000000000010011;
    assign weights1[52][659] = 16'b0000000000010011;
    assign weights1[52][660] = 16'b0000000000010001;
    assign weights1[52][661] = 16'b0000000000010001;
    assign weights1[52][662] = 16'b0000000000011101;
    assign weights1[52][663] = 16'b0000000000001111;
    assign weights1[52][664] = 16'b1111111111111011;
    assign weights1[52][665] = 16'b0000000000000011;
    assign weights1[52][666] = 16'b1111111111110010;
    assign weights1[52][667] = 16'b0000000000000001;
    assign weights1[52][668] = 16'b0000000000000000;
    assign weights1[52][669] = 16'b1111111111111100;
    assign weights1[52][670] = 16'b1111111111111110;
    assign weights1[52][671] = 16'b1111111111111110;
    assign weights1[52][672] = 16'b0000000000001010;
    assign weights1[52][673] = 16'b0000000000001010;
    assign weights1[52][674] = 16'b0000000000001011;
    assign weights1[52][675] = 16'b0000000000001110;
    assign weights1[52][676] = 16'b0000000000010101;
    assign weights1[52][677] = 16'b0000000000001111;
    assign weights1[52][678] = 16'b0000000000101100;
    assign weights1[52][679] = 16'b0000000000010110;
    assign weights1[52][680] = 16'b0000000000101101;
    assign weights1[52][681] = 16'b0000000000011011;
    assign weights1[52][682] = 16'b0000000000100111;
    assign weights1[52][683] = 16'b0000000000011110;
    assign weights1[52][684] = 16'b0000000000100111;
    assign weights1[52][685] = 16'b0000000000011111;
    assign weights1[52][686] = 16'b0000000000010001;
    assign weights1[52][687] = 16'b0000000000001111;
    assign weights1[52][688] = 16'b0000000000001100;
    assign weights1[52][689] = 16'b0000000000001010;
    assign weights1[52][690] = 16'b0000000000001000;
    assign weights1[52][691] = 16'b0000000000000011;
    assign weights1[52][692] = 16'b1111111111111010;
    assign weights1[52][693] = 16'b1111111111111010;
    assign weights1[52][694] = 16'b1111111111101101;
    assign weights1[52][695] = 16'b1111111111011010;
    assign weights1[52][696] = 16'b1111111111110111;
    assign weights1[52][697] = 16'b1111111111111010;
    assign weights1[52][698] = 16'b1111111111111011;
    assign weights1[52][699] = 16'b1111111111111101;
    assign weights1[52][700] = 16'b0000000000001001;
    assign weights1[52][701] = 16'b0000000000010000;
    assign weights1[52][702] = 16'b0000000000001010;
    assign weights1[52][703] = 16'b0000000000000101;
    assign weights1[52][704] = 16'b0000000000010100;
    assign weights1[52][705] = 16'b0000000000010110;
    assign weights1[52][706] = 16'b0000000000100110;
    assign weights1[52][707] = 16'b0000000000000110;
    assign weights1[52][708] = 16'b0000000000010101;
    assign weights1[52][709] = 16'b0000000000001110;
    assign weights1[52][710] = 16'b0000000000011010;
    assign weights1[52][711] = 16'b0000000000001011;
    assign weights1[52][712] = 16'b0000000000000111;
    assign weights1[52][713] = 16'b0000000000010010;
    assign weights1[52][714] = 16'b0000000000011100;
    assign weights1[52][715] = 16'b0000000000000000;
    assign weights1[52][716] = 16'b0000000000010101;
    assign weights1[52][717] = 16'b1111111111111100;
    assign weights1[52][718] = 16'b0000000000000100;
    assign weights1[52][719] = 16'b0000000000010110;
    assign weights1[52][720] = 16'b1111111111111001;
    assign weights1[52][721] = 16'b0000000000001101;
    assign weights1[52][722] = 16'b1111111111111010;
    assign weights1[52][723] = 16'b1111111111111100;
    assign weights1[52][724] = 16'b1111111111111101;
    assign weights1[52][725] = 16'b1111111111101000;
    assign weights1[52][726] = 16'b1111111111110110;
    assign weights1[52][727] = 16'b1111111111111100;
    assign weights1[52][728] = 16'b0000000000001001;
    assign weights1[52][729] = 16'b0000000000001110;
    assign weights1[52][730] = 16'b0000000000001001;
    assign weights1[52][731] = 16'b0000000000001010;
    assign weights1[52][732] = 16'b0000000000010100;
    assign weights1[52][733] = 16'b0000000000010010;
    assign weights1[52][734] = 16'b0000000000011111;
    assign weights1[52][735] = 16'b0000000000000110;
    assign weights1[52][736] = 16'b0000000000000110;
    assign weights1[52][737] = 16'b0000000000001011;
    assign weights1[52][738] = 16'b1111111111110100;
    assign weights1[52][739] = 16'b0000000000001000;
    assign weights1[52][740] = 16'b0000000000001000;
    assign weights1[52][741] = 16'b1111111111111011;
    assign weights1[52][742] = 16'b1111111111111010;
    assign weights1[52][743] = 16'b0000000000001010;
    assign weights1[52][744] = 16'b0000000000000000;
    assign weights1[52][745] = 16'b1111111111111101;
    assign weights1[52][746] = 16'b0000000000001001;
    assign weights1[52][747] = 16'b0000000000011010;
    assign weights1[52][748] = 16'b1111111111111010;
    assign weights1[52][749] = 16'b0000000000000100;
    assign weights1[52][750] = 16'b0000000000001010;
    assign weights1[52][751] = 16'b0000000000001101;
    assign weights1[52][752] = 16'b1111111111111011;
    assign weights1[52][753] = 16'b1111111111110001;
    assign weights1[52][754] = 16'b1111111111110111;
    assign weights1[52][755] = 16'b1111111111111101;
    assign weights1[52][756] = 16'b0000000000000010;
    assign weights1[52][757] = 16'b0000000000001100;
    assign weights1[52][758] = 16'b1111111111111111;
    assign weights1[52][759] = 16'b1111111111111100;
    assign weights1[52][760] = 16'b0000000000000010;
    assign weights1[52][761] = 16'b0000000000010101;
    assign weights1[52][762] = 16'b0000000000011010;
    assign weights1[52][763] = 16'b1111111111111111;
    assign weights1[52][764] = 16'b0000000000010000;
    assign weights1[52][765] = 16'b0000000000000000;
    assign weights1[52][766] = 16'b0000000000001110;
    assign weights1[52][767] = 16'b0000000000001100;
    assign weights1[52][768] = 16'b1111111111111110;
    assign weights1[52][769] = 16'b0000000000001010;
    assign weights1[52][770] = 16'b0000000000001101;
    assign weights1[52][771] = 16'b0000000000000010;
    assign weights1[52][772] = 16'b0000000000001111;
    assign weights1[52][773] = 16'b0000000000010001;
    assign weights1[52][774] = 16'b1111111111111000;
    assign weights1[52][775] = 16'b1111111111111001;
    assign weights1[52][776] = 16'b0000000000000101;
    assign weights1[52][777] = 16'b0000000000000110;
    assign weights1[52][778] = 16'b0000000000000101;
    assign weights1[52][779] = 16'b1111111111111111;
    assign weights1[52][780] = 16'b1111111111111101;
    assign weights1[52][781] = 16'b1111111111111010;
    assign weights1[52][782] = 16'b1111111111111101;
    assign weights1[52][783] = 16'b0000000000000000;
    assign weights1[53][0] = 16'b0000000000000001;
    assign weights1[53][1] = 16'b0000000000000001;
    assign weights1[53][2] = 16'b1111111111111100;
    assign weights1[53][3] = 16'b1111111111110100;
    assign weights1[53][4] = 16'b1111111111110011;
    assign weights1[53][5] = 16'b1111111111101001;
    assign weights1[53][6] = 16'b1111111111100101;
    assign weights1[53][7] = 16'b1111111111011010;
    assign weights1[53][8] = 16'b1111111111010000;
    assign weights1[53][9] = 16'b1111111111010001;
    assign weights1[53][10] = 16'b1111111111010000;
    assign weights1[53][11] = 16'b1111111111010110;
    assign weights1[53][12] = 16'b1111111111001110;
    assign weights1[53][13] = 16'b1111111111010000;
    assign weights1[53][14] = 16'b1111111111100010;
    assign weights1[53][15] = 16'b1111111111010111;
    assign weights1[53][16] = 16'b1111111111010100;
    assign weights1[53][17] = 16'b1111111111011110;
    assign weights1[53][18] = 16'b1111111111101100;
    assign weights1[53][19] = 16'b1111111111100010;
    assign weights1[53][20] = 16'b1111111111101000;
    assign weights1[53][21] = 16'b1111111111110011;
    assign weights1[53][22] = 16'b1111111111111001;
    assign weights1[53][23] = 16'b1111111111111000;
    assign weights1[53][24] = 16'b1111111111111011;
    assign weights1[53][25] = 16'b1111111111111011;
    assign weights1[53][26] = 16'b1111111111111101;
    assign weights1[53][27] = 16'b1111111111111101;
    assign weights1[53][28] = 16'b0000000000000000;
    assign weights1[53][29] = 16'b1111111111111111;
    assign weights1[53][30] = 16'b1111111111111010;
    assign weights1[53][31] = 16'b1111111111110000;
    assign weights1[53][32] = 16'b1111111111100110;
    assign weights1[53][33] = 16'b1111111111011111;
    assign weights1[53][34] = 16'b1111111111010110;
    assign weights1[53][35] = 16'b1111111111001101;
    assign weights1[53][36] = 16'b1111111111001010;
    assign weights1[53][37] = 16'b1111111111000011;
    assign weights1[53][38] = 16'b1111111110111111;
    assign weights1[53][39] = 16'b1111111110111101;
    assign weights1[53][40] = 16'b1111111110111101;
    assign weights1[53][41] = 16'b1111111110111101;
    assign weights1[53][42] = 16'b1111111111001110;
    assign weights1[53][43] = 16'b1111111111010011;
    assign weights1[53][44] = 16'b1111111111010011;
    assign weights1[53][45] = 16'b1111111111001111;
    assign weights1[53][46] = 16'b1111111111100001;
    assign weights1[53][47] = 16'b1111111111100100;
    assign weights1[53][48] = 16'b1111111111100101;
    assign weights1[53][49] = 16'b1111111111101010;
    assign weights1[53][50] = 16'b1111111111101001;
    assign weights1[53][51] = 16'b1111111111100111;
    assign weights1[53][52] = 16'b1111111111101111;
    assign weights1[53][53] = 16'b1111111111111100;
    assign weights1[53][54] = 16'b1111111111111111;
    assign weights1[53][55] = 16'b1111111111111011;
    assign weights1[53][56] = 16'b1111111111111100;
    assign weights1[53][57] = 16'b1111111111111110;
    assign weights1[53][58] = 16'b1111111111111000;
    assign weights1[53][59] = 16'b1111111111101010;
    assign weights1[53][60] = 16'b1111111111010101;
    assign weights1[53][61] = 16'b1111111111010010;
    assign weights1[53][62] = 16'b1111111110111110;
    assign weights1[53][63] = 16'b1111111110111000;
    assign weights1[53][64] = 16'b1111111111000011;
    assign weights1[53][65] = 16'b1111111110110100;
    assign weights1[53][66] = 16'b1111111110101101;
    assign weights1[53][67] = 16'b1111111110110110;
    assign weights1[53][68] = 16'b1111111110111101;
    assign weights1[53][69] = 16'b1111111111001001;
    assign weights1[53][70] = 16'b1111111111001100;
    assign weights1[53][71] = 16'b1111111111001011;
    assign weights1[53][72] = 16'b1111111110111101;
    assign weights1[53][73] = 16'b1111111110111100;
    assign weights1[53][74] = 16'b1111111111010111;
    assign weights1[53][75] = 16'b1111111111011011;
    assign weights1[53][76] = 16'b1111111111011101;
    assign weights1[53][77] = 16'b1111111111100000;
    assign weights1[53][78] = 16'b1111111111100001;
    assign weights1[53][79] = 16'b1111111111101000;
    assign weights1[53][80] = 16'b1111111111011101;
    assign weights1[53][81] = 16'b1111111111101110;
    assign weights1[53][82] = 16'b1111111111110010;
    assign weights1[53][83] = 16'b1111111111111000;
    assign weights1[53][84] = 16'b1111111111111100;
    assign weights1[53][85] = 16'b1111111111111010;
    assign weights1[53][86] = 16'b1111111111110010;
    assign weights1[53][87] = 16'b1111111111100011;
    assign weights1[53][88] = 16'b1111111111010100;
    assign weights1[53][89] = 16'b1111111111001000;
    assign weights1[53][90] = 16'b1111111111000010;
    assign weights1[53][91] = 16'b1111111110110110;
    assign weights1[53][92] = 16'b1111111110111010;
    assign weights1[53][93] = 16'b1111111110111010;
    assign weights1[53][94] = 16'b1111111111000100;
    assign weights1[53][95] = 16'b1111111111001101;
    assign weights1[53][96] = 16'b1111111111010000;
    assign weights1[53][97] = 16'b1111111110110111;
    assign weights1[53][98] = 16'b1111111111011000;
    assign weights1[53][99] = 16'b1111111111001011;
    assign weights1[53][100] = 16'b1111111111001001;
    assign weights1[53][101] = 16'b1111111111011100;
    assign weights1[53][102] = 16'b1111111111010100;
    assign weights1[53][103] = 16'b1111111110111111;
    assign weights1[53][104] = 16'b1111111111001111;
    assign weights1[53][105] = 16'b1111111111010000;
    assign weights1[53][106] = 16'b1111111111001101;
    assign weights1[53][107] = 16'b1111111111011010;
    assign weights1[53][108] = 16'b1111111111011101;
    assign weights1[53][109] = 16'b1111111111100111;
    assign weights1[53][110] = 16'b1111111111110000;
    assign weights1[53][111] = 16'b1111111111110100;
    assign weights1[53][112] = 16'b1111111111111110;
    assign weights1[53][113] = 16'b1111111111110111;
    assign weights1[53][114] = 16'b1111111111110011;
    assign weights1[53][115] = 16'b1111111111101001;
    assign weights1[53][116] = 16'b1111111111010101;
    assign weights1[53][117] = 16'b1111111111000101;
    assign weights1[53][118] = 16'b1111111111011011;
    assign weights1[53][119] = 16'b1111111111000111;
    assign weights1[53][120] = 16'b1111111111010111;
    assign weights1[53][121] = 16'b1111111111001011;
    assign weights1[53][122] = 16'b1111111110111010;
    assign weights1[53][123] = 16'b1111111111010001;
    assign weights1[53][124] = 16'b1111111111010111;
    assign weights1[53][125] = 16'b1111111111011000;
    assign weights1[53][126] = 16'b1111111111001101;
    assign weights1[53][127] = 16'b1111111111100101;
    assign weights1[53][128] = 16'b1111111111111001;
    assign weights1[53][129] = 16'b1111111111011001;
    assign weights1[53][130] = 16'b1111111111010011;
    assign weights1[53][131] = 16'b1111111111010000;
    assign weights1[53][132] = 16'b1111111111010100;
    assign weights1[53][133] = 16'b1111111111100111;
    assign weights1[53][134] = 16'b1111111111100000;
    assign weights1[53][135] = 16'b1111111111011110;
    assign weights1[53][136] = 16'b1111111111101110;
    assign weights1[53][137] = 16'b1111111111101000;
    assign weights1[53][138] = 16'b1111111111111011;
    assign weights1[53][139] = 16'b1111111111111110;
    assign weights1[53][140] = 16'b1111111111111111;
    assign weights1[53][141] = 16'b1111111111111001;
    assign weights1[53][142] = 16'b1111111111110110;
    assign weights1[53][143] = 16'b1111111111100101;
    assign weights1[53][144] = 16'b1111111111011011;
    assign weights1[53][145] = 16'b1111111111010100;
    assign weights1[53][146] = 16'b1111111111011111;
    assign weights1[53][147] = 16'b1111111111010001;
    assign weights1[53][148] = 16'b1111111111111101;
    assign weights1[53][149] = 16'b1111111111111100;
    assign weights1[53][150] = 16'b1111111111100001;
    assign weights1[53][151] = 16'b1111111111111100;
    assign weights1[53][152] = 16'b0000000000000001;
    assign weights1[53][153] = 16'b1111111111001100;
    assign weights1[53][154] = 16'b1111111111010101;
    assign weights1[53][155] = 16'b1111111111001110;
    assign weights1[53][156] = 16'b1111111111010101;
    assign weights1[53][157] = 16'b1111111111100010;
    assign weights1[53][158] = 16'b1111111111001000;
    assign weights1[53][159] = 16'b1111111111000110;
    assign weights1[53][160] = 16'b1111111111000101;
    assign weights1[53][161] = 16'b1111111111001010;
    assign weights1[53][162] = 16'b1111111111101000;
    assign weights1[53][163] = 16'b1111111111110101;
    assign weights1[53][164] = 16'b1111111111111001;
    assign weights1[53][165] = 16'b1111111111101110;
    assign weights1[53][166] = 16'b1111111111111001;
    assign weights1[53][167] = 16'b0000000000000001;
    assign weights1[53][168] = 16'b0000000000000000;
    assign weights1[53][169] = 16'b0000000000000001;
    assign weights1[53][170] = 16'b1111111111111010;
    assign weights1[53][171] = 16'b1111111111110011;
    assign weights1[53][172] = 16'b1111111111101000;
    assign weights1[53][173] = 16'b1111111111100001;
    assign weights1[53][174] = 16'b1111111111100111;
    assign weights1[53][175] = 16'b1111111111111101;
    assign weights1[53][176] = 16'b0000000000000010;
    assign weights1[53][177] = 16'b0000000000000001;
    assign weights1[53][178] = 16'b1111111111111101;
    assign weights1[53][179] = 16'b1111111111011110;
    assign weights1[53][180] = 16'b1111111111111101;
    assign weights1[53][181] = 16'b1111111111110011;
    assign weights1[53][182] = 16'b0000000000001111;
    assign weights1[53][183] = 16'b1111111111111000;
    assign weights1[53][184] = 16'b1111111111100010;
    assign weights1[53][185] = 16'b0000000000010101;
    assign weights1[53][186] = 16'b1111111111101101;
    assign weights1[53][187] = 16'b1111111111110011;
    assign weights1[53][188] = 16'b1111111111100101;
    assign weights1[53][189] = 16'b0000000000000100;
    assign weights1[53][190] = 16'b0000000000000001;
    assign weights1[53][191] = 16'b0000000000000010;
    assign weights1[53][192] = 16'b1111111111111101;
    assign weights1[53][193] = 16'b0000000000001011;
    assign weights1[53][194] = 16'b1111111111101100;
    assign weights1[53][195] = 16'b1111111111111111;
    assign weights1[53][196] = 16'b0000000000000010;
    assign weights1[53][197] = 16'b0000000000000000;
    assign weights1[53][198] = 16'b1111111111111101;
    assign weights1[53][199] = 16'b1111111111110011;
    assign weights1[53][200] = 16'b1111111111100100;
    assign weights1[53][201] = 16'b1111111111110000;
    assign weights1[53][202] = 16'b1111111111100000;
    assign weights1[53][203] = 16'b0000000000001000;
    assign weights1[53][204] = 16'b1111111111110101;
    assign weights1[53][205] = 16'b0000000000000111;
    assign weights1[53][206] = 16'b0000000000011010;
    assign weights1[53][207] = 16'b0000000000010111;
    assign weights1[53][208] = 16'b0000000000001101;
    assign weights1[53][209] = 16'b0000000000011001;
    assign weights1[53][210] = 16'b0000000000000101;
    assign weights1[53][211] = 16'b0000000000000010;
    assign weights1[53][212] = 16'b0000000000100100;
    assign weights1[53][213] = 16'b0000000000010010;
    assign weights1[53][214] = 16'b0000000000010110;
    assign weights1[53][215] = 16'b0000000000100001;
    assign weights1[53][216] = 16'b0000000000001000;
    assign weights1[53][217] = 16'b0000000000010000;
    assign weights1[53][218] = 16'b0000000000010001;
    assign weights1[53][219] = 16'b1111111111110101;
    assign weights1[53][220] = 16'b0000000000000101;
    assign weights1[53][221] = 16'b1111111111110100;
    assign weights1[53][222] = 16'b1111111111101111;
    assign weights1[53][223] = 16'b1111111111111110;
    assign weights1[53][224] = 16'b0000000000000000;
    assign weights1[53][225] = 16'b0000000000000100;
    assign weights1[53][226] = 16'b0000000000000101;
    assign weights1[53][227] = 16'b1111111111111101;
    assign weights1[53][228] = 16'b1111111111101111;
    assign weights1[53][229] = 16'b0000000000000011;
    assign weights1[53][230] = 16'b0000000000000000;
    assign weights1[53][231] = 16'b1111111111110001;
    assign weights1[53][232] = 16'b0000000000001010;
    assign weights1[53][233] = 16'b0000000000000000;
    assign weights1[53][234] = 16'b1111111111100111;
    assign weights1[53][235] = 16'b0000000000000101;
    assign weights1[53][236] = 16'b0000000000010110;
    assign weights1[53][237] = 16'b0000000000001100;
    assign weights1[53][238] = 16'b0000000000000010;
    assign weights1[53][239] = 16'b0000000000001100;
    assign weights1[53][240] = 16'b0000000000000101;
    assign weights1[53][241] = 16'b0000000000010011;
    assign weights1[53][242] = 16'b1111111111110101;
    assign weights1[53][243] = 16'b0000000000001001;
    assign weights1[53][244] = 16'b1111111111100011;
    assign weights1[53][245] = 16'b0000000000001110;
    assign weights1[53][246] = 16'b1111111111111001;
    assign weights1[53][247] = 16'b1111111111110010;
    assign weights1[53][248] = 16'b1111111111111000;
    assign weights1[53][249] = 16'b0000000000000100;
    assign weights1[53][250] = 16'b1111111111101100;
    assign weights1[53][251] = 16'b1111111111111011;
    assign weights1[53][252] = 16'b0000000000000010;
    assign weights1[53][253] = 16'b0000000000000101;
    assign weights1[53][254] = 16'b0000000000010100;
    assign weights1[53][255] = 16'b0000000000001110;
    assign weights1[53][256] = 16'b1111111111110110;
    assign weights1[53][257] = 16'b1111111111101010;
    assign weights1[53][258] = 16'b0000000000001000;
    assign weights1[53][259] = 16'b1111111111101101;
    assign weights1[53][260] = 16'b1111111111101110;
    assign weights1[53][261] = 16'b1111111111101100;
    assign weights1[53][262] = 16'b1111111111101111;
    assign weights1[53][263] = 16'b1111111111111100;
    assign weights1[53][264] = 16'b1111111111111110;
    assign weights1[53][265] = 16'b0000000000001010;
    assign weights1[53][266] = 16'b0000000000001011;
    assign weights1[53][267] = 16'b0000000000001011;
    assign weights1[53][268] = 16'b0000000000000110;
    assign weights1[53][269] = 16'b0000000000011000;
    assign weights1[53][270] = 16'b0000000000001100;
    assign weights1[53][271] = 16'b0000000000001000;
    assign weights1[53][272] = 16'b1111111111101100;
    assign weights1[53][273] = 16'b1111111111111011;
    assign weights1[53][274] = 16'b1111111111111000;
    assign weights1[53][275] = 16'b1111111111110001;
    assign weights1[53][276] = 16'b1111111111111111;
    assign weights1[53][277] = 16'b0000000000001010;
    assign weights1[53][278] = 16'b1111111111111001;
    assign weights1[53][279] = 16'b0000000000000010;
    assign weights1[53][280] = 16'b0000000000000111;
    assign weights1[53][281] = 16'b0000000000001000;
    assign weights1[53][282] = 16'b0000000000001010;
    assign weights1[53][283] = 16'b0000000000001110;
    assign weights1[53][284] = 16'b0000000000010011;
    assign weights1[53][285] = 16'b0000000000001011;
    assign weights1[53][286] = 16'b0000000000011111;
    assign weights1[53][287] = 16'b0000000000000110;
    assign weights1[53][288] = 16'b0000000000001000;
    assign weights1[53][289] = 16'b0000000000000101;
    assign weights1[53][290] = 16'b0000000000010011;
    assign weights1[53][291] = 16'b1111111111101001;
    assign weights1[53][292] = 16'b1111111111111101;
    assign weights1[53][293] = 16'b1111111111111101;
    assign weights1[53][294] = 16'b1111111111110110;
    assign weights1[53][295] = 16'b1111111111111000;
    assign weights1[53][296] = 16'b0000000000001101;
    assign weights1[53][297] = 16'b0000000000000000;
    assign weights1[53][298] = 16'b1111111111110000;
    assign weights1[53][299] = 16'b1111111111111010;
    assign weights1[53][300] = 16'b0000000000001011;
    assign weights1[53][301] = 16'b0000000000001000;
    assign weights1[53][302] = 16'b1111111111111110;
    assign weights1[53][303] = 16'b1111111111101101;
    assign weights1[53][304] = 16'b1111111111110111;
    assign weights1[53][305] = 16'b0000000000001111;
    assign weights1[53][306] = 16'b0000000000000001;
    assign weights1[53][307] = 16'b0000000000000110;
    assign weights1[53][308] = 16'b0000000000001111;
    assign weights1[53][309] = 16'b0000000000010000;
    assign weights1[53][310] = 16'b0000000000110000;
    assign weights1[53][311] = 16'b0000000000101100;
    assign weights1[53][312] = 16'b0000000000011110;
    assign weights1[53][313] = 16'b0000000000010010;
    assign weights1[53][314] = 16'b0000000000000101;
    assign weights1[53][315] = 16'b0000000000000110;
    assign weights1[53][316] = 16'b0000000000011100;
    assign weights1[53][317] = 16'b0000000000010011;
    assign weights1[53][318] = 16'b0000000000001110;
    assign weights1[53][319] = 16'b0000000000001000;
    assign weights1[53][320] = 16'b0000000000000101;
    assign weights1[53][321] = 16'b1111111111101100;
    assign weights1[53][322] = 16'b1111111111110111;
    assign weights1[53][323] = 16'b1111111111111001;
    assign weights1[53][324] = 16'b1111111111111101;
    assign weights1[53][325] = 16'b1111111111111110;
    assign weights1[53][326] = 16'b0000000000001001;
    assign weights1[53][327] = 16'b1111111111110000;
    assign weights1[53][328] = 16'b0000000000001010;
    assign weights1[53][329] = 16'b1111111111111100;
    assign weights1[53][330] = 16'b1111111111101100;
    assign weights1[53][331] = 16'b1111111111011000;
    assign weights1[53][332] = 16'b0000000000000110;
    assign weights1[53][333] = 16'b0000000000000110;
    assign weights1[53][334] = 16'b0000000000001101;
    assign weights1[53][335] = 16'b0000000000011100;
    assign weights1[53][336] = 16'b0000000000001101;
    assign weights1[53][337] = 16'b0000000000001011;
    assign weights1[53][338] = 16'b0000000000101111;
    assign weights1[53][339] = 16'b0000000000100111;
    assign weights1[53][340] = 16'b0000000000101011;
    assign weights1[53][341] = 16'b0000000000100001;
    assign weights1[53][342] = 16'b0000000000100000;
    assign weights1[53][343] = 16'b0000000000100100;
    assign weights1[53][344] = 16'b0000000000000011;
    assign weights1[53][345] = 16'b0000000000100111;
    assign weights1[53][346] = 16'b0000000000001100;
    assign weights1[53][347] = 16'b0000000000001011;
    assign weights1[53][348] = 16'b1111111111111101;
    assign weights1[53][349] = 16'b0000000000001001;
    assign weights1[53][350] = 16'b1111111111111111;
    assign weights1[53][351] = 16'b1111111111110011;
    assign weights1[53][352] = 16'b0000000000000010;
    assign weights1[53][353] = 16'b0000000000001001;
    assign weights1[53][354] = 16'b1111111111111100;
    assign weights1[53][355] = 16'b1111111111111000;
    assign weights1[53][356] = 16'b1111111111101011;
    assign weights1[53][357] = 16'b1111111111111111;
    assign weights1[53][358] = 16'b1111111111110000;
    assign weights1[53][359] = 16'b1111111111110011;
    assign weights1[53][360] = 16'b1111111111101111;
    assign weights1[53][361] = 16'b1111111111111011;
    assign weights1[53][362] = 16'b0000000000010010;
    assign weights1[53][363] = 16'b0000000000001000;
    assign weights1[53][364] = 16'b0000000000001110;
    assign weights1[53][365] = 16'b0000000000011100;
    assign weights1[53][366] = 16'b0000000000101100;
    assign weights1[53][367] = 16'b0000000000100001;
    assign weights1[53][368] = 16'b0000000000100111;
    assign weights1[53][369] = 16'b0000000001000001;
    assign weights1[53][370] = 16'b0000000000010100;
    assign weights1[53][371] = 16'b0000000000011111;
    assign weights1[53][372] = 16'b0000000000001001;
    assign weights1[53][373] = 16'b0000000000011000;
    assign weights1[53][374] = 16'b0000000000100101;
    assign weights1[53][375] = 16'b0000000000010101;
    assign weights1[53][376] = 16'b0000000000000111;
    assign weights1[53][377] = 16'b0000000000010010;
    assign weights1[53][378] = 16'b1111111111110011;
    assign weights1[53][379] = 16'b0000000000011000;
    assign weights1[53][380] = 16'b0000000000001010;
    assign weights1[53][381] = 16'b0000000000010011;
    assign weights1[53][382] = 16'b0000000000001101;
    assign weights1[53][383] = 16'b1111111111111111;
    assign weights1[53][384] = 16'b0000000000101001;
    assign weights1[53][385] = 16'b1111111111111011;
    assign weights1[53][386] = 16'b0000000000000100;
    assign weights1[53][387] = 16'b0000000000000101;
    assign weights1[53][388] = 16'b1111111111111110;
    assign weights1[53][389] = 16'b0000000000000110;
    assign weights1[53][390] = 16'b0000000000000011;
    assign weights1[53][391] = 16'b0000000000010000;
    assign weights1[53][392] = 16'b0000000000001001;
    assign weights1[53][393] = 16'b0000000000011010;
    assign weights1[53][394] = 16'b0000000000110001;
    assign weights1[53][395] = 16'b0000000000011111;
    assign weights1[53][396] = 16'b0000000000011101;
    assign weights1[53][397] = 16'b0000000000101110;
    assign weights1[53][398] = 16'b0000000000101100;
    assign weights1[53][399] = 16'b0000000000111101;
    assign weights1[53][400] = 16'b0000000000100110;
    assign weights1[53][401] = 16'b0000000000110111;
    assign weights1[53][402] = 16'b0000000000000100;
    assign weights1[53][403] = 16'b0000000000001011;
    assign weights1[53][404] = 16'b0000000000000110;
    assign weights1[53][405] = 16'b0000000000010010;
    assign weights1[53][406] = 16'b0000000000010001;
    assign weights1[53][407] = 16'b0000000000001001;
    assign weights1[53][408] = 16'b0000000000001111;
    assign weights1[53][409] = 16'b0000000000001100;
    assign weights1[53][410] = 16'b0000000000001110;
    assign weights1[53][411] = 16'b0000000000011011;
    assign weights1[53][412] = 16'b0000000000010001;
    assign weights1[53][413] = 16'b0000000000001111;
    assign weights1[53][414] = 16'b0000000000011000;
    assign weights1[53][415] = 16'b0000000000100111;
    assign weights1[53][416] = 16'b0000000000001100;
    assign weights1[53][417] = 16'b0000000000011100;
    assign weights1[53][418] = 16'b0000000000010001;
    assign weights1[53][419] = 16'b0000000000000000;
    assign weights1[53][420] = 16'b0000000000001001;
    assign weights1[53][421] = 16'b0000000000001010;
    assign weights1[53][422] = 16'b0000000000011001;
    assign weights1[53][423] = 16'b0000000000011000;
    assign weights1[53][424] = 16'b0000000000101101;
    assign weights1[53][425] = 16'b0000000000110011;
    assign weights1[53][426] = 16'b0000000000011000;
    assign weights1[53][427] = 16'b0000000000110010;
    assign weights1[53][428] = 16'b0000000000101011;
    assign weights1[53][429] = 16'b0000000000011110;
    assign weights1[53][430] = 16'b0000000000010010;
    assign weights1[53][431] = 16'b0000000000010100;
    assign weights1[53][432] = 16'b0000000000001100;
    assign weights1[53][433] = 16'b0000000000000101;
    assign weights1[53][434] = 16'b0000000000011000;
    assign weights1[53][435] = 16'b0000000000100010;
    assign weights1[53][436] = 16'b0000000000011100;
    assign weights1[53][437] = 16'b0000000000100011;
    assign weights1[53][438] = 16'b0000000000011101;
    assign weights1[53][439] = 16'b0000000000010100;
    assign weights1[53][440] = 16'b0000000000101010;
    assign weights1[53][441] = 16'b0000000000101000;
    assign weights1[53][442] = 16'b0000000000010101;
    assign weights1[53][443] = 16'b0000000000011100;
    assign weights1[53][444] = 16'b0000000000001011;
    assign weights1[53][445] = 16'b1111111111111101;
    assign weights1[53][446] = 16'b0000000000001001;
    assign weights1[53][447] = 16'b0000000000001001;
    assign weights1[53][448] = 16'b1111111111111111;
    assign weights1[53][449] = 16'b0000000000000011;
    assign weights1[53][450] = 16'b0000000000000100;
    assign weights1[53][451] = 16'b0000000000000011;
    assign weights1[53][452] = 16'b0000000000010011;
    assign weights1[53][453] = 16'b0000000000011001;
    assign weights1[53][454] = 16'b0000000000010010;
    assign weights1[53][455] = 16'b0000000000010110;
    assign weights1[53][456] = 16'b0000000000100011;
    assign weights1[53][457] = 16'b0000000000001000;
    assign weights1[53][458] = 16'b0000000000010001;
    assign weights1[53][459] = 16'b0000000000001000;
    assign weights1[53][460] = 16'b0000000000011101;
    assign weights1[53][461] = 16'b0000000000010100;
    assign weights1[53][462] = 16'b0000000000001111;
    assign weights1[53][463] = 16'b0000000000011010;
    assign weights1[53][464] = 16'b0000000000011001;
    assign weights1[53][465] = 16'b0000000000100010;
    assign weights1[53][466] = 16'b0000000000001011;
    assign weights1[53][467] = 16'b0000000000001111;
    assign weights1[53][468] = 16'b0000000000010000;
    assign weights1[53][469] = 16'b0000000000011000;
    assign weights1[53][470] = 16'b1111111111111011;
    assign weights1[53][471] = 16'b0000000000001010;
    assign weights1[53][472] = 16'b0000000000001010;
    assign weights1[53][473] = 16'b0000000000000000;
    assign weights1[53][474] = 16'b1111111111111110;
    assign weights1[53][475] = 16'b0000000000000000;
    assign weights1[53][476] = 16'b1111111111101111;
    assign weights1[53][477] = 16'b1111111111101001;
    assign weights1[53][478] = 16'b1111111111100111;
    assign weights1[53][479] = 16'b1111111111101111;
    assign weights1[53][480] = 16'b1111111111110011;
    assign weights1[53][481] = 16'b1111111111110111;
    assign weights1[53][482] = 16'b1111111111110110;
    assign weights1[53][483] = 16'b1111111111110011;
    assign weights1[53][484] = 16'b1111111111110101;
    assign weights1[53][485] = 16'b1111111111100111;
    assign weights1[53][486] = 16'b1111111111110010;
    assign weights1[53][487] = 16'b0000000000011001;
    assign weights1[53][488] = 16'b1111111111111111;
    assign weights1[53][489] = 16'b0000000000001000;
    assign weights1[53][490] = 16'b0000000000000110;
    assign weights1[53][491] = 16'b0000000000001000;
    assign weights1[53][492] = 16'b0000000000000000;
    assign weights1[53][493] = 16'b0000000000000110;
    assign weights1[53][494] = 16'b0000000000001011;
    assign weights1[53][495] = 16'b1111111111110110;
    assign weights1[53][496] = 16'b0000000000000011;
    assign weights1[53][497] = 16'b0000000000000110;
    assign weights1[53][498] = 16'b1111111111101011;
    assign weights1[53][499] = 16'b1111111111111000;
    assign weights1[53][500] = 16'b1111111111101101;
    assign weights1[53][501] = 16'b1111111111111000;
    assign weights1[53][502] = 16'b1111111111111011;
    assign weights1[53][503] = 16'b1111111111111110;
    assign weights1[53][504] = 16'b1111111111100001;
    assign weights1[53][505] = 16'b1111111111010100;
    assign weights1[53][506] = 16'b1111111111001110;
    assign weights1[53][507] = 16'b1111111111000100;
    assign weights1[53][508] = 16'b1111111111011110;
    assign weights1[53][509] = 16'b1111111111010101;
    assign weights1[53][510] = 16'b1111111111010011;
    assign weights1[53][511] = 16'b1111111111001010;
    assign weights1[53][512] = 16'b1111111111000111;
    assign weights1[53][513] = 16'b1111111110111101;
    assign weights1[53][514] = 16'b1111111111010000;
    assign weights1[53][515] = 16'b1111111111011000;
    assign weights1[53][516] = 16'b1111111111011011;
    assign weights1[53][517] = 16'b1111111111100100;
    assign weights1[53][518] = 16'b1111111111101111;
    assign weights1[53][519] = 16'b1111111111111011;
    assign weights1[53][520] = 16'b1111111111110100;
    assign weights1[53][521] = 16'b1111111111110011;
    assign weights1[53][522] = 16'b1111111111110011;
    assign weights1[53][523] = 16'b1111111111100111;
    assign weights1[53][524] = 16'b1111111111110101;
    assign weights1[53][525] = 16'b1111111111101100;
    assign weights1[53][526] = 16'b1111111111001111;
    assign weights1[53][527] = 16'b1111111111011111;
    assign weights1[53][528] = 16'b1111111111011011;
    assign weights1[53][529] = 16'b1111111111101111;
    assign weights1[53][530] = 16'b1111111111110000;
    assign weights1[53][531] = 16'b1111111111111110;
    assign weights1[53][532] = 16'b1111111111011100;
    assign weights1[53][533] = 16'b1111111111010000;
    assign weights1[53][534] = 16'b1111111111000001;
    assign weights1[53][535] = 16'b1111111110101010;
    assign weights1[53][536] = 16'b1111111110110000;
    assign weights1[53][537] = 16'b1111111110001110;
    assign weights1[53][538] = 16'b1111111101110000;
    assign weights1[53][539] = 16'b1111111101111000;
    assign weights1[53][540] = 16'b1111111101111000;
    assign weights1[53][541] = 16'b1111111110101110;
    assign weights1[53][542] = 16'b1111111111000110;
    assign weights1[53][543] = 16'b1111111111001100;
    assign weights1[53][544] = 16'b1111111111001111;
    assign weights1[53][545] = 16'b1111111111100111;
    assign weights1[53][546] = 16'b1111111111111010;
    assign weights1[53][547] = 16'b1111111111100110;
    assign weights1[53][548] = 16'b1111111111101010;
    assign weights1[53][549] = 16'b1111111111111110;
    assign weights1[53][550] = 16'b1111111111100000;
    assign weights1[53][551] = 16'b1111111111110011;
    assign weights1[53][552] = 16'b1111111111100010;
    assign weights1[53][553] = 16'b1111111111011100;
    assign weights1[53][554] = 16'b1111111111010010;
    assign weights1[53][555] = 16'b1111111111010110;
    assign weights1[53][556] = 16'b1111111111011111;
    assign weights1[53][557] = 16'b1111111111111100;
    assign weights1[53][558] = 16'b1111111111110111;
    assign weights1[53][559] = 16'b1111111111111110;
    assign weights1[53][560] = 16'b1111111111011001;
    assign weights1[53][561] = 16'b1111111111010010;
    assign weights1[53][562] = 16'b1111111111000101;
    assign weights1[53][563] = 16'b1111111110110000;
    assign weights1[53][564] = 16'b1111111110011011;
    assign weights1[53][565] = 16'b1111111110010011;
    assign weights1[53][566] = 16'b1111111110010011;
    assign weights1[53][567] = 16'b1111111110100111;
    assign weights1[53][568] = 16'b1111111111010000;
    assign weights1[53][569] = 16'b1111111111111000;
    assign weights1[53][570] = 16'b1111111111111100;
    assign weights1[53][571] = 16'b0000000000000000;
    assign weights1[53][572] = 16'b0000000000000011;
    assign weights1[53][573] = 16'b0000000000000101;
    assign weights1[53][574] = 16'b0000000000001100;
    assign weights1[53][575] = 16'b0000000000010011;
    assign weights1[53][576] = 16'b1111111111100111;
    assign weights1[53][577] = 16'b1111111111111010;
    assign weights1[53][578] = 16'b0000000000000101;
    assign weights1[53][579] = 16'b1111111111011001;
    assign weights1[53][580] = 16'b1111111111010010;
    assign weights1[53][581] = 16'b1111111111100011;
    assign weights1[53][582] = 16'b1111111111101001;
    assign weights1[53][583] = 16'b1111111111100010;
    assign weights1[53][584] = 16'b0000000000000001;
    assign weights1[53][585] = 16'b1111111111111011;
    assign weights1[53][586] = 16'b1111111111110111;
    assign weights1[53][587] = 16'b1111111111111011;
    assign weights1[53][588] = 16'b1111111111100011;
    assign weights1[53][589] = 16'b1111111111011000;
    assign weights1[53][590] = 16'b1111111111001110;
    assign weights1[53][591] = 16'b1111111110110111;
    assign weights1[53][592] = 16'b1111111110101101;
    assign weights1[53][593] = 16'b1111111110101100;
    assign weights1[53][594] = 16'b1111111111000101;
    assign weights1[53][595] = 16'b0000000000000100;
    assign weights1[53][596] = 16'b0000000000010100;
    assign weights1[53][597] = 16'b0000000000100011;
    assign weights1[53][598] = 16'b0000000000011000;
    assign weights1[53][599] = 16'b0000000000001101;
    assign weights1[53][600] = 16'b0000000000001000;
    assign weights1[53][601] = 16'b1111111111101010;
    assign weights1[53][602] = 16'b1111111111101110;
    assign weights1[53][603] = 16'b1111111111110111;
    assign weights1[53][604] = 16'b1111111111011101;
    assign weights1[53][605] = 16'b1111111111100100;
    assign weights1[53][606] = 16'b1111111111110100;
    assign weights1[53][607] = 16'b1111111111011111;
    assign weights1[53][608] = 16'b1111111111101010;
    assign weights1[53][609] = 16'b1111111111111111;
    assign weights1[53][610] = 16'b1111111111100000;
    assign weights1[53][611] = 16'b1111111111011111;
    assign weights1[53][612] = 16'b1111111111111000;
    assign weights1[53][613] = 16'b1111111111111000;
    assign weights1[53][614] = 16'b1111111111110100;
    assign weights1[53][615] = 16'b1111111111111110;
    assign weights1[53][616] = 16'b1111111111100001;
    assign weights1[53][617] = 16'b1111111111010000;
    assign weights1[53][618] = 16'b1111111111001010;
    assign weights1[53][619] = 16'b1111111111000100;
    assign weights1[53][620] = 16'b1111111111001110;
    assign weights1[53][621] = 16'b1111111111101000;
    assign weights1[53][622] = 16'b0000000000000000;
    assign weights1[53][623] = 16'b0000000000100110;
    assign weights1[53][624] = 16'b0000000000110100;
    assign weights1[53][625] = 16'b0000000000000111;
    assign weights1[53][626] = 16'b0000000000011000;
    assign weights1[53][627] = 16'b1111111111111001;
    assign weights1[53][628] = 16'b1111111111110110;
    assign weights1[53][629] = 16'b1111111111110011;
    assign weights1[53][630] = 16'b1111111111111010;
    assign weights1[53][631] = 16'b1111111111110101;
    assign weights1[53][632] = 16'b1111111111111010;
    assign weights1[53][633] = 16'b1111111111111101;
    assign weights1[53][634] = 16'b1111111111110111;
    assign weights1[53][635] = 16'b1111111111101100;
    assign weights1[53][636] = 16'b1111111111110001;
    assign weights1[53][637] = 16'b1111111111111101;
    assign weights1[53][638] = 16'b1111111111101101;
    assign weights1[53][639] = 16'b1111111111100110;
    assign weights1[53][640] = 16'b1111111111111001;
    assign weights1[53][641] = 16'b1111111111101101;
    assign weights1[53][642] = 16'b0000000000000000;
    assign weights1[53][643] = 16'b0000000000000000;
    assign weights1[53][644] = 16'b1111111111011111;
    assign weights1[53][645] = 16'b1111111111011111;
    assign weights1[53][646] = 16'b1111111111010101;
    assign weights1[53][647] = 16'b1111111111001110;
    assign weights1[53][648] = 16'b1111111111011010;
    assign weights1[53][649] = 16'b1111111111111010;
    assign weights1[53][650] = 16'b0000000000100000;
    assign weights1[53][651] = 16'b0000000000011011;
    assign weights1[53][652] = 16'b0000000000000100;
    assign weights1[53][653] = 16'b1111111111110111;
    assign weights1[53][654] = 16'b1111111111110101;
    assign weights1[53][655] = 16'b0000000000000111;
    assign weights1[53][656] = 16'b1111111111111000;
    assign weights1[53][657] = 16'b0000000000001100;
    assign weights1[53][658] = 16'b1111111111111000;
    assign weights1[53][659] = 16'b1111111111011001;
    assign weights1[53][660] = 16'b1111111111101111;
    assign weights1[53][661] = 16'b0000000000010111;
    assign weights1[53][662] = 16'b1111111111111001;
    assign weights1[53][663] = 16'b1111111111100101;
    assign weights1[53][664] = 16'b1111111111011100;
    assign weights1[53][665] = 16'b1111111111101010;
    assign weights1[53][666] = 16'b1111111111011100;
    assign weights1[53][667] = 16'b1111111111011111;
    assign weights1[53][668] = 16'b1111111111110011;
    assign weights1[53][669] = 16'b1111111111111111;
    assign weights1[53][670] = 16'b0000000000000000;
    assign weights1[53][671] = 16'b1111111111111111;
    assign weights1[53][672] = 16'b1111111111101110;
    assign weights1[53][673] = 16'b1111111111101000;
    assign weights1[53][674] = 16'b1111111111100000;
    assign weights1[53][675] = 16'b1111111111110110;
    assign weights1[53][676] = 16'b1111111111111011;
    assign weights1[53][677] = 16'b0000000000010011;
    assign weights1[53][678] = 16'b0000000000100000;
    assign weights1[53][679] = 16'b0000000000100100;
    assign weights1[53][680] = 16'b0000000000001101;
    assign weights1[53][681] = 16'b0000000000001100;
    assign weights1[53][682] = 16'b1111111111110101;
    assign weights1[53][683] = 16'b1111111111110101;
    assign weights1[53][684] = 16'b1111111111110101;
    assign weights1[53][685] = 16'b0000000000000100;
    assign weights1[53][686] = 16'b1111111111111100;
    assign weights1[53][687] = 16'b1111111111010101;
    assign weights1[53][688] = 16'b1111111111111000;
    assign weights1[53][689] = 16'b1111111111110100;
    assign weights1[53][690] = 16'b1111111111111010;
    assign weights1[53][691] = 16'b1111111111010101;
    assign weights1[53][692] = 16'b1111111111111011;
    assign weights1[53][693] = 16'b1111111111110111;
    assign weights1[53][694] = 16'b1111111111110111;
    assign weights1[53][695] = 16'b1111111111111100;
    assign weights1[53][696] = 16'b1111111111110011;
    assign weights1[53][697] = 16'b1111111111110101;
    assign weights1[53][698] = 16'b1111111111111011;
    assign weights1[53][699] = 16'b1111111111111110;
    assign weights1[53][700] = 16'b1111111111111001;
    assign weights1[53][701] = 16'b1111111111110010;
    assign weights1[53][702] = 16'b1111111111110101;
    assign weights1[53][703] = 16'b1111111111111010;
    assign weights1[53][704] = 16'b0000000000011101;
    assign weights1[53][705] = 16'b0000000000010111;
    assign weights1[53][706] = 16'b0000000000010111;
    assign weights1[53][707] = 16'b0000000000000011;
    assign weights1[53][708] = 16'b0000000000001100;
    assign weights1[53][709] = 16'b1111111111110010;
    assign weights1[53][710] = 16'b1111111111110101;
    assign weights1[53][711] = 16'b1111111111110111;
    assign weights1[53][712] = 16'b1111111111011111;
    assign weights1[53][713] = 16'b0000000000001001;
    assign weights1[53][714] = 16'b1111111111111100;
    assign weights1[53][715] = 16'b0000000000000101;
    assign weights1[53][716] = 16'b0000000000011001;
    assign weights1[53][717] = 16'b0000000000000100;
    assign weights1[53][718] = 16'b0000000000000100;
    assign weights1[53][719] = 16'b1111111111110110;
    assign weights1[53][720] = 16'b1111111111101110;
    assign weights1[53][721] = 16'b1111111111111000;
    assign weights1[53][722] = 16'b0000000000000001;
    assign weights1[53][723] = 16'b0000000000000100;
    assign weights1[53][724] = 16'b1111111111111101;
    assign weights1[53][725] = 16'b1111111111111101;
    assign weights1[53][726] = 16'b1111111111111111;
    assign weights1[53][727] = 16'b1111111111111101;
    assign weights1[53][728] = 16'b1111111111111100;
    assign weights1[53][729] = 16'b1111111111111010;
    assign weights1[53][730] = 16'b1111111111111111;
    assign weights1[53][731] = 16'b0000000000000100;
    assign weights1[53][732] = 16'b0000000000011001;
    assign weights1[53][733] = 16'b0000000000010010;
    assign weights1[53][734] = 16'b0000000000010000;
    assign weights1[53][735] = 16'b1111111111110101;
    assign weights1[53][736] = 16'b1111111111101111;
    assign weights1[53][737] = 16'b1111111111111010;
    assign weights1[53][738] = 16'b1111111111101110;
    assign weights1[53][739] = 16'b1111111111110011;
    assign weights1[53][740] = 16'b0000000000000111;
    assign weights1[53][741] = 16'b0000000000000110;
    assign weights1[53][742] = 16'b1111111111111100;
    assign weights1[53][743] = 16'b1111111111101110;
    assign weights1[53][744] = 16'b0000000000000111;
    assign weights1[53][745] = 16'b1111111111111110;
    assign weights1[53][746] = 16'b1111111111110000;
    assign weights1[53][747] = 16'b1111111111110011;
    assign weights1[53][748] = 16'b1111111111101110;
    assign weights1[53][749] = 16'b1111111111110010;
    assign weights1[53][750] = 16'b1111111111110100;
    assign weights1[53][751] = 16'b1111111111111011;
    assign weights1[53][752] = 16'b1111111111111110;
    assign weights1[53][753] = 16'b0000000000000001;
    assign weights1[53][754] = 16'b0000000000000000;
    assign weights1[53][755] = 16'b0000000000000000;
    assign weights1[53][756] = 16'b1111111111111111;
    assign weights1[53][757] = 16'b1111111111111111;
    assign weights1[53][758] = 16'b0000000000000101;
    assign weights1[53][759] = 16'b0000000000001000;
    assign weights1[53][760] = 16'b0000000000010000;
    assign weights1[53][761] = 16'b0000000000000011;
    assign weights1[53][762] = 16'b1111111111110110;
    assign weights1[53][763] = 16'b1111111111110010;
    assign weights1[53][764] = 16'b1111111111101000;
    assign weights1[53][765] = 16'b1111111111101101;
    assign weights1[53][766] = 16'b1111111111111000;
    assign weights1[53][767] = 16'b1111111111110001;
    assign weights1[53][768] = 16'b1111111111100100;
    assign weights1[53][769] = 16'b1111111111101110;
    assign weights1[53][770] = 16'b1111111111110000;
    assign weights1[53][771] = 16'b1111111111101101;
    assign weights1[53][772] = 16'b1111111111111001;
    assign weights1[53][773] = 16'b1111111111111101;
    assign weights1[53][774] = 16'b1111111111110100;
    assign weights1[53][775] = 16'b1111111111110111;
    assign weights1[53][776] = 16'b1111111111111000;
    assign weights1[53][777] = 16'b1111111111110001;
    assign weights1[53][778] = 16'b1111111111111000;
    assign weights1[53][779] = 16'b1111111111110111;
    assign weights1[53][780] = 16'b1111111111111011;
    assign weights1[53][781] = 16'b1111111111111101;
    assign weights1[53][782] = 16'b1111111111111111;
    assign weights1[53][783] = 16'b0000000000000001;
    assign weights1[54][0] = 16'b0000000000000000;
    assign weights1[54][1] = 16'b0000000000000000;
    assign weights1[54][2] = 16'b0000000000000000;
    assign weights1[54][3] = 16'b0000000000000000;
    assign weights1[54][4] = 16'b0000000000000000;
    assign weights1[54][5] = 16'b0000000000000000;
    assign weights1[54][6] = 16'b0000000000000000;
    assign weights1[54][7] = 16'b0000000000000000;
    assign weights1[54][8] = 16'b0000000000000000;
    assign weights1[54][9] = 16'b0000000000000000;
    assign weights1[54][10] = 16'b0000000000000000;
    assign weights1[54][11] = 16'b0000000000000000;
    assign weights1[54][12] = 16'b0000000000000000;
    assign weights1[54][13] = 16'b0000000000000000;
    assign weights1[54][14] = 16'b0000000000000000;
    assign weights1[54][15] = 16'b0000000000000000;
    assign weights1[54][16] = 16'b0000000000000000;
    assign weights1[54][17] = 16'b0000000000000000;
    assign weights1[54][18] = 16'b0000000000000000;
    assign weights1[54][19] = 16'b0000000000000000;
    assign weights1[54][20] = 16'b0000000000000000;
    assign weights1[54][21] = 16'b0000000000000000;
    assign weights1[54][22] = 16'b0000000000000000;
    assign weights1[54][23] = 16'b0000000000000000;
    assign weights1[54][24] = 16'b0000000000000000;
    assign weights1[54][25] = 16'b0000000000000000;
    assign weights1[54][26] = 16'b0000000000000000;
    assign weights1[54][27] = 16'b0000000000000000;
    assign weights1[54][28] = 16'b0000000000000000;
    assign weights1[54][29] = 16'b0000000000000000;
    assign weights1[54][30] = 16'b0000000000000000;
    assign weights1[54][31] = 16'b0000000000000000;
    assign weights1[54][32] = 16'b0000000000000000;
    assign weights1[54][33] = 16'b0000000000000000;
    assign weights1[54][34] = 16'b0000000000000000;
    assign weights1[54][35] = 16'b0000000000000000;
    assign weights1[54][36] = 16'b0000000000000000;
    assign weights1[54][37] = 16'b0000000000000000;
    assign weights1[54][38] = 16'b0000000000000000;
    assign weights1[54][39] = 16'b0000000000000000;
    assign weights1[54][40] = 16'b0000000000000000;
    assign weights1[54][41] = 16'b0000000000000000;
    assign weights1[54][42] = 16'b0000000000000000;
    assign weights1[54][43] = 16'b0000000000000000;
    assign weights1[54][44] = 16'b0000000000000000;
    assign weights1[54][45] = 16'b0000000000000000;
    assign weights1[54][46] = 16'b0000000000000000;
    assign weights1[54][47] = 16'b0000000000000000;
    assign weights1[54][48] = 16'b0000000000000000;
    assign weights1[54][49] = 16'b0000000000000000;
    assign weights1[54][50] = 16'b0000000000000000;
    assign weights1[54][51] = 16'b0000000000000000;
    assign weights1[54][52] = 16'b0000000000000000;
    assign weights1[54][53] = 16'b0000000000000000;
    assign weights1[54][54] = 16'b0000000000000000;
    assign weights1[54][55] = 16'b0000000000000000;
    assign weights1[54][56] = 16'b0000000000000000;
    assign weights1[54][57] = 16'b0000000000000000;
    assign weights1[54][58] = 16'b0000000000000000;
    assign weights1[54][59] = 16'b0000000000000000;
    assign weights1[54][60] = 16'b0000000000000000;
    assign weights1[54][61] = 16'b0000000000000000;
    assign weights1[54][62] = 16'b0000000000000000;
    assign weights1[54][63] = 16'b0000000000000000;
    assign weights1[54][64] = 16'b0000000000000000;
    assign weights1[54][65] = 16'b0000000000000000;
    assign weights1[54][66] = 16'b0000000000000000;
    assign weights1[54][67] = 16'b0000000000000000;
    assign weights1[54][68] = 16'b0000000000000000;
    assign weights1[54][69] = 16'b0000000000000000;
    assign weights1[54][70] = 16'b0000000000000000;
    assign weights1[54][71] = 16'b0000000000000000;
    assign weights1[54][72] = 16'b0000000000000000;
    assign weights1[54][73] = 16'b0000000000000000;
    assign weights1[54][74] = 16'b0000000000000000;
    assign weights1[54][75] = 16'b0000000000000000;
    assign weights1[54][76] = 16'b0000000000000000;
    assign weights1[54][77] = 16'b0000000000000000;
    assign weights1[54][78] = 16'b0000000000000000;
    assign weights1[54][79] = 16'b0000000000000000;
    assign weights1[54][80] = 16'b0000000000000000;
    assign weights1[54][81] = 16'b0000000000000000;
    assign weights1[54][82] = 16'b0000000000000000;
    assign weights1[54][83] = 16'b0000000000000000;
    assign weights1[54][84] = 16'b0000000000000000;
    assign weights1[54][85] = 16'b0000000000000000;
    assign weights1[54][86] = 16'b0000000000000000;
    assign weights1[54][87] = 16'b0000000000000000;
    assign weights1[54][88] = 16'b0000000000000000;
    assign weights1[54][89] = 16'b0000000000000000;
    assign weights1[54][90] = 16'b0000000000000000;
    assign weights1[54][91] = 16'b0000000000000000;
    assign weights1[54][92] = 16'b0000000000000000;
    assign weights1[54][93] = 16'b0000000000000000;
    assign weights1[54][94] = 16'b0000000000000000;
    assign weights1[54][95] = 16'b0000000000000000;
    assign weights1[54][96] = 16'b0000000000000000;
    assign weights1[54][97] = 16'b0000000000000000;
    assign weights1[54][98] = 16'b0000000000000000;
    assign weights1[54][99] = 16'b0000000000000000;
    assign weights1[54][100] = 16'b0000000000000000;
    assign weights1[54][101] = 16'b0000000000000000;
    assign weights1[54][102] = 16'b0000000000000000;
    assign weights1[54][103] = 16'b0000000000000000;
    assign weights1[54][104] = 16'b0000000000000000;
    assign weights1[54][105] = 16'b0000000000000000;
    assign weights1[54][106] = 16'b0000000000000000;
    assign weights1[54][107] = 16'b0000000000000000;
    assign weights1[54][108] = 16'b0000000000000000;
    assign weights1[54][109] = 16'b0000000000000000;
    assign weights1[54][110] = 16'b0000000000000000;
    assign weights1[54][111] = 16'b0000000000000000;
    assign weights1[54][112] = 16'b0000000000000000;
    assign weights1[54][113] = 16'b0000000000000000;
    assign weights1[54][114] = 16'b0000000000000000;
    assign weights1[54][115] = 16'b0000000000000000;
    assign weights1[54][116] = 16'b0000000000000000;
    assign weights1[54][117] = 16'b0000000000000000;
    assign weights1[54][118] = 16'b0000000000000000;
    assign weights1[54][119] = 16'b0000000000000000;
    assign weights1[54][120] = 16'b0000000000000000;
    assign weights1[54][121] = 16'b0000000000000000;
    assign weights1[54][122] = 16'b0000000000000000;
    assign weights1[54][123] = 16'b0000000000000000;
    assign weights1[54][124] = 16'b0000000000000000;
    assign weights1[54][125] = 16'b0000000000000000;
    assign weights1[54][126] = 16'b0000000000000000;
    assign weights1[54][127] = 16'b0000000000000000;
    assign weights1[54][128] = 16'b0000000000000000;
    assign weights1[54][129] = 16'b0000000000000000;
    assign weights1[54][130] = 16'b0000000000000000;
    assign weights1[54][131] = 16'b0000000000000000;
    assign weights1[54][132] = 16'b0000000000000000;
    assign weights1[54][133] = 16'b0000000000000000;
    assign weights1[54][134] = 16'b0000000000000000;
    assign weights1[54][135] = 16'b0000000000000000;
    assign weights1[54][136] = 16'b0000000000000000;
    assign weights1[54][137] = 16'b0000000000000000;
    assign weights1[54][138] = 16'b0000000000000000;
    assign weights1[54][139] = 16'b0000000000000000;
    assign weights1[54][140] = 16'b0000000000000000;
    assign weights1[54][141] = 16'b0000000000000000;
    assign weights1[54][142] = 16'b0000000000000000;
    assign weights1[54][143] = 16'b0000000000000000;
    assign weights1[54][144] = 16'b0000000000000000;
    assign weights1[54][145] = 16'b0000000000000000;
    assign weights1[54][146] = 16'b0000000000000000;
    assign weights1[54][147] = 16'b0000000000000000;
    assign weights1[54][148] = 16'b0000000000000000;
    assign weights1[54][149] = 16'b0000000000000000;
    assign weights1[54][150] = 16'b0000000000000000;
    assign weights1[54][151] = 16'b0000000000000000;
    assign weights1[54][152] = 16'b0000000000000000;
    assign weights1[54][153] = 16'b0000000000000000;
    assign weights1[54][154] = 16'b0000000000000000;
    assign weights1[54][155] = 16'b0000000000000000;
    assign weights1[54][156] = 16'b0000000000000000;
    assign weights1[54][157] = 16'b0000000000000000;
    assign weights1[54][158] = 16'b0000000000000000;
    assign weights1[54][159] = 16'b0000000000000000;
    assign weights1[54][160] = 16'b0000000000000000;
    assign weights1[54][161] = 16'b0000000000000000;
    assign weights1[54][162] = 16'b0000000000000000;
    assign weights1[54][163] = 16'b0000000000000000;
    assign weights1[54][164] = 16'b0000000000000000;
    assign weights1[54][165] = 16'b0000000000000000;
    assign weights1[54][166] = 16'b0000000000000000;
    assign weights1[54][167] = 16'b0000000000000000;
    assign weights1[54][168] = 16'b0000000000000000;
    assign weights1[54][169] = 16'b0000000000000000;
    assign weights1[54][170] = 16'b0000000000000000;
    assign weights1[54][171] = 16'b0000000000000000;
    assign weights1[54][172] = 16'b0000000000000000;
    assign weights1[54][173] = 16'b0000000000000000;
    assign weights1[54][174] = 16'b0000000000000000;
    assign weights1[54][175] = 16'b0000000000000000;
    assign weights1[54][176] = 16'b0000000000000000;
    assign weights1[54][177] = 16'b0000000000000000;
    assign weights1[54][178] = 16'b0000000000000000;
    assign weights1[54][179] = 16'b0000000000000000;
    assign weights1[54][180] = 16'b0000000000000000;
    assign weights1[54][181] = 16'b0000000000000000;
    assign weights1[54][182] = 16'b0000000000000000;
    assign weights1[54][183] = 16'b0000000000000000;
    assign weights1[54][184] = 16'b0000000000000000;
    assign weights1[54][185] = 16'b0000000000000000;
    assign weights1[54][186] = 16'b0000000000000000;
    assign weights1[54][187] = 16'b0000000000000000;
    assign weights1[54][188] = 16'b0000000000000000;
    assign weights1[54][189] = 16'b0000000000000000;
    assign weights1[54][190] = 16'b0000000000000000;
    assign weights1[54][191] = 16'b0000000000000000;
    assign weights1[54][192] = 16'b0000000000000000;
    assign weights1[54][193] = 16'b0000000000000000;
    assign weights1[54][194] = 16'b0000000000000000;
    assign weights1[54][195] = 16'b0000000000000000;
    assign weights1[54][196] = 16'b0000000000000000;
    assign weights1[54][197] = 16'b0000000000000000;
    assign weights1[54][198] = 16'b0000000000000000;
    assign weights1[54][199] = 16'b0000000000000000;
    assign weights1[54][200] = 16'b0000000000000000;
    assign weights1[54][201] = 16'b0000000000000000;
    assign weights1[54][202] = 16'b0000000000000000;
    assign weights1[54][203] = 16'b0000000000000000;
    assign weights1[54][204] = 16'b0000000000000000;
    assign weights1[54][205] = 16'b0000000000000000;
    assign weights1[54][206] = 16'b0000000000000000;
    assign weights1[54][207] = 16'b0000000000000000;
    assign weights1[54][208] = 16'b0000000000000000;
    assign weights1[54][209] = 16'b0000000000000000;
    assign weights1[54][210] = 16'b0000000000000000;
    assign weights1[54][211] = 16'b0000000000000000;
    assign weights1[54][212] = 16'b0000000000000000;
    assign weights1[54][213] = 16'b0000000000000000;
    assign weights1[54][214] = 16'b0000000000000000;
    assign weights1[54][215] = 16'b0000000000000000;
    assign weights1[54][216] = 16'b0000000000000000;
    assign weights1[54][217] = 16'b0000000000000000;
    assign weights1[54][218] = 16'b0000000000000000;
    assign weights1[54][219] = 16'b0000000000000000;
    assign weights1[54][220] = 16'b0000000000000000;
    assign weights1[54][221] = 16'b0000000000000000;
    assign weights1[54][222] = 16'b0000000000000000;
    assign weights1[54][223] = 16'b0000000000000000;
    assign weights1[54][224] = 16'b0000000000000000;
    assign weights1[54][225] = 16'b0000000000000000;
    assign weights1[54][226] = 16'b0000000000000000;
    assign weights1[54][227] = 16'b0000000000000000;
    assign weights1[54][228] = 16'b0000000000000000;
    assign weights1[54][229] = 16'b0000000000000000;
    assign weights1[54][230] = 16'b0000000000000000;
    assign weights1[54][231] = 16'b0000000000000000;
    assign weights1[54][232] = 16'b0000000000000000;
    assign weights1[54][233] = 16'b0000000000000000;
    assign weights1[54][234] = 16'b0000000000000000;
    assign weights1[54][235] = 16'b0000000000000000;
    assign weights1[54][236] = 16'b0000000000000000;
    assign weights1[54][237] = 16'b0000000000000000;
    assign weights1[54][238] = 16'b0000000000000000;
    assign weights1[54][239] = 16'b0000000000000000;
    assign weights1[54][240] = 16'b0000000000000000;
    assign weights1[54][241] = 16'b0000000000000000;
    assign weights1[54][242] = 16'b0000000000000000;
    assign weights1[54][243] = 16'b0000000000000000;
    assign weights1[54][244] = 16'b0000000000000000;
    assign weights1[54][245] = 16'b0000000000000000;
    assign weights1[54][246] = 16'b0000000000000000;
    assign weights1[54][247] = 16'b0000000000000000;
    assign weights1[54][248] = 16'b0000000000000000;
    assign weights1[54][249] = 16'b0000000000000000;
    assign weights1[54][250] = 16'b0000000000000000;
    assign weights1[54][251] = 16'b0000000000000000;
    assign weights1[54][252] = 16'b0000000000000000;
    assign weights1[54][253] = 16'b0000000000000000;
    assign weights1[54][254] = 16'b0000000000000000;
    assign weights1[54][255] = 16'b0000000000000000;
    assign weights1[54][256] = 16'b0000000000000000;
    assign weights1[54][257] = 16'b0000000000000000;
    assign weights1[54][258] = 16'b0000000000000000;
    assign weights1[54][259] = 16'b0000000000000000;
    assign weights1[54][260] = 16'b0000000000000000;
    assign weights1[54][261] = 16'b0000000000000000;
    assign weights1[54][262] = 16'b0000000000000000;
    assign weights1[54][263] = 16'b0000000000000000;
    assign weights1[54][264] = 16'b0000000000000000;
    assign weights1[54][265] = 16'b0000000000000000;
    assign weights1[54][266] = 16'b0000000000000000;
    assign weights1[54][267] = 16'b0000000000000000;
    assign weights1[54][268] = 16'b0000000000000000;
    assign weights1[54][269] = 16'b0000000000000000;
    assign weights1[54][270] = 16'b0000000000000000;
    assign weights1[54][271] = 16'b0000000000000000;
    assign weights1[54][272] = 16'b0000000000000000;
    assign weights1[54][273] = 16'b0000000000000000;
    assign weights1[54][274] = 16'b0000000000000000;
    assign weights1[54][275] = 16'b0000000000000000;
    assign weights1[54][276] = 16'b0000000000000000;
    assign weights1[54][277] = 16'b0000000000000000;
    assign weights1[54][278] = 16'b0000000000000000;
    assign weights1[54][279] = 16'b0000000000000000;
    assign weights1[54][280] = 16'b0000000000000000;
    assign weights1[54][281] = 16'b0000000000000000;
    assign weights1[54][282] = 16'b0000000000000000;
    assign weights1[54][283] = 16'b0000000000000000;
    assign weights1[54][284] = 16'b0000000000000000;
    assign weights1[54][285] = 16'b0000000000000000;
    assign weights1[54][286] = 16'b0000000000000000;
    assign weights1[54][287] = 16'b0000000000000000;
    assign weights1[54][288] = 16'b0000000000000000;
    assign weights1[54][289] = 16'b0000000000000000;
    assign weights1[54][290] = 16'b0000000000000000;
    assign weights1[54][291] = 16'b0000000000000000;
    assign weights1[54][292] = 16'b0000000000000000;
    assign weights1[54][293] = 16'b0000000000000000;
    assign weights1[54][294] = 16'b0000000000000000;
    assign weights1[54][295] = 16'b0000000000000000;
    assign weights1[54][296] = 16'b0000000000000000;
    assign weights1[54][297] = 16'b0000000000000000;
    assign weights1[54][298] = 16'b0000000000000000;
    assign weights1[54][299] = 16'b0000000000000000;
    assign weights1[54][300] = 16'b0000000000000000;
    assign weights1[54][301] = 16'b0000000000000000;
    assign weights1[54][302] = 16'b0000000000000000;
    assign weights1[54][303] = 16'b0000000000000000;
    assign weights1[54][304] = 16'b0000000000000000;
    assign weights1[54][305] = 16'b0000000000000000;
    assign weights1[54][306] = 16'b0000000000000000;
    assign weights1[54][307] = 16'b0000000000000000;
    assign weights1[54][308] = 16'b0000000000000000;
    assign weights1[54][309] = 16'b0000000000000000;
    assign weights1[54][310] = 16'b0000000000000000;
    assign weights1[54][311] = 16'b0000000000000000;
    assign weights1[54][312] = 16'b0000000000000000;
    assign weights1[54][313] = 16'b0000000000000000;
    assign weights1[54][314] = 16'b0000000000000000;
    assign weights1[54][315] = 16'b0000000000000000;
    assign weights1[54][316] = 16'b0000000000000000;
    assign weights1[54][317] = 16'b0000000000000000;
    assign weights1[54][318] = 16'b0000000000000000;
    assign weights1[54][319] = 16'b0000000000000000;
    assign weights1[54][320] = 16'b0000000000000000;
    assign weights1[54][321] = 16'b0000000000000000;
    assign weights1[54][322] = 16'b0000000000000000;
    assign weights1[54][323] = 16'b0000000000000000;
    assign weights1[54][324] = 16'b0000000000000000;
    assign weights1[54][325] = 16'b0000000000000000;
    assign weights1[54][326] = 16'b0000000000000000;
    assign weights1[54][327] = 16'b0000000000000000;
    assign weights1[54][328] = 16'b0000000000000000;
    assign weights1[54][329] = 16'b0000000000000000;
    assign weights1[54][330] = 16'b0000000000000000;
    assign weights1[54][331] = 16'b0000000000000000;
    assign weights1[54][332] = 16'b0000000000000000;
    assign weights1[54][333] = 16'b0000000000000000;
    assign weights1[54][334] = 16'b0000000000000000;
    assign weights1[54][335] = 16'b0000000000000000;
    assign weights1[54][336] = 16'b0000000000000000;
    assign weights1[54][337] = 16'b0000000000000000;
    assign weights1[54][338] = 16'b0000000000000000;
    assign weights1[54][339] = 16'b0000000000000000;
    assign weights1[54][340] = 16'b0000000000000000;
    assign weights1[54][341] = 16'b0000000000000000;
    assign weights1[54][342] = 16'b0000000000000000;
    assign weights1[54][343] = 16'b0000000000000000;
    assign weights1[54][344] = 16'b0000000000000000;
    assign weights1[54][345] = 16'b0000000000000000;
    assign weights1[54][346] = 16'b0000000000000000;
    assign weights1[54][347] = 16'b0000000000000000;
    assign weights1[54][348] = 16'b0000000000000000;
    assign weights1[54][349] = 16'b0000000000000000;
    assign weights1[54][350] = 16'b0000000000000000;
    assign weights1[54][351] = 16'b0000000000000000;
    assign weights1[54][352] = 16'b0000000000000000;
    assign weights1[54][353] = 16'b0000000000000000;
    assign weights1[54][354] = 16'b0000000000000000;
    assign weights1[54][355] = 16'b0000000000000000;
    assign weights1[54][356] = 16'b0000000000000000;
    assign weights1[54][357] = 16'b0000000000000000;
    assign weights1[54][358] = 16'b0000000000000000;
    assign weights1[54][359] = 16'b0000000000000000;
    assign weights1[54][360] = 16'b0000000000000000;
    assign weights1[54][361] = 16'b0000000000000000;
    assign weights1[54][362] = 16'b0000000000000000;
    assign weights1[54][363] = 16'b0000000000000000;
    assign weights1[54][364] = 16'b0000000000000000;
    assign weights1[54][365] = 16'b0000000000000000;
    assign weights1[54][366] = 16'b0000000000000000;
    assign weights1[54][367] = 16'b0000000000000000;
    assign weights1[54][368] = 16'b0000000000000000;
    assign weights1[54][369] = 16'b0000000000000000;
    assign weights1[54][370] = 16'b0000000000000000;
    assign weights1[54][371] = 16'b0000000000000000;
    assign weights1[54][372] = 16'b0000000000000000;
    assign weights1[54][373] = 16'b0000000000000000;
    assign weights1[54][374] = 16'b0000000000000000;
    assign weights1[54][375] = 16'b0000000000000000;
    assign weights1[54][376] = 16'b0000000000000000;
    assign weights1[54][377] = 16'b0000000000000000;
    assign weights1[54][378] = 16'b0000000000000000;
    assign weights1[54][379] = 16'b0000000000000000;
    assign weights1[54][380] = 16'b0000000000000000;
    assign weights1[54][381] = 16'b0000000000000000;
    assign weights1[54][382] = 16'b0000000000000000;
    assign weights1[54][383] = 16'b0000000000000000;
    assign weights1[54][384] = 16'b0000000000000000;
    assign weights1[54][385] = 16'b0000000000000000;
    assign weights1[54][386] = 16'b0000000000000000;
    assign weights1[54][387] = 16'b0000000000000000;
    assign weights1[54][388] = 16'b0000000000000000;
    assign weights1[54][389] = 16'b0000000000000000;
    assign weights1[54][390] = 16'b0000000000000000;
    assign weights1[54][391] = 16'b0000000000000000;
    assign weights1[54][392] = 16'b0000000000000000;
    assign weights1[54][393] = 16'b0000000000000000;
    assign weights1[54][394] = 16'b0000000000000000;
    assign weights1[54][395] = 16'b0000000000000000;
    assign weights1[54][396] = 16'b0000000000000000;
    assign weights1[54][397] = 16'b0000000000000000;
    assign weights1[54][398] = 16'b0000000000000000;
    assign weights1[54][399] = 16'b0000000000000000;
    assign weights1[54][400] = 16'b0000000000000000;
    assign weights1[54][401] = 16'b0000000000000000;
    assign weights1[54][402] = 16'b0000000000000000;
    assign weights1[54][403] = 16'b0000000000000000;
    assign weights1[54][404] = 16'b0000000000000000;
    assign weights1[54][405] = 16'b0000000000000000;
    assign weights1[54][406] = 16'b0000000000000000;
    assign weights1[54][407] = 16'b0000000000000000;
    assign weights1[54][408] = 16'b0000000000000000;
    assign weights1[54][409] = 16'b0000000000000000;
    assign weights1[54][410] = 16'b0000000000000000;
    assign weights1[54][411] = 16'b0000000000000000;
    assign weights1[54][412] = 16'b0000000000000000;
    assign weights1[54][413] = 16'b0000000000000000;
    assign weights1[54][414] = 16'b0000000000000000;
    assign weights1[54][415] = 16'b0000000000000000;
    assign weights1[54][416] = 16'b0000000000000000;
    assign weights1[54][417] = 16'b0000000000000000;
    assign weights1[54][418] = 16'b0000000000000000;
    assign weights1[54][419] = 16'b0000000000000000;
    assign weights1[54][420] = 16'b0000000000000000;
    assign weights1[54][421] = 16'b0000000000000000;
    assign weights1[54][422] = 16'b0000000000000000;
    assign weights1[54][423] = 16'b0000000000000000;
    assign weights1[54][424] = 16'b0000000000000000;
    assign weights1[54][425] = 16'b0000000000000000;
    assign weights1[54][426] = 16'b0000000000000000;
    assign weights1[54][427] = 16'b0000000000000000;
    assign weights1[54][428] = 16'b0000000000000000;
    assign weights1[54][429] = 16'b0000000000000000;
    assign weights1[54][430] = 16'b0000000000000000;
    assign weights1[54][431] = 16'b0000000000000000;
    assign weights1[54][432] = 16'b0000000000000000;
    assign weights1[54][433] = 16'b0000000000000000;
    assign weights1[54][434] = 16'b0000000000000000;
    assign weights1[54][435] = 16'b0000000000000000;
    assign weights1[54][436] = 16'b0000000000000000;
    assign weights1[54][437] = 16'b0000000000000000;
    assign weights1[54][438] = 16'b0000000000000000;
    assign weights1[54][439] = 16'b0000000000000000;
    assign weights1[54][440] = 16'b0000000000000000;
    assign weights1[54][441] = 16'b0000000000000000;
    assign weights1[54][442] = 16'b0000000000000000;
    assign weights1[54][443] = 16'b0000000000000000;
    assign weights1[54][444] = 16'b0000000000000000;
    assign weights1[54][445] = 16'b0000000000000000;
    assign weights1[54][446] = 16'b0000000000000000;
    assign weights1[54][447] = 16'b0000000000000000;
    assign weights1[54][448] = 16'b0000000000000000;
    assign weights1[54][449] = 16'b0000000000000000;
    assign weights1[54][450] = 16'b0000000000000000;
    assign weights1[54][451] = 16'b0000000000000000;
    assign weights1[54][452] = 16'b0000000000000000;
    assign weights1[54][453] = 16'b0000000000000000;
    assign weights1[54][454] = 16'b0000000000000000;
    assign weights1[54][455] = 16'b0000000000000000;
    assign weights1[54][456] = 16'b0000000000000000;
    assign weights1[54][457] = 16'b0000000000000000;
    assign weights1[54][458] = 16'b0000000000000000;
    assign weights1[54][459] = 16'b0000000000000000;
    assign weights1[54][460] = 16'b0000000000000000;
    assign weights1[54][461] = 16'b0000000000000000;
    assign weights1[54][462] = 16'b0000000000000000;
    assign weights1[54][463] = 16'b0000000000000000;
    assign weights1[54][464] = 16'b0000000000000000;
    assign weights1[54][465] = 16'b0000000000000000;
    assign weights1[54][466] = 16'b0000000000000000;
    assign weights1[54][467] = 16'b0000000000000000;
    assign weights1[54][468] = 16'b0000000000000000;
    assign weights1[54][469] = 16'b0000000000000000;
    assign weights1[54][470] = 16'b0000000000000000;
    assign weights1[54][471] = 16'b0000000000000000;
    assign weights1[54][472] = 16'b0000000000000000;
    assign weights1[54][473] = 16'b0000000000000000;
    assign weights1[54][474] = 16'b0000000000000000;
    assign weights1[54][475] = 16'b0000000000000000;
    assign weights1[54][476] = 16'b0000000000000000;
    assign weights1[54][477] = 16'b0000000000000000;
    assign weights1[54][478] = 16'b0000000000000000;
    assign weights1[54][479] = 16'b0000000000000000;
    assign weights1[54][480] = 16'b0000000000000000;
    assign weights1[54][481] = 16'b0000000000000000;
    assign weights1[54][482] = 16'b0000000000000000;
    assign weights1[54][483] = 16'b0000000000000000;
    assign weights1[54][484] = 16'b0000000000000000;
    assign weights1[54][485] = 16'b0000000000000000;
    assign weights1[54][486] = 16'b0000000000000000;
    assign weights1[54][487] = 16'b0000000000000000;
    assign weights1[54][488] = 16'b0000000000000000;
    assign weights1[54][489] = 16'b0000000000000000;
    assign weights1[54][490] = 16'b0000000000000000;
    assign weights1[54][491] = 16'b0000000000000000;
    assign weights1[54][492] = 16'b0000000000000000;
    assign weights1[54][493] = 16'b0000000000000000;
    assign weights1[54][494] = 16'b0000000000000000;
    assign weights1[54][495] = 16'b0000000000000000;
    assign weights1[54][496] = 16'b0000000000000000;
    assign weights1[54][497] = 16'b0000000000000000;
    assign weights1[54][498] = 16'b0000000000000000;
    assign weights1[54][499] = 16'b0000000000000000;
    assign weights1[54][500] = 16'b0000000000000000;
    assign weights1[54][501] = 16'b0000000000000000;
    assign weights1[54][502] = 16'b0000000000000000;
    assign weights1[54][503] = 16'b0000000000000000;
    assign weights1[54][504] = 16'b0000000000000000;
    assign weights1[54][505] = 16'b0000000000000000;
    assign weights1[54][506] = 16'b0000000000000000;
    assign weights1[54][507] = 16'b0000000000000000;
    assign weights1[54][508] = 16'b0000000000000000;
    assign weights1[54][509] = 16'b0000000000000000;
    assign weights1[54][510] = 16'b0000000000000000;
    assign weights1[54][511] = 16'b0000000000000000;
    assign weights1[54][512] = 16'b0000000000000000;
    assign weights1[54][513] = 16'b0000000000000000;
    assign weights1[54][514] = 16'b0000000000000000;
    assign weights1[54][515] = 16'b0000000000000000;
    assign weights1[54][516] = 16'b0000000000000000;
    assign weights1[54][517] = 16'b0000000000000000;
    assign weights1[54][518] = 16'b0000000000000000;
    assign weights1[54][519] = 16'b0000000000000000;
    assign weights1[54][520] = 16'b0000000000000000;
    assign weights1[54][521] = 16'b0000000000000000;
    assign weights1[54][522] = 16'b0000000000000000;
    assign weights1[54][523] = 16'b0000000000000000;
    assign weights1[54][524] = 16'b0000000000000000;
    assign weights1[54][525] = 16'b0000000000000000;
    assign weights1[54][526] = 16'b0000000000000000;
    assign weights1[54][527] = 16'b0000000000000000;
    assign weights1[54][528] = 16'b0000000000000000;
    assign weights1[54][529] = 16'b0000000000000000;
    assign weights1[54][530] = 16'b0000000000000000;
    assign weights1[54][531] = 16'b0000000000000000;
    assign weights1[54][532] = 16'b0000000000000000;
    assign weights1[54][533] = 16'b0000000000000000;
    assign weights1[54][534] = 16'b0000000000000000;
    assign weights1[54][535] = 16'b0000000000000000;
    assign weights1[54][536] = 16'b0000000000000000;
    assign weights1[54][537] = 16'b0000000000000000;
    assign weights1[54][538] = 16'b0000000000000000;
    assign weights1[54][539] = 16'b0000000000000000;
    assign weights1[54][540] = 16'b0000000000000000;
    assign weights1[54][541] = 16'b0000000000000000;
    assign weights1[54][542] = 16'b0000000000000000;
    assign weights1[54][543] = 16'b0000000000000000;
    assign weights1[54][544] = 16'b0000000000000000;
    assign weights1[54][545] = 16'b0000000000000000;
    assign weights1[54][546] = 16'b0000000000000000;
    assign weights1[54][547] = 16'b0000000000000000;
    assign weights1[54][548] = 16'b0000000000000000;
    assign weights1[54][549] = 16'b0000000000000000;
    assign weights1[54][550] = 16'b0000000000000000;
    assign weights1[54][551] = 16'b0000000000000000;
    assign weights1[54][552] = 16'b0000000000000000;
    assign weights1[54][553] = 16'b0000000000000000;
    assign weights1[54][554] = 16'b0000000000000000;
    assign weights1[54][555] = 16'b0000000000000000;
    assign weights1[54][556] = 16'b0000000000000000;
    assign weights1[54][557] = 16'b0000000000000000;
    assign weights1[54][558] = 16'b0000000000000000;
    assign weights1[54][559] = 16'b0000000000000000;
    assign weights1[54][560] = 16'b0000000000000000;
    assign weights1[54][561] = 16'b0000000000000000;
    assign weights1[54][562] = 16'b0000000000000000;
    assign weights1[54][563] = 16'b0000000000000000;
    assign weights1[54][564] = 16'b0000000000000000;
    assign weights1[54][565] = 16'b0000000000000000;
    assign weights1[54][566] = 16'b0000000000000000;
    assign weights1[54][567] = 16'b0000000000000000;
    assign weights1[54][568] = 16'b0000000000000000;
    assign weights1[54][569] = 16'b0000000000000000;
    assign weights1[54][570] = 16'b0000000000000000;
    assign weights1[54][571] = 16'b0000000000000000;
    assign weights1[54][572] = 16'b0000000000000000;
    assign weights1[54][573] = 16'b0000000000000000;
    assign weights1[54][574] = 16'b0000000000000000;
    assign weights1[54][575] = 16'b0000000000000000;
    assign weights1[54][576] = 16'b0000000000000000;
    assign weights1[54][577] = 16'b0000000000000000;
    assign weights1[54][578] = 16'b0000000000000000;
    assign weights1[54][579] = 16'b0000000000000000;
    assign weights1[54][580] = 16'b0000000000000000;
    assign weights1[54][581] = 16'b0000000000000000;
    assign weights1[54][582] = 16'b0000000000000000;
    assign weights1[54][583] = 16'b0000000000000000;
    assign weights1[54][584] = 16'b0000000000000000;
    assign weights1[54][585] = 16'b0000000000000000;
    assign weights1[54][586] = 16'b0000000000000000;
    assign weights1[54][587] = 16'b0000000000000000;
    assign weights1[54][588] = 16'b0000000000000000;
    assign weights1[54][589] = 16'b0000000000000000;
    assign weights1[54][590] = 16'b0000000000000000;
    assign weights1[54][591] = 16'b0000000000000000;
    assign weights1[54][592] = 16'b0000000000000000;
    assign weights1[54][593] = 16'b0000000000000000;
    assign weights1[54][594] = 16'b0000000000000000;
    assign weights1[54][595] = 16'b0000000000000000;
    assign weights1[54][596] = 16'b0000000000000000;
    assign weights1[54][597] = 16'b0000000000000000;
    assign weights1[54][598] = 16'b0000000000000000;
    assign weights1[54][599] = 16'b0000000000000000;
    assign weights1[54][600] = 16'b0000000000000000;
    assign weights1[54][601] = 16'b0000000000000000;
    assign weights1[54][602] = 16'b0000000000000000;
    assign weights1[54][603] = 16'b0000000000000000;
    assign weights1[54][604] = 16'b0000000000000000;
    assign weights1[54][605] = 16'b0000000000000000;
    assign weights1[54][606] = 16'b0000000000000000;
    assign weights1[54][607] = 16'b0000000000000000;
    assign weights1[54][608] = 16'b0000000000000000;
    assign weights1[54][609] = 16'b0000000000000000;
    assign weights1[54][610] = 16'b0000000000000000;
    assign weights1[54][611] = 16'b0000000000000000;
    assign weights1[54][612] = 16'b0000000000000000;
    assign weights1[54][613] = 16'b0000000000000000;
    assign weights1[54][614] = 16'b0000000000000000;
    assign weights1[54][615] = 16'b0000000000000000;
    assign weights1[54][616] = 16'b0000000000000000;
    assign weights1[54][617] = 16'b0000000000000000;
    assign weights1[54][618] = 16'b0000000000000000;
    assign weights1[54][619] = 16'b0000000000000000;
    assign weights1[54][620] = 16'b0000000000000000;
    assign weights1[54][621] = 16'b0000000000000000;
    assign weights1[54][622] = 16'b0000000000000000;
    assign weights1[54][623] = 16'b0000000000000000;
    assign weights1[54][624] = 16'b0000000000000000;
    assign weights1[54][625] = 16'b0000000000000000;
    assign weights1[54][626] = 16'b0000000000000000;
    assign weights1[54][627] = 16'b0000000000000000;
    assign weights1[54][628] = 16'b0000000000000000;
    assign weights1[54][629] = 16'b0000000000000000;
    assign weights1[54][630] = 16'b0000000000000000;
    assign weights1[54][631] = 16'b0000000000000000;
    assign weights1[54][632] = 16'b0000000000000000;
    assign weights1[54][633] = 16'b0000000000000000;
    assign weights1[54][634] = 16'b0000000000000000;
    assign weights1[54][635] = 16'b0000000000000000;
    assign weights1[54][636] = 16'b0000000000000000;
    assign weights1[54][637] = 16'b0000000000000000;
    assign weights1[54][638] = 16'b0000000000000000;
    assign weights1[54][639] = 16'b0000000000000000;
    assign weights1[54][640] = 16'b0000000000000000;
    assign weights1[54][641] = 16'b0000000000000000;
    assign weights1[54][642] = 16'b0000000000000000;
    assign weights1[54][643] = 16'b0000000000000000;
    assign weights1[54][644] = 16'b0000000000000000;
    assign weights1[54][645] = 16'b0000000000000000;
    assign weights1[54][646] = 16'b0000000000000000;
    assign weights1[54][647] = 16'b0000000000000000;
    assign weights1[54][648] = 16'b0000000000000000;
    assign weights1[54][649] = 16'b0000000000000000;
    assign weights1[54][650] = 16'b0000000000000000;
    assign weights1[54][651] = 16'b0000000000000000;
    assign weights1[54][652] = 16'b0000000000000000;
    assign weights1[54][653] = 16'b0000000000000000;
    assign weights1[54][654] = 16'b0000000000000000;
    assign weights1[54][655] = 16'b0000000000000000;
    assign weights1[54][656] = 16'b0000000000000000;
    assign weights1[54][657] = 16'b0000000000000000;
    assign weights1[54][658] = 16'b0000000000000000;
    assign weights1[54][659] = 16'b0000000000000000;
    assign weights1[54][660] = 16'b0000000000000000;
    assign weights1[54][661] = 16'b0000000000000000;
    assign weights1[54][662] = 16'b0000000000000000;
    assign weights1[54][663] = 16'b0000000000000000;
    assign weights1[54][664] = 16'b0000000000000000;
    assign weights1[54][665] = 16'b0000000000000000;
    assign weights1[54][666] = 16'b0000000000000000;
    assign weights1[54][667] = 16'b0000000000000000;
    assign weights1[54][668] = 16'b0000000000000000;
    assign weights1[54][669] = 16'b0000000000000000;
    assign weights1[54][670] = 16'b0000000000000000;
    assign weights1[54][671] = 16'b0000000000000000;
    assign weights1[54][672] = 16'b0000000000000000;
    assign weights1[54][673] = 16'b0000000000000000;
    assign weights1[54][674] = 16'b0000000000000000;
    assign weights1[54][675] = 16'b0000000000000000;
    assign weights1[54][676] = 16'b0000000000000000;
    assign weights1[54][677] = 16'b0000000000000000;
    assign weights1[54][678] = 16'b0000000000000000;
    assign weights1[54][679] = 16'b0000000000000000;
    assign weights1[54][680] = 16'b0000000000000000;
    assign weights1[54][681] = 16'b0000000000000000;
    assign weights1[54][682] = 16'b0000000000000000;
    assign weights1[54][683] = 16'b0000000000000000;
    assign weights1[54][684] = 16'b0000000000000000;
    assign weights1[54][685] = 16'b0000000000000000;
    assign weights1[54][686] = 16'b0000000000000000;
    assign weights1[54][687] = 16'b0000000000000000;
    assign weights1[54][688] = 16'b0000000000000000;
    assign weights1[54][689] = 16'b0000000000000000;
    assign weights1[54][690] = 16'b0000000000000000;
    assign weights1[54][691] = 16'b0000000000000000;
    assign weights1[54][692] = 16'b0000000000000000;
    assign weights1[54][693] = 16'b0000000000000000;
    assign weights1[54][694] = 16'b0000000000000000;
    assign weights1[54][695] = 16'b0000000000000000;
    assign weights1[54][696] = 16'b0000000000000000;
    assign weights1[54][697] = 16'b0000000000000000;
    assign weights1[54][698] = 16'b0000000000000000;
    assign weights1[54][699] = 16'b0000000000000000;
    assign weights1[54][700] = 16'b0000000000000000;
    assign weights1[54][701] = 16'b0000000000000000;
    assign weights1[54][702] = 16'b0000000000000000;
    assign weights1[54][703] = 16'b0000000000000000;
    assign weights1[54][704] = 16'b0000000000000000;
    assign weights1[54][705] = 16'b0000000000000000;
    assign weights1[54][706] = 16'b0000000000000000;
    assign weights1[54][707] = 16'b0000000000000000;
    assign weights1[54][708] = 16'b0000000000000000;
    assign weights1[54][709] = 16'b0000000000000000;
    assign weights1[54][710] = 16'b0000000000000000;
    assign weights1[54][711] = 16'b0000000000000000;
    assign weights1[54][712] = 16'b0000000000000000;
    assign weights1[54][713] = 16'b0000000000000000;
    assign weights1[54][714] = 16'b0000000000000000;
    assign weights1[54][715] = 16'b0000000000000000;
    assign weights1[54][716] = 16'b0000000000000000;
    assign weights1[54][717] = 16'b0000000000000000;
    assign weights1[54][718] = 16'b0000000000000000;
    assign weights1[54][719] = 16'b0000000000000000;
    assign weights1[54][720] = 16'b0000000000000000;
    assign weights1[54][721] = 16'b0000000000000000;
    assign weights1[54][722] = 16'b0000000000000000;
    assign weights1[54][723] = 16'b0000000000000000;
    assign weights1[54][724] = 16'b0000000000000000;
    assign weights1[54][725] = 16'b0000000000000000;
    assign weights1[54][726] = 16'b0000000000000000;
    assign weights1[54][727] = 16'b0000000000000000;
    assign weights1[54][728] = 16'b0000000000000000;
    assign weights1[54][729] = 16'b0000000000000000;
    assign weights1[54][730] = 16'b0000000000000000;
    assign weights1[54][731] = 16'b0000000000000000;
    assign weights1[54][732] = 16'b0000000000000000;
    assign weights1[54][733] = 16'b0000000000000000;
    assign weights1[54][734] = 16'b0000000000000000;
    assign weights1[54][735] = 16'b0000000000000000;
    assign weights1[54][736] = 16'b0000000000000000;
    assign weights1[54][737] = 16'b0000000000000000;
    assign weights1[54][738] = 16'b0000000000000000;
    assign weights1[54][739] = 16'b0000000000000000;
    assign weights1[54][740] = 16'b0000000000000000;
    assign weights1[54][741] = 16'b0000000000000000;
    assign weights1[54][742] = 16'b0000000000000000;
    assign weights1[54][743] = 16'b0000000000000000;
    assign weights1[54][744] = 16'b0000000000000000;
    assign weights1[54][745] = 16'b0000000000000000;
    assign weights1[54][746] = 16'b0000000000000000;
    assign weights1[54][747] = 16'b0000000000000000;
    assign weights1[54][748] = 16'b0000000000000000;
    assign weights1[54][749] = 16'b0000000000000000;
    assign weights1[54][750] = 16'b0000000000000000;
    assign weights1[54][751] = 16'b0000000000000000;
    assign weights1[54][752] = 16'b0000000000000000;
    assign weights1[54][753] = 16'b0000000000000000;
    assign weights1[54][754] = 16'b0000000000000000;
    assign weights1[54][755] = 16'b0000000000000000;
    assign weights1[54][756] = 16'b0000000000000000;
    assign weights1[54][757] = 16'b0000000000000000;
    assign weights1[54][758] = 16'b0000000000000000;
    assign weights1[54][759] = 16'b0000000000000000;
    assign weights1[54][760] = 16'b0000000000000000;
    assign weights1[54][761] = 16'b0000000000000000;
    assign weights1[54][762] = 16'b0000000000000000;
    assign weights1[54][763] = 16'b0000000000000000;
    assign weights1[54][764] = 16'b0000000000000000;
    assign weights1[54][765] = 16'b0000000000000000;
    assign weights1[54][766] = 16'b0000000000000000;
    assign weights1[54][767] = 16'b0000000000000000;
    assign weights1[54][768] = 16'b0000000000000000;
    assign weights1[54][769] = 16'b0000000000000000;
    assign weights1[54][770] = 16'b0000000000000000;
    assign weights1[54][771] = 16'b0000000000000000;
    assign weights1[54][772] = 16'b0000000000000000;
    assign weights1[54][773] = 16'b0000000000000000;
    assign weights1[54][774] = 16'b0000000000000000;
    assign weights1[54][775] = 16'b0000000000000000;
    assign weights1[54][776] = 16'b0000000000000000;
    assign weights1[54][777] = 16'b0000000000000000;
    assign weights1[54][778] = 16'b0000000000000000;
    assign weights1[54][779] = 16'b0000000000000000;
    assign weights1[54][780] = 16'b0000000000000000;
    assign weights1[54][781] = 16'b0000000000000000;
    assign weights1[54][782] = 16'b0000000000000000;
    assign weights1[54][783] = 16'b0000000000000000;
    assign weights1[55][0] = 16'b0000000000000000;
    assign weights1[55][1] = 16'b1111111111111111;
    assign weights1[55][2] = 16'b1111111111111111;
    assign weights1[55][3] = 16'b0000000000000000;
    assign weights1[55][4] = 16'b0000000000000000;
    assign weights1[55][5] = 16'b0000000000000000;
    assign weights1[55][6] = 16'b0000000000000000;
    assign weights1[55][7] = 16'b1111111111111111;
    assign weights1[55][8] = 16'b1111111111111111;
    assign weights1[55][9] = 16'b1111111111111110;
    assign weights1[55][10] = 16'b0000000000000001;
    assign weights1[55][11] = 16'b1111111111111010;
    assign weights1[55][12] = 16'b1111111111111010;
    assign weights1[55][13] = 16'b1111111111111101;
    assign weights1[55][14] = 16'b1111111111111110;
    assign weights1[55][15] = 16'b1111111111111100;
    assign weights1[55][16] = 16'b1111111111110110;
    assign weights1[55][17] = 16'b1111111111110100;
    assign weights1[55][18] = 16'b1111111111110110;
    assign weights1[55][19] = 16'b1111111111110110;
    assign weights1[55][20] = 16'b1111111111110101;
    assign weights1[55][21] = 16'b1111111111111000;
    assign weights1[55][22] = 16'b1111111111111010;
    assign weights1[55][23] = 16'b1111111111111100;
    assign weights1[55][24] = 16'b1111111111111101;
    assign weights1[55][25] = 16'b1111111111111111;
    assign weights1[55][26] = 16'b0000000000000000;
    assign weights1[55][27] = 16'b0000000000000000;
    assign weights1[55][28] = 16'b0000000000000000;
    assign weights1[55][29] = 16'b1111111111111110;
    assign weights1[55][30] = 16'b1111111111111110;
    assign weights1[55][31] = 16'b1111111111111111;
    assign weights1[55][32] = 16'b0000000000000000;
    assign weights1[55][33] = 16'b0000000000000100;
    assign weights1[55][34] = 16'b0000000000000101;
    assign weights1[55][35] = 16'b0000000000000010;
    assign weights1[55][36] = 16'b1111111111111100;
    assign weights1[55][37] = 16'b1111111111110111;
    assign weights1[55][38] = 16'b1111111111111011;
    assign weights1[55][39] = 16'b1111111111111011;
    assign weights1[55][40] = 16'b1111111111111010;
    assign weights1[55][41] = 16'b1111111111101111;
    assign weights1[55][42] = 16'b1111111111101110;
    assign weights1[55][43] = 16'b1111111111101100;
    assign weights1[55][44] = 16'b1111111111101111;
    assign weights1[55][45] = 16'b1111111111100111;
    assign weights1[55][46] = 16'b1111111111101001;
    assign weights1[55][47] = 16'b1111111111101110;
    assign weights1[55][48] = 16'b1111111111110001;
    assign weights1[55][49] = 16'b1111111111110101;
    assign weights1[55][50] = 16'b1111111111111000;
    assign weights1[55][51] = 16'b1111111111111001;
    assign weights1[55][52] = 16'b1111111111111100;
    assign weights1[55][53] = 16'b1111111111111111;
    assign weights1[55][54] = 16'b0000000000000001;
    assign weights1[55][55] = 16'b0000000000000000;
    assign weights1[55][56] = 16'b1111111111111111;
    assign weights1[55][57] = 16'b1111111111111111;
    assign weights1[55][58] = 16'b0000000000000001;
    assign weights1[55][59] = 16'b0000000000000000;
    assign weights1[55][60] = 16'b0000000000000010;
    assign weights1[55][61] = 16'b0000000000000100;
    assign weights1[55][62] = 16'b0000000000001011;
    assign weights1[55][63] = 16'b1111111111111110;
    assign weights1[55][64] = 16'b1111111111111001;
    assign weights1[55][65] = 16'b1111111111111000;
    assign weights1[55][66] = 16'b1111111111111010;
    assign weights1[55][67] = 16'b1111111111111000;
    assign weights1[55][68] = 16'b1111111111110001;
    assign weights1[55][69] = 16'b1111111111101011;
    assign weights1[55][70] = 16'b1111111111101100;
    assign weights1[55][71] = 16'b1111111111100100;
    assign weights1[55][72] = 16'b1111111111101010;
    assign weights1[55][73] = 16'b1111111111100110;
    assign weights1[55][74] = 16'b1111111111101100;
    assign weights1[55][75] = 16'b1111111111100101;
    assign weights1[55][76] = 16'b1111111111101001;
    assign weights1[55][77] = 16'b1111111111101001;
    assign weights1[55][78] = 16'b1111111111110001;
    assign weights1[55][79] = 16'b1111111111110111;
    assign weights1[55][80] = 16'b1111111111111111;
    assign weights1[55][81] = 16'b1111111111111111;
    assign weights1[55][82] = 16'b1111111111111110;
    assign weights1[55][83] = 16'b1111111111111110;
    assign weights1[55][84] = 16'b1111111111111111;
    assign weights1[55][85] = 16'b1111111111111110;
    assign weights1[55][86] = 16'b1111111111111111;
    assign weights1[55][87] = 16'b1111111111111110;
    assign weights1[55][88] = 16'b0000000000000000;
    assign weights1[55][89] = 16'b0000000000000010;
    assign weights1[55][90] = 16'b1111111111111111;
    assign weights1[55][91] = 16'b1111111111111110;
    assign weights1[55][92] = 16'b1111111111110100;
    assign weights1[55][93] = 16'b1111111111111110;
    assign weights1[55][94] = 16'b1111111111110101;
    assign weights1[55][95] = 16'b0000000000000010;
    assign weights1[55][96] = 16'b1111111111111100;
    assign weights1[55][97] = 16'b0000000000000110;
    assign weights1[55][98] = 16'b1111111111111101;
    assign weights1[55][99] = 16'b1111111111110001;
    assign weights1[55][100] = 16'b1111111111100011;
    assign weights1[55][101] = 16'b1111111111100011;
    assign weights1[55][102] = 16'b1111111111011100;
    assign weights1[55][103] = 16'b1111111111010111;
    assign weights1[55][104] = 16'b1111111111011110;
    assign weights1[55][105] = 16'b1111111111100011;
    assign weights1[55][106] = 16'b1111111111100101;
    assign weights1[55][107] = 16'b1111111111110110;
    assign weights1[55][108] = 16'b1111111111111000;
    assign weights1[55][109] = 16'b1111111111111011;
    assign weights1[55][110] = 16'b1111111111111000;
    assign weights1[55][111] = 16'b1111111111111010;
    assign weights1[55][112] = 16'b1111111111111111;
    assign weights1[55][113] = 16'b1111111111111110;
    assign weights1[55][114] = 16'b1111111111111110;
    assign weights1[55][115] = 16'b0000000000000001;
    assign weights1[55][116] = 16'b1111111111111100;
    assign weights1[55][117] = 16'b1111111111111100;
    assign weights1[55][118] = 16'b1111111111110111;
    assign weights1[55][119] = 16'b1111111111111000;
    assign weights1[55][120] = 16'b1111111111111000;
    assign weights1[55][121] = 16'b1111111111100011;
    assign weights1[55][122] = 16'b1111111111101000;
    assign weights1[55][123] = 16'b1111111111100100;
    assign weights1[55][124] = 16'b1111111111100010;
    assign weights1[55][125] = 16'b0000000000000001;
    assign weights1[55][126] = 16'b0000000000010001;
    assign weights1[55][127] = 16'b1111111111101010;
    assign weights1[55][128] = 16'b1111111111100000;
    assign weights1[55][129] = 16'b1111111111110011;
    assign weights1[55][130] = 16'b1111111111110100;
    assign weights1[55][131] = 16'b1111111111110000;
    assign weights1[55][132] = 16'b1111111111110010;
    assign weights1[55][133] = 16'b1111111111011110;
    assign weights1[55][134] = 16'b1111111111100101;
    assign weights1[55][135] = 16'b1111111111101001;
    assign weights1[55][136] = 16'b1111111111101101;
    assign weights1[55][137] = 16'b1111111111110010;
    assign weights1[55][138] = 16'b1111111111110100;
    assign weights1[55][139] = 16'b1111111111111100;
    assign weights1[55][140] = 16'b1111111111111111;
    assign weights1[55][141] = 16'b0000000000000001;
    assign weights1[55][142] = 16'b1111111111111010;
    assign weights1[55][143] = 16'b1111111111111010;
    assign weights1[55][144] = 16'b1111111111111100;
    assign weights1[55][145] = 16'b1111111111100101;
    assign weights1[55][146] = 16'b1111111111111000;
    assign weights1[55][147] = 16'b1111111111101110;
    assign weights1[55][148] = 16'b1111111111100000;
    assign weights1[55][149] = 16'b1111111111101010;
    assign weights1[55][150] = 16'b0000000000000010;
    assign weights1[55][151] = 16'b0000000000001101;
    assign weights1[55][152] = 16'b0000000000000100;
    assign weights1[55][153] = 16'b0000000000010000;
    assign weights1[55][154] = 16'b1111111111101000;
    assign weights1[55][155] = 16'b1111111111011011;
    assign weights1[55][156] = 16'b1111111111101010;
    assign weights1[55][157] = 16'b0000000000000000;
    assign weights1[55][158] = 16'b0000000000010011;
    assign weights1[55][159] = 16'b1111111111100100;
    assign weights1[55][160] = 16'b1111111111101100;
    assign weights1[55][161] = 16'b1111111111110111;
    assign weights1[55][162] = 16'b1111111111011111;
    assign weights1[55][163] = 16'b1111111111101010;
    assign weights1[55][164] = 16'b1111111111101011;
    assign weights1[55][165] = 16'b1111111111110011;
    assign weights1[55][166] = 16'b1111111111110100;
    assign weights1[55][167] = 16'b0000000000000000;
    assign weights1[55][168] = 16'b1111111111111111;
    assign weights1[55][169] = 16'b1111111111111111;
    assign weights1[55][170] = 16'b1111111111101010;
    assign weights1[55][171] = 16'b1111111111101111;
    assign weights1[55][172] = 16'b1111111111110100;
    assign weights1[55][173] = 16'b1111111111101010;
    assign weights1[55][174] = 16'b0000000000001111;
    assign weights1[55][175] = 16'b1111111111111111;
    assign weights1[55][176] = 16'b1111111111101101;
    assign weights1[55][177] = 16'b0000000000000001;
    assign weights1[55][178] = 16'b0000000000010111;
    assign weights1[55][179] = 16'b1111111111111011;
    assign weights1[55][180] = 16'b1111111111110011;
    assign weights1[55][181] = 16'b1111111111111100;
    assign weights1[55][182] = 16'b1111111111111111;
    assign weights1[55][183] = 16'b1111111111100000;
    assign weights1[55][184] = 16'b1111111111101111;
    assign weights1[55][185] = 16'b1111111111111100;
    assign weights1[55][186] = 16'b1111111111011011;
    assign weights1[55][187] = 16'b0000000000000101;
    assign weights1[55][188] = 16'b1111111111101110;
    assign weights1[55][189] = 16'b1111111111101101;
    assign weights1[55][190] = 16'b1111111111011000;
    assign weights1[55][191] = 16'b1111111111011011;
    assign weights1[55][192] = 16'b1111111111110000;
    assign weights1[55][193] = 16'b1111111111100100;
    assign weights1[55][194] = 16'b1111111111110011;
    assign weights1[55][195] = 16'b1111111111111100;
    assign weights1[55][196] = 16'b0000000000000000;
    assign weights1[55][197] = 16'b1111111111111110;
    assign weights1[55][198] = 16'b1111111111110001;
    assign weights1[55][199] = 16'b1111111111110011;
    assign weights1[55][200] = 16'b1111111111101000;
    assign weights1[55][201] = 16'b1111111111111000;
    assign weights1[55][202] = 16'b0000000000001101;
    assign weights1[55][203] = 16'b1111111111100100;
    assign weights1[55][204] = 16'b0000000000011000;
    assign weights1[55][205] = 16'b1111111111110101;
    assign weights1[55][206] = 16'b0000000000001000;
    assign weights1[55][207] = 16'b0000000000000010;
    assign weights1[55][208] = 16'b0000000000001001;
    assign weights1[55][209] = 16'b0000000000010010;
    assign weights1[55][210] = 16'b0000000000000100;
    assign weights1[55][211] = 16'b1111111111111011;
    assign weights1[55][212] = 16'b0000000000011001;
    assign weights1[55][213] = 16'b1111111111101101;
    assign weights1[55][214] = 16'b1111111111110010;
    assign weights1[55][215] = 16'b1111111111110010;
    assign weights1[55][216] = 16'b0000000000000010;
    assign weights1[55][217] = 16'b0000000000000011;
    assign weights1[55][218] = 16'b1111111111110001;
    assign weights1[55][219] = 16'b1111111111101101;
    assign weights1[55][220] = 16'b1111111111110000;
    assign weights1[55][221] = 16'b1111111111100011;
    assign weights1[55][222] = 16'b1111111111110001;
    assign weights1[55][223] = 16'b1111111111110100;
    assign weights1[55][224] = 16'b0000000000000001;
    assign weights1[55][225] = 16'b1111111111111100;
    assign weights1[55][226] = 16'b0000000000000000;
    assign weights1[55][227] = 16'b1111111111101010;
    assign weights1[55][228] = 16'b1111111111110110;
    assign weights1[55][229] = 16'b1111111111110010;
    assign weights1[55][230] = 16'b1111111111111011;
    assign weights1[55][231] = 16'b1111111111111001;
    assign weights1[55][232] = 16'b1111111111111111;
    assign weights1[55][233] = 16'b1111111111110011;
    assign weights1[55][234] = 16'b1111111111110011;
    assign weights1[55][235] = 16'b0000000000000110;
    assign weights1[55][236] = 16'b0000000000000010;
    assign weights1[55][237] = 16'b0000000000001100;
    assign weights1[55][238] = 16'b1111111111111001;
    assign weights1[55][239] = 16'b0000000000010000;
    assign weights1[55][240] = 16'b0000000000001101;
    assign weights1[55][241] = 16'b0000000000001100;
    assign weights1[55][242] = 16'b1111111111100100;
    assign weights1[55][243] = 16'b0000000000010011;
    assign weights1[55][244] = 16'b1111111111101100;
    assign weights1[55][245] = 16'b1111111111110000;
    assign weights1[55][246] = 16'b0000000000000010;
    assign weights1[55][247] = 16'b0000000000001001;
    assign weights1[55][248] = 16'b1111111111101100;
    assign weights1[55][249] = 16'b1111111111110110;
    assign weights1[55][250] = 16'b1111111111101100;
    assign weights1[55][251] = 16'b1111111111110110;
    assign weights1[55][252] = 16'b0000000000000000;
    assign weights1[55][253] = 16'b1111111111111101;
    assign weights1[55][254] = 16'b1111111111111110;
    assign weights1[55][255] = 16'b1111111111110011;
    assign weights1[55][256] = 16'b1111111111110111;
    assign weights1[55][257] = 16'b0000000000000110;
    assign weights1[55][258] = 16'b1111111111011000;
    assign weights1[55][259] = 16'b1111111111110001;
    assign weights1[55][260] = 16'b0000000000000000;
    assign weights1[55][261] = 16'b1111111111111000;
    assign weights1[55][262] = 16'b1111111111111011;
    assign weights1[55][263] = 16'b1111111111111110;
    assign weights1[55][264] = 16'b1111111111100101;
    assign weights1[55][265] = 16'b1111111111110001;
    assign weights1[55][266] = 16'b0000000000001011;
    assign weights1[55][267] = 16'b0000000000000000;
    assign weights1[55][268] = 16'b1111111111111111;
    assign weights1[55][269] = 16'b1111111111110001;
    assign weights1[55][270] = 16'b1111111111111010;
    assign weights1[55][271] = 16'b1111111111111011;
    assign weights1[55][272] = 16'b1111111111110111;
    assign weights1[55][273] = 16'b0000000000001101;
    assign weights1[55][274] = 16'b0000000000010001;
    assign weights1[55][275] = 16'b1111111111111011;
    assign weights1[55][276] = 16'b1111111111011110;
    assign weights1[55][277] = 16'b1111111111101010;
    assign weights1[55][278] = 16'b1111111111110010;
    assign weights1[55][279] = 16'b0000000000000001;
    assign weights1[55][280] = 16'b1111111111111111;
    assign weights1[55][281] = 16'b1111111111111101;
    assign weights1[55][282] = 16'b1111111111110010;
    assign weights1[55][283] = 16'b1111111111101111;
    assign weights1[55][284] = 16'b1111111111111001;
    assign weights1[55][285] = 16'b0000000000000111;
    assign weights1[55][286] = 16'b1111111111110111;
    assign weights1[55][287] = 16'b1111111111111010;
    assign weights1[55][288] = 16'b1111111111111110;
    assign weights1[55][289] = 16'b1111111111110111;
    assign weights1[55][290] = 16'b1111111111101100;
    assign weights1[55][291] = 16'b0000000000000001;
    assign weights1[55][292] = 16'b1111111111111010;
    assign weights1[55][293] = 16'b1111111111100110;
    assign weights1[55][294] = 16'b1111111111101001;
    assign weights1[55][295] = 16'b0000000000000100;
    assign weights1[55][296] = 16'b1111111111101110;
    assign weights1[55][297] = 16'b0000000000010110;
    assign weights1[55][298] = 16'b1111111111110001;
    assign weights1[55][299] = 16'b1111111111110100;
    assign weights1[55][300] = 16'b1111111111101111;
    assign weights1[55][301] = 16'b1111111111100110;
    assign weights1[55][302] = 16'b0000000000001101;
    assign weights1[55][303] = 16'b1111111111110001;
    assign weights1[55][304] = 16'b1111111111111010;
    assign weights1[55][305] = 16'b1111111111111100;
    assign weights1[55][306] = 16'b1111111111111010;
    assign weights1[55][307] = 16'b1111111111111111;
    assign weights1[55][308] = 16'b1111111111111001;
    assign weights1[55][309] = 16'b1111111111111110;
    assign weights1[55][310] = 16'b1111111111110010;
    assign weights1[55][311] = 16'b1111111111110000;
    assign weights1[55][312] = 16'b0000000000010011;
    assign weights1[55][313] = 16'b1111111111100110;
    assign weights1[55][314] = 16'b1111111111101101;
    assign weights1[55][315] = 16'b1111111111110110;
    assign weights1[55][316] = 16'b1111111111110001;
    assign weights1[55][317] = 16'b1111111111110111;
    assign weights1[55][318] = 16'b1111111111100110;
    assign weights1[55][319] = 16'b1111111111100111;
    assign weights1[55][320] = 16'b1111111111100110;
    assign weights1[55][321] = 16'b1111111111111111;
    assign weights1[55][322] = 16'b1111111111100011;
    assign weights1[55][323] = 16'b1111111111101111;
    assign weights1[55][324] = 16'b1111111111110100;
    assign weights1[55][325] = 16'b1111111111111000;
    assign weights1[55][326] = 16'b0000000000001110;
    assign weights1[55][327] = 16'b1111111111110001;
    assign weights1[55][328] = 16'b0000000000001000;
    assign weights1[55][329] = 16'b0000000000001101;
    assign weights1[55][330] = 16'b0000000000001001;
    assign weights1[55][331] = 16'b1111111111110010;
    assign weights1[55][332] = 16'b1111111111101100;
    assign weights1[55][333] = 16'b0000000000000001;
    assign weights1[55][334] = 16'b0000000000000010;
    assign weights1[55][335] = 16'b0000000000000011;
    assign weights1[55][336] = 16'b1111111111111100;
    assign weights1[55][337] = 16'b0000000000000011;
    assign weights1[55][338] = 16'b1111111111111010;
    assign weights1[55][339] = 16'b0000000000000000;
    assign weights1[55][340] = 16'b0000000000000000;
    assign weights1[55][341] = 16'b1111111111100010;
    assign weights1[55][342] = 16'b1111111111101110;
    assign weights1[55][343] = 16'b1111111111111001;
    assign weights1[55][344] = 16'b1111111111100101;
    assign weights1[55][345] = 16'b1111111111110011;
    assign weights1[55][346] = 16'b1111111111110011;
    assign weights1[55][347] = 16'b1111111111110110;
    assign weights1[55][348] = 16'b1111111111101111;
    assign weights1[55][349] = 16'b1111111111101001;
    assign weights1[55][350] = 16'b1111111111100000;
    assign weights1[55][351] = 16'b1111111111101100;
    assign weights1[55][352] = 16'b1111111111111001;
    assign weights1[55][353] = 16'b1111111111101000;
    assign weights1[55][354] = 16'b1111111111101101;
    assign weights1[55][355] = 16'b0000000000000100;
    assign weights1[55][356] = 16'b1111111111110000;
    assign weights1[55][357] = 16'b1111111111110010;
    assign weights1[55][358] = 16'b0000000000001011;
    assign weights1[55][359] = 16'b0000000000001100;
    assign weights1[55][360] = 16'b0000000000000000;
    assign weights1[55][361] = 16'b1111111111110110;
    assign weights1[55][362] = 16'b1111111111101000;
    assign weights1[55][363] = 16'b1111111111101111;
    assign weights1[55][364] = 16'b1111111111111011;
    assign weights1[55][365] = 16'b1111111111111000;
    assign weights1[55][366] = 16'b1111111111101101;
    assign weights1[55][367] = 16'b1111111111110010;
    assign weights1[55][368] = 16'b1111111111111111;
    assign weights1[55][369] = 16'b1111111111100101;
    assign weights1[55][370] = 16'b1111111111101000;
    assign weights1[55][371] = 16'b1111111111110101;
    assign weights1[55][372] = 16'b1111111111101110;
    assign weights1[55][373] = 16'b1111111111101000;
    assign weights1[55][374] = 16'b1111111111100100;
    assign weights1[55][375] = 16'b1111111111001111;
    assign weights1[55][376] = 16'b1111111111010000;
    assign weights1[55][377] = 16'b1111111111001101;
    assign weights1[55][378] = 16'b1111111111100101;
    assign weights1[55][379] = 16'b1111111111011000;
    assign weights1[55][380] = 16'b1111111111001000;
    assign weights1[55][381] = 16'b1111111111110100;
    assign weights1[55][382] = 16'b1111111111101101;
    assign weights1[55][383] = 16'b1111111111110111;
    assign weights1[55][384] = 16'b1111111111110001;
    assign weights1[55][385] = 16'b1111111111111001;
    assign weights1[55][386] = 16'b1111111111111010;
    assign weights1[55][387] = 16'b1111111111110101;
    assign weights1[55][388] = 16'b1111111111101101;
    assign weights1[55][389] = 16'b1111111111111000;
    assign weights1[55][390] = 16'b0000000000000011;
    assign weights1[55][391] = 16'b1111111111110110;
    assign weights1[55][392] = 16'b0000000000000110;
    assign weights1[55][393] = 16'b1111111111110110;
    assign weights1[55][394] = 16'b1111111111110000;
    assign weights1[55][395] = 16'b1111111111101000;
    assign weights1[55][396] = 16'b1111111111110000;
    assign weights1[55][397] = 16'b1111111111110010;
    assign weights1[55][398] = 16'b1111111111110000;
    assign weights1[55][399] = 16'b1111111111100111;
    assign weights1[55][400] = 16'b1111111111111111;
    assign weights1[55][401] = 16'b1111111111000100;
    assign weights1[55][402] = 16'b1111111111011010;
    assign weights1[55][403] = 16'b1111111111100011;
    assign weights1[55][404] = 16'b1111111111011101;
    assign weights1[55][405] = 16'b1111111111100100;
    assign weights1[55][406] = 16'b1111111111001001;
    assign weights1[55][407] = 16'b1111111111000110;
    assign weights1[55][408] = 16'b1111111111011011;
    assign weights1[55][409] = 16'b1111111111010111;
    assign weights1[55][410] = 16'b1111111111001101;
    assign weights1[55][411] = 16'b1111111110110111;
    assign weights1[55][412] = 16'b1111111111000101;
    assign weights1[55][413] = 16'b1111111111011101;
    assign weights1[55][414] = 16'b1111111111011111;
    assign weights1[55][415] = 16'b1111111111101100;
    assign weights1[55][416] = 16'b1111111111011110;
    assign weights1[55][417] = 16'b1111111111110001;
    assign weights1[55][418] = 16'b1111111111110100;
    assign weights1[55][419] = 16'b1111111111110101;
    assign weights1[55][420] = 16'b0000000000000001;
    assign weights1[55][421] = 16'b1111111111111000;
    assign weights1[55][422] = 16'b1111111111111000;
    assign weights1[55][423] = 16'b1111111111110010;
    assign weights1[55][424] = 16'b1111111111011110;
    assign weights1[55][425] = 16'b1111111111101100;
    assign weights1[55][426] = 16'b1111111111110011;
    assign weights1[55][427] = 16'b1111111111100111;
    assign weights1[55][428] = 16'b1111111111001010;
    assign weights1[55][429] = 16'b1111111110111111;
    assign weights1[55][430] = 16'b1111111110111111;
    assign weights1[55][431] = 16'b1111111111001000;
    assign weights1[55][432] = 16'b1111111110111101;
    assign weights1[55][433] = 16'b1111111111000111;
    assign weights1[55][434] = 16'b1111111111010100;
    assign weights1[55][435] = 16'b1111111110101111;
    assign weights1[55][436] = 16'b1111111111010000;
    assign weights1[55][437] = 16'b1111111110110001;
    assign weights1[55][438] = 16'b1111111110111000;
    assign weights1[55][439] = 16'b1111111110111100;
    assign weights1[55][440] = 16'b1111111111000011;
    assign weights1[55][441] = 16'b1111111111001001;
    assign weights1[55][442] = 16'b1111111111011110;
    assign weights1[55][443] = 16'b1111111111001111;
    assign weights1[55][444] = 16'b1111111111110000;
    assign weights1[55][445] = 16'b1111111111101010;
    assign weights1[55][446] = 16'b1111111111101111;
    assign weights1[55][447] = 16'b1111111111110111;
    assign weights1[55][448] = 16'b0000000000001001;
    assign weights1[55][449] = 16'b0000000000000011;
    assign weights1[55][450] = 16'b0000000000000110;
    assign weights1[55][451] = 16'b0000000000000000;
    assign weights1[55][452] = 16'b0000000000000000;
    assign weights1[55][453] = 16'b1111111111111011;
    assign weights1[55][454] = 16'b1111111111100101;
    assign weights1[55][455] = 16'b1111111110111110;
    assign weights1[55][456] = 16'b1111111111001001;
    assign weights1[55][457] = 16'b1111111110101011;
    assign weights1[55][458] = 16'b1111111110110111;
    assign weights1[55][459] = 16'b1111111110111101;
    assign weights1[55][460] = 16'b1111111111011100;
    assign weights1[55][461] = 16'b1111111111001111;
    assign weights1[55][462] = 16'b1111111111001101;
    assign weights1[55][463] = 16'b1111111110111110;
    assign weights1[55][464] = 16'b1111111111100101;
    assign weights1[55][465] = 16'b1111111110111000;
    assign weights1[55][466] = 16'b1111111111010010;
    assign weights1[55][467] = 16'b1111111111000110;
    assign weights1[55][468] = 16'b1111111111000110;
    assign weights1[55][469] = 16'b1111111111000011;
    assign weights1[55][470] = 16'b1111111111001001;
    assign weights1[55][471] = 16'b1111111111001110;
    assign weights1[55][472] = 16'b1111111111100101;
    assign weights1[55][473] = 16'b1111111111101100;
    assign weights1[55][474] = 16'b1111111111111001;
    assign weights1[55][475] = 16'b1111111111111111;
    assign weights1[55][476] = 16'b0000000000000101;
    assign weights1[55][477] = 16'b0000000000010110;
    assign weights1[55][478] = 16'b0000000000011100;
    assign weights1[55][479] = 16'b0000000000010011;
    assign weights1[55][480] = 16'b0000000000011111;
    assign weights1[55][481] = 16'b0000000000011110;
    assign weights1[55][482] = 16'b0000000000010001;
    assign weights1[55][483] = 16'b0000000000100100;
    assign weights1[55][484] = 16'b1111111111101110;
    assign weights1[55][485] = 16'b1111111111101111;
    assign weights1[55][486] = 16'b1111111111011010;
    assign weights1[55][487] = 16'b1111111111010001;
    assign weights1[55][488] = 16'b1111111111101011;
    assign weights1[55][489] = 16'b1111111111011010;
    assign weights1[55][490] = 16'b1111111110111000;
    assign weights1[55][491] = 16'b1111111111010001;
    assign weights1[55][492] = 16'b1111111110110101;
    assign weights1[55][493] = 16'b1111111111000011;
    assign weights1[55][494] = 16'b1111111111001001;
    assign weights1[55][495] = 16'b1111111111001110;
    assign weights1[55][496] = 16'b1111111110111001;
    assign weights1[55][497] = 16'b1111111110111011;
    assign weights1[55][498] = 16'b1111111111011011;
    assign weights1[55][499] = 16'b1111111111101001;
    assign weights1[55][500] = 16'b1111111111100011;
    assign weights1[55][501] = 16'b1111111111110100;
    assign weights1[55][502] = 16'b0000000000010010;
    assign weights1[55][503] = 16'b0000000000010110;
    assign weights1[55][504] = 16'b0000000000010000;
    assign weights1[55][505] = 16'b0000000000100011;
    assign weights1[55][506] = 16'b0000000000101101;
    assign weights1[55][507] = 16'b0000000000011110;
    assign weights1[55][508] = 16'b0000000000101001;
    assign weights1[55][509] = 16'b0000000000110100;
    assign weights1[55][510] = 16'b0000000000010000;
    assign weights1[55][511] = 16'b0000000000100101;
    assign weights1[55][512] = 16'b0000000000100110;
    assign weights1[55][513] = 16'b0000000000011001;
    assign weights1[55][514] = 16'b0000000000000010;
    assign weights1[55][515] = 16'b1111111111110101;
    assign weights1[55][516] = 16'b1111111111111001;
    assign weights1[55][517] = 16'b1111111111110011;
    assign weights1[55][518] = 16'b1111111110111100;
    assign weights1[55][519] = 16'b1111111111010001;
    assign weights1[55][520] = 16'b1111111111100101;
    assign weights1[55][521] = 16'b1111111111001101;
    assign weights1[55][522] = 16'b1111111111011100;
    assign weights1[55][523] = 16'b1111111111010111;
    assign weights1[55][524] = 16'b1111111111100000;
    assign weights1[55][525] = 16'b1111111111011011;
    assign weights1[55][526] = 16'b1111111111111010;
    assign weights1[55][527] = 16'b1111111111110000;
    assign weights1[55][528] = 16'b1111111111100111;
    assign weights1[55][529] = 16'b0000000000000101;
    assign weights1[55][530] = 16'b0000000000011011;
    assign weights1[55][531] = 16'b0000000000100010;
    assign weights1[55][532] = 16'b0000000000011011;
    assign weights1[55][533] = 16'b0000000000101000;
    assign weights1[55][534] = 16'b0000000000101101;
    assign weights1[55][535] = 16'b0000000000100111;
    assign weights1[55][536] = 16'b0000000000101000;
    assign weights1[55][537] = 16'b0000000000010001;
    assign weights1[55][538] = 16'b0000000000011111;
    assign weights1[55][539] = 16'b0000000000101111;
    assign weights1[55][540] = 16'b0000000000100000;
    assign weights1[55][541] = 16'b0000000000001000;
    assign weights1[55][542] = 16'b0000000000001111;
    assign weights1[55][543] = 16'b0000000000001100;
    assign weights1[55][544] = 16'b0000000000000101;
    assign weights1[55][545] = 16'b1111111111111111;
    assign weights1[55][546] = 16'b1111111111110110;
    assign weights1[55][547] = 16'b1111111111110001;
    assign weights1[55][548] = 16'b1111111111100110;
    assign weights1[55][549] = 16'b1111111111101000;
    assign weights1[55][550] = 16'b1111111111110011;
    assign weights1[55][551] = 16'b1111111111111011;
    assign weights1[55][552] = 16'b0000000000000111;
    assign weights1[55][553] = 16'b1111111111110101;
    assign weights1[55][554] = 16'b1111111111110100;
    assign weights1[55][555] = 16'b1111111111111100;
    assign weights1[55][556] = 16'b0000000000001111;
    assign weights1[55][557] = 16'b0000000000100001;
    assign weights1[55][558] = 16'b0000000000011110;
    assign weights1[55][559] = 16'b0000000000100011;
    assign weights1[55][560] = 16'b0000000000011100;
    assign weights1[55][561] = 16'b0000000000101000;
    assign weights1[55][562] = 16'b0000000000011011;
    assign weights1[55][563] = 16'b0000000000110010;
    assign weights1[55][564] = 16'b0000000000100010;
    assign weights1[55][565] = 16'b0000000000101111;
    assign weights1[55][566] = 16'b0000000000101100;
    assign weights1[55][567] = 16'b0000000000100100;
    assign weights1[55][568] = 16'b0000000000011010;
    assign weights1[55][569] = 16'b0000000000111001;
    assign weights1[55][570] = 16'b0000000001001001;
    assign weights1[55][571] = 16'b0000000000010110;
    assign weights1[55][572] = 16'b0000000000111100;
    assign weights1[55][573] = 16'b0000000000111001;
    assign weights1[55][574] = 16'b0000000000111101;
    assign weights1[55][575] = 16'b0000000000011001;
    assign weights1[55][576] = 16'b0000000000101010;
    assign weights1[55][577] = 16'b1111111111111111;
    assign weights1[55][578] = 16'b0000000000101010;
    assign weights1[55][579] = 16'b0000000000100000;
    assign weights1[55][580] = 16'b0000000000001001;
    assign weights1[55][581] = 16'b0000000000010010;
    assign weights1[55][582] = 16'b0000000000110000;
    assign weights1[55][583] = 16'b0000000000101010;
    assign weights1[55][584] = 16'b0000000000101100;
    assign weights1[55][585] = 16'b0000000000110000;
    assign weights1[55][586] = 16'b0000000000100100;
    assign weights1[55][587] = 16'b0000000000100000;
    assign weights1[55][588] = 16'b0000000000011111;
    assign weights1[55][589] = 16'b0000000000101001;
    assign weights1[55][590] = 16'b0000000000101000;
    assign weights1[55][591] = 16'b0000000000101000;
    assign weights1[55][592] = 16'b0000000000011100;
    assign weights1[55][593] = 16'b0000000000100111;
    assign weights1[55][594] = 16'b0000000001000001;
    assign weights1[55][595] = 16'b0000000000101000;
    assign weights1[55][596] = 16'b0000000000100110;
    assign weights1[55][597] = 16'b0000000000110000;
    assign weights1[55][598] = 16'b0000000000111010;
    assign weights1[55][599] = 16'b0000000001010011;
    assign weights1[55][600] = 16'b0000000000111101;
    assign weights1[55][601] = 16'b0000000000111110;
    assign weights1[55][602] = 16'b0000000001011011;
    assign weights1[55][603] = 16'b0000000001011001;
    assign weights1[55][604] = 16'b0000000001001001;
    assign weights1[55][605] = 16'b0000000001001110;
    assign weights1[55][606] = 16'b0000000001001010;
    assign weights1[55][607] = 16'b0000000001000101;
    assign weights1[55][608] = 16'b0000000000111111;
    assign weights1[55][609] = 16'b0000000000101110;
    assign weights1[55][610] = 16'b0000000000111000;
    assign weights1[55][611] = 16'b0000000000111001;
    assign weights1[55][612] = 16'b0000000000110010;
    assign weights1[55][613] = 16'b0000000000111001;
    assign weights1[55][614] = 16'b0000000000101100;
    assign weights1[55][615] = 16'b0000000000100101;
    assign weights1[55][616] = 16'b0000000000011011;
    assign weights1[55][617] = 16'b0000000000100011;
    assign weights1[55][618] = 16'b0000000000100011;
    assign weights1[55][619] = 16'b0000000000100011;
    assign weights1[55][620] = 16'b0000000000100000;
    assign weights1[55][621] = 16'b0000000000110000;
    assign weights1[55][622] = 16'b0000000000111101;
    assign weights1[55][623] = 16'b0000000000100111;
    assign weights1[55][624] = 16'b0000000000111111;
    assign weights1[55][625] = 16'b0000000001000101;
    assign weights1[55][626] = 16'b0000000000011110;
    assign weights1[55][627] = 16'b0000000001000000;
    assign weights1[55][628] = 16'b0000000000101111;
    assign weights1[55][629] = 16'b0000000000110110;
    assign weights1[55][630] = 16'b0000000000110100;
    assign weights1[55][631] = 16'b0000000001000010;
    assign weights1[55][632] = 16'b0000000000110011;
    assign weights1[55][633] = 16'b0000000001000011;
    assign weights1[55][634] = 16'b0000000000011001;
    assign weights1[55][635] = 16'b0000000000011010;
    assign weights1[55][636] = 16'b0000000001001100;
    assign weights1[55][637] = 16'b0000000000101110;
    assign weights1[55][638] = 16'b0000000000111010;
    assign weights1[55][639] = 16'b0000000000101101;
    assign weights1[55][640] = 16'b0000000000111001;
    assign weights1[55][641] = 16'b0000000000111100;
    assign weights1[55][642] = 16'b0000000000101101;
    assign weights1[55][643] = 16'b0000000000011100;
    assign weights1[55][644] = 16'b0000000000011010;
    assign weights1[55][645] = 16'b0000000000011101;
    assign weights1[55][646] = 16'b0000000000101110;
    assign weights1[55][647] = 16'b0000000000001101;
    assign weights1[55][648] = 16'b0000000000101000;
    assign weights1[55][649] = 16'b0000000000100111;
    assign weights1[55][650] = 16'b0000000000010111;
    assign weights1[55][651] = 16'b0000000000101001;
    assign weights1[55][652] = 16'b0000000000100110;
    assign weights1[55][653] = 16'b0000000000110101;
    assign weights1[55][654] = 16'b0000000000100000;
    assign weights1[55][655] = 16'b0000000000110101;
    assign weights1[55][656] = 16'b0000000000111100;
    assign weights1[55][657] = 16'b0000000000101110;
    assign weights1[55][658] = 16'b0000000000100000;
    assign weights1[55][659] = 16'b0000000001001101;
    assign weights1[55][660] = 16'b0000000001000011;
    assign weights1[55][661] = 16'b0000000000111001;
    assign weights1[55][662] = 16'b0000000000101000;
    assign weights1[55][663] = 16'b0000000001001011;
    assign weights1[55][664] = 16'b0000000000111100;
    assign weights1[55][665] = 16'b0000000000101110;
    assign weights1[55][666] = 16'b0000000000101111;
    assign weights1[55][667] = 16'b0000000000101111;
    assign weights1[55][668] = 16'b0000000000110010;
    assign weights1[55][669] = 16'b0000000000111010;
    assign weights1[55][670] = 16'b0000000000101001;
    assign weights1[55][671] = 16'b0000000000011001;
    assign weights1[55][672] = 16'b0000000000010001;
    assign weights1[55][673] = 16'b0000000000001110;
    assign weights1[55][674] = 16'b0000000000011000;
    assign weights1[55][675] = 16'b0000000000010011;
    assign weights1[55][676] = 16'b0000000000010100;
    assign weights1[55][677] = 16'b0000000000001010;
    assign weights1[55][678] = 16'b0000000000100100;
    assign weights1[55][679] = 16'b0000000000110000;
    assign weights1[55][680] = 16'b0000000000010001;
    assign weights1[55][681] = 16'b0000000000001110;
    assign weights1[55][682] = 16'b0000000000001010;
    assign weights1[55][683] = 16'b0000000000100110;
    assign weights1[55][684] = 16'b0000000000100001;
    assign weights1[55][685] = 16'b0000000000111110;
    assign weights1[55][686] = 16'b0000000001000010;
    assign weights1[55][687] = 16'b0000000000101001;
    assign weights1[55][688] = 16'b0000000000101011;
    assign weights1[55][689] = 16'b0000000001000101;
    assign weights1[55][690] = 16'b0000000001000000;
    assign weights1[55][691] = 16'b0000000000110100;
    assign weights1[55][692] = 16'b0000000000110100;
    assign weights1[55][693] = 16'b0000000001000011;
    assign weights1[55][694] = 16'b0000000000110011;
    assign weights1[55][695] = 16'b0000000000101110;
    assign weights1[55][696] = 16'b0000000000101111;
    assign weights1[55][697] = 16'b0000000000100010;
    assign weights1[55][698] = 16'b0000000000100000;
    assign weights1[55][699] = 16'b0000000000010010;
    assign weights1[55][700] = 16'b0000000000000100;
    assign weights1[55][701] = 16'b0000000000001011;
    assign weights1[55][702] = 16'b0000000000001111;
    assign weights1[55][703] = 16'b0000000000001100;
    assign weights1[55][704] = 16'b0000000000011001;
    assign weights1[55][705] = 16'b0000000000000011;
    assign weights1[55][706] = 16'b0000000000010011;
    assign weights1[55][707] = 16'b1111111111110110;
    assign weights1[55][708] = 16'b0000000000100010;
    assign weights1[55][709] = 16'b0000000000010001;
    assign weights1[55][710] = 16'b0000000000011101;
    assign weights1[55][711] = 16'b0000000000100100;
    assign weights1[55][712] = 16'b0000000000010100;
    assign weights1[55][713] = 16'b0000000000011011;
    assign weights1[55][714] = 16'b0000000000001101;
    assign weights1[55][715] = 16'b0000000000100000;
    assign weights1[55][716] = 16'b0000000000101001;
    assign weights1[55][717] = 16'b0000000000111010;
    assign weights1[55][718] = 16'b0000000000110011;
    assign weights1[55][719] = 16'b0000000001001011;
    assign weights1[55][720] = 16'b0000000000101011;
    assign weights1[55][721] = 16'b0000000000011000;
    assign weights1[55][722] = 16'b0000000000101010;
    assign weights1[55][723] = 16'b0000000000110010;
    assign weights1[55][724] = 16'b0000000000100011;
    assign weights1[55][725] = 16'b0000000000100001;
    assign weights1[55][726] = 16'b0000000000010110;
    assign weights1[55][727] = 16'b0000000000000110;
    assign weights1[55][728] = 16'b0000000000000011;
    assign weights1[55][729] = 16'b0000000000000111;
    assign weights1[55][730] = 16'b1111111111111111;
    assign weights1[55][731] = 16'b0000000000000010;
    assign weights1[55][732] = 16'b0000000000010110;
    assign weights1[55][733] = 16'b0000000000000111;
    assign weights1[55][734] = 16'b0000000000000110;
    assign weights1[55][735] = 16'b0000000000000100;
    assign weights1[55][736] = 16'b0000000000010011;
    assign weights1[55][737] = 16'b0000000000001001;
    assign weights1[55][738] = 16'b0000000000010101;
    assign weights1[55][739] = 16'b0000000000011011;
    assign weights1[55][740] = 16'b0000000000001100;
    assign weights1[55][741] = 16'b1111111111111011;
    assign weights1[55][742] = 16'b0000000000001110;
    assign weights1[55][743] = 16'b0000000000001101;
    assign weights1[55][744] = 16'b0000000000000011;
    assign weights1[55][745] = 16'b1111111111110110;
    assign weights1[55][746] = 16'b1111111111111110;
    assign weights1[55][747] = 16'b0000000000001111;
    assign weights1[55][748] = 16'b0000000000001010;
    assign weights1[55][749] = 16'b0000000000100001;
    assign weights1[55][750] = 16'b0000000000100000;
    assign weights1[55][751] = 16'b0000000000011001;
    assign weights1[55][752] = 16'b0000000000001111;
    assign weights1[55][753] = 16'b0000000000000001;
    assign weights1[55][754] = 16'b0000000000000111;
    assign weights1[55][755] = 16'b0000000000000001;
    assign weights1[55][756] = 16'b1111111111111101;
    assign weights1[55][757] = 16'b1111111111111010;
    assign weights1[55][758] = 16'b0000000000000010;
    assign weights1[55][759] = 16'b0000000000000111;
    assign weights1[55][760] = 16'b0000000000001001;
    assign weights1[55][761] = 16'b1111111111111101;
    assign weights1[55][762] = 16'b0000000000010000;
    assign weights1[55][763] = 16'b0000000000001000;
    assign weights1[55][764] = 16'b1111111111111110;
    assign weights1[55][765] = 16'b1111111111101011;
    assign weights1[55][766] = 16'b1111111111110101;
    assign weights1[55][767] = 16'b1111111111110101;
    assign weights1[55][768] = 16'b1111111111110001;
    assign weights1[55][769] = 16'b1111111111100110;
    assign weights1[55][770] = 16'b1111111111101101;
    assign weights1[55][771] = 16'b1111111111110110;
    assign weights1[55][772] = 16'b1111111111111111;
    assign weights1[55][773] = 16'b0000000000000100;
    assign weights1[55][774] = 16'b0000000000001110;
    assign weights1[55][775] = 16'b0000000000000110;
    assign weights1[55][776] = 16'b1111111111101101;
    assign weights1[55][777] = 16'b0000000000001010;
    assign weights1[55][778] = 16'b0000000000011011;
    assign weights1[55][779] = 16'b0000000000001000;
    assign weights1[55][780] = 16'b0000000000000110;
    assign weights1[55][781] = 16'b0000000000000010;
    assign weights1[55][782] = 16'b0000000000000001;
    assign weights1[55][783] = 16'b0000000000000000;
    assign weights1[56][0] = 16'b0000000000000000;
    assign weights1[56][1] = 16'b1111111111111111;
    assign weights1[56][2] = 16'b1111111111111011;
    assign weights1[56][3] = 16'b1111111111110101;
    assign weights1[56][4] = 16'b1111111111110010;
    assign weights1[56][5] = 16'b1111111111110001;
    assign weights1[56][6] = 16'b1111111111101110;
    assign weights1[56][7] = 16'b1111111111100111;
    assign weights1[56][8] = 16'b1111111111100100;
    assign weights1[56][9] = 16'b1111111111100101;
    assign weights1[56][10] = 16'b1111111111101000;
    assign weights1[56][11] = 16'b1111111111101100;
    assign weights1[56][12] = 16'b1111111111101111;
    assign weights1[56][13] = 16'b1111111111110111;
    assign weights1[56][14] = 16'b1111111111111010;
    assign weights1[56][15] = 16'b1111111111110100;
    assign weights1[56][16] = 16'b1111111111110010;
    assign weights1[56][17] = 16'b1111111111101010;
    assign weights1[56][18] = 16'b1111111111110001;
    assign weights1[56][19] = 16'b1111111111101011;
    assign weights1[56][20] = 16'b1111111111110011;
    assign weights1[56][21] = 16'b1111111111111000;
    assign weights1[56][22] = 16'b0000000000000011;
    assign weights1[56][23] = 16'b1111111111111010;
    assign weights1[56][24] = 16'b0000000000000101;
    assign weights1[56][25] = 16'b1111111111111110;
    assign weights1[56][26] = 16'b0000000000000001;
    assign weights1[56][27] = 16'b1111111111111100;
    assign weights1[56][28] = 16'b0000000000000000;
    assign weights1[56][29] = 16'b1111111111111101;
    assign weights1[56][30] = 16'b1111111111110101;
    assign weights1[56][31] = 16'b1111111111101110;
    assign weights1[56][32] = 16'b1111111111101100;
    assign weights1[56][33] = 16'b1111111111101010;
    assign weights1[56][34] = 16'b1111111111100010;
    assign weights1[56][35] = 16'b1111111111011100;
    assign weights1[56][36] = 16'b1111111111100001;
    assign weights1[56][37] = 16'b1111111111011000;
    assign weights1[56][38] = 16'b1111111111011000;
    assign weights1[56][39] = 16'b1111111111011000;
    assign weights1[56][40] = 16'b1111111111100010;
    assign weights1[56][41] = 16'b1111111111100011;
    assign weights1[56][42] = 16'b1111111111101000;
    assign weights1[56][43] = 16'b1111111111011100;
    assign weights1[56][44] = 16'b1111111111010011;
    assign weights1[56][45] = 16'b1111111111011110;
    assign weights1[56][46] = 16'b1111111111100100;
    assign weights1[56][47] = 16'b1111111111100110;
    assign weights1[56][48] = 16'b1111111111101010;
    assign weights1[56][49] = 16'b1111111111110010;
    assign weights1[56][50] = 16'b1111111111101011;
    assign weights1[56][51] = 16'b1111111111110010;
    assign weights1[56][52] = 16'b1111111111111101;
    assign weights1[56][53] = 16'b0000000000000011;
    assign weights1[56][54] = 16'b1111111111111001;
    assign weights1[56][55] = 16'b1111111111110110;
    assign weights1[56][56] = 16'b1111111111111101;
    assign weights1[56][57] = 16'b1111111111111001;
    assign weights1[56][58] = 16'b1111111111110010;
    assign weights1[56][59] = 16'b1111111111101001;
    assign weights1[56][60] = 16'b1111111111100100;
    assign weights1[56][61] = 16'b1111111111011111;
    assign weights1[56][62] = 16'b1111111111011001;
    assign weights1[56][63] = 16'b1111111111010000;
    assign weights1[56][64] = 16'b1111111111001100;
    assign weights1[56][65] = 16'b1111111111000100;
    assign weights1[56][66] = 16'b1111111111001000;
    assign weights1[56][67] = 16'b1111111111001000;
    assign weights1[56][68] = 16'b1111111111001011;
    assign weights1[56][69] = 16'b1111111111000010;
    assign weights1[56][70] = 16'b1111111110110110;
    assign weights1[56][71] = 16'b1111111110111110;
    assign weights1[56][72] = 16'b1111111111000100;
    assign weights1[56][73] = 16'b1111111111001111;
    assign weights1[56][74] = 16'b1111111111001011;
    assign weights1[56][75] = 16'b1111111111001001;
    assign weights1[56][76] = 16'b1111111111011001;
    assign weights1[56][77] = 16'b1111111111011100;
    assign weights1[56][78] = 16'b1111111111100000;
    assign weights1[56][79] = 16'b1111111111110011;
    assign weights1[56][80] = 16'b1111111111101001;
    assign weights1[56][81] = 16'b1111111111101001;
    assign weights1[56][82] = 16'b1111111111110010;
    assign weights1[56][83] = 16'b1111111111110000;
    assign weights1[56][84] = 16'b1111111111111101;
    assign weights1[56][85] = 16'b1111111111110010;
    assign weights1[56][86] = 16'b1111111111101100;
    assign weights1[56][87] = 16'b1111111111100010;
    assign weights1[56][88] = 16'b1111111111011110;
    assign weights1[56][89] = 16'b1111111111010111;
    assign weights1[56][90] = 16'b1111111111001100;
    assign weights1[56][91] = 16'b1111111111000011;
    assign weights1[56][92] = 16'b1111111111000010;
    assign weights1[56][93] = 16'b1111111110111100;
    assign weights1[56][94] = 16'b1111111110110001;
    assign weights1[56][95] = 16'b1111111110101101;
    assign weights1[56][96] = 16'b1111111110101100;
    assign weights1[56][97] = 16'b1111111110111001;
    assign weights1[56][98] = 16'b1111111111001110;
    assign weights1[56][99] = 16'b1111111110111010;
    assign weights1[56][100] = 16'b1111111111001110;
    assign weights1[56][101] = 16'b1111111111010100;
    assign weights1[56][102] = 16'b1111111111100000;
    assign weights1[56][103] = 16'b1111111111001101;
    assign weights1[56][104] = 16'b1111111111001110;
    assign weights1[56][105] = 16'b1111111111010101;
    assign weights1[56][106] = 16'b1111111111010000;
    assign weights1[56][107] = 16'b1111111111100011;
    assign weights1[56][108] = 16'b1111111111101110;
    assign weights1[56][109] = 16'b1111111111101110;
    assign weights1[56][110] = 16'b1111111111111010;
    assign weights1[56][111] = 16'b0000000000000011;
    assign weights1[56][112] = 16'b1111111111111001;
    assign weights1[56][113] = 16'b1111111111110000;
    assign weights1[56][114] = 16'b1111111111101010;
    assign weights1[56][115] = 16'b1111111111100110;
    assign weights1[56][116] = 16'b1111111111100011;
    assign weights1[56][117] = 16'b1111111111010000;
    assign weights1[56][118] = 16'b1111111111000010;
    assign weights1[56][119] = 16'b1111111110110010;
    assign weights1[56][120] = 16'b1111111111000000;
    assign weights1[56][121] = 16'b1111111111000010;
    assign weights1[56][122] = 16'b1111111111000110;
    assign weights1[56][123] = 16'b1111111111001010;
    assign weights1[56][124] = 16'b1111111111011000;
    assign weights1[56][125] = 16'b1111111111001010;
    assign weights1[56][126] = 16'b1111111111110101;
    assign weights1[56][127] = 16'b1111111111101011;
    assign weights1[56][128] = 16'b1111111111111001;
    assign weights1[56][129] = 16'b1111111111011000;
    assign weights1[56][130] = 16'b1111111111100100;
    assign weights1[56][131] = 16'b1111111111101001;
    assign weights1[56][132] = 16'b1111111111001110;
    assign weights1[56][133] = 16'b1111111111010111;
    assign weights1[56][134] = 16'b1111111111010001;
    assign weights1[56][135] = 16'b0000000000001010;
    assign weights1[56][136] = 16'b1111111111111000;
    assign weights1[56][137] = 16'b1111111111110101;
    assign weights1[56][138] = 16'b0000000000000110;
    assign weights1[56][139] = 16'b0000000000001001;
    assign weights1[56][140] = 16'b1111111111111100;
    assign weights1[56][141] = 16'b1111111111110010;
    assign weights1[56][142] = 16'b1111111111100110;
    assign weights1[56][143] = 16'b1111111111101001;
    assign weights1[56][144] = 16'b1111111111100111;
    assign weights1[56][145] = 16'b1111111111110010;
    assign weights1[56][146] = 16'b1111111111011011;
    assign weights1[56][147] = 16'b1111111111110110;
    assign weights1[56][148] = 16'b1111111111111001;
    assign weights1[56][149] = 16'b0000000000000001;
    assign weights1[56][150] = 16'b0000000000001100;
    assign weights1[56][151] = 16'b0000000000010101;
    assign weights1[56][152] = 16'b1111111111111110;
    assign weights1[56][153] = 16'b1111111111110011;
    assign weights1[56][154] = 16'b1111111111110000;
    assign weights1[56][155] = 16'b1111111111111101;
    assign weights1[56][156] = 16'b1111111111110100;
    assign weights1[56][157] = 16'b0000000000000111;
    assign weights1[56][158] = 16'b1111111111111000;
    assign weights1[56][159] = 16'b1111111111111101;
    assign weights1[56][160] = 16'b1111111111111111;
    assign weights1[56][161] = 16'b1111111111100110;
    assign weights1[56][162] = 16'b1111111111110011;
    assign weights1[56][163] = 16'b1111111111110001;
    assign weights1[56][164] = 16'b1111111111100000;
    assign weights1[56][165] = 16'b1111111111110011;
    assign weights1[56][166] = 16'b0000000000001101;
    assign weights1[56][167] = 16'b0000000000010101;
    assign weights1[56][168] = 16'b1111111111111100;
    assign weights1[56][169] = 16'b1111111111111000;
    assign weights1[56][170] = 16'b1111111111111001;
    assign weights1[56][171] = 16'b1111111111111000;
    assign weights1[56][172] = 16'b0000000000000100;
    assign weights1[56][173] = 16'b1111111111100100;
    assign weights1[56][174] = 16'b1111111111111110;
    assign weights1[56][175] = 16'b0000000000001111;
    assign weights1[56][176] = 16'b0000000000011110;
    assign weights1[56][177] = 16'b0000000000000100;
    assign weights1[56][178] = 16'b1111111111110011;
    assign weights1[56][179] = 16'b1111111111110111;
    assign weights1[56][180] = 16'b0000000000001111;
    assign weights1[56][181] = 16'b0000000000001001;
    assign weights1[56][182] = 16'b0000000000010000;
    assign weights1[56][183] = 16'b1111111111111111;
    assign weights1[56][184] = 16'b1111111111110001;
    assign weights1[56][185] = 16'b0000000000000001;
    assign weights1[56][186] = 16'b1111111111111011;
    assign weights1[56][187] = 16'b1111111111110110;
    assign weights1[56][188] = 16'b0000000000000110;
    assign weights1[56][189] = 16'b0000000000011001;
    assign weights1[56][190] = 16'b1111111111111101;
    assign weights1[56][191] = 16'b1111111111111001;
    assign weights1[56][192] = 16'b1111111111101101;
    assign weights1[56][193] = 16'b0000000000000111;
    assign weights1[56][194] = 16'b0000000000000011;
    assign weights1[56][195] = 16'b0000000000001000;
    assign weights1[56][196] = 16'b1111111111111110;
    assign weights1[56][197] = 16'b0000000000000000;
    assign weights1[56][198] = 16'b1111111111111101;
    assign weights1[56][199] = 16'b0000000000000100;
    assign weights1[56][200] = 16'b0000000000000100;
    assign weights1[56][201] = 16'b0000000000000101;
    assign weights1[56][202] = 16'b0000000000000010;
    assign weights1[56][203] = 16'b1111111111110001;
    assign weights1[56][204] = 16'b1111111111111101;
    assign weights1[56][205] = 16'b1111111111101011;
    assign weights1[56][206] = 16'b0000000000010001;
    assign weights1[56][207] = 16'b1111111111110111;
    assign weights1[56][208] = 16'b0000000000001011;
    assign weights1[56][209] = 16'b0000000000001110;
    assign weights1[56][210] = 16'b0000000000000101;
    assign weights1[56][211] = 16'b0000000000001100;
    assign weights1[56][212] = 16'b0000000000000111;
    assign weights1[56][213] = 16'b0000000000001001;
    assign weights1[56][214] = 16'b0000000000001101;
    assign weights1[56][215] = 16'b0000000000000001;
    assign weights1[56][216] = 16'b1111111111111110;
    assign weights1[56][217] = 16'b1111111111101110;
    assign weights1[56][218] = 16'b1111111111111010;
    assign weights1[56][219] = 16'b1111111111111011;
    assign weights1[56][220] = 16'b0000000000000001;
    assign weights1[56][221] = 16'b1111111111110101;
    assign weights1[56][222] = 16'b0000000000000011;
    assign weights1[56][223] = 16'b0000000000000101;
    assign weights1[56][224] = 16'b1111111111111100;
    assign weights1[56][225] = 16'b0000000000000110;
    assign weights1[56][226] = 16'b0000000000000000;
    assign weights1[56][227] = 16'b0000000000001000;
    assign weights1[56][228] = 16'b0000000000000010;
    assign weights1[56][229] = 16'b0000000000001110;
    assign weights1[56][230] = 16'b0000000000010101;
    assign weights1[56][231] = 16'b0000000000000010;
    assign weights1[56][232] = 16'b1111111111110011;
    assign weights1[56][233] = 16'b0000000000001111;
    assign weights1[56][234] = 16'b1111111111110010;
    assign weights1[56][235] = 16'b0000000000000001;
    assign weights1[56][236] = 16'b1111111111101110;
    assign weights1[56][237] = 16'b0000000000000001;
    assign weights1[56][238] = 16'b1111111111111110;
    assign weights1[56][239] = 16'b1111111111110100;
    assign weights1[56][240] = 16'b1111111111111111;
    assign weights1[56][241] = 16'b1111111111110111;
    assign weights1[56][242] = 16'b0000000000000011;
    assign weights1[56][243] = 16'b1111111111111110;
    assign weights1[56][244] = 16'b1111111111111000;
    assign weights1[56][245] = 16'b1111111111110010;
    assign weights1[56][246] = 16'b1111111111111100;
    assign weights1[56][247] = 16'b0000000000001000;
    assign weights1[56][248] = 16'b1111111111110100;
    assign weights1[56][249] = 16'b0000000000001010;
    assign weights1[56][250] = 16'b1111111111111110;
    assign weights1[56][251] = 16'b0000000000001010;
    assign weights1[56][252] = 16'b0000000000000111;
    assign weights1[56][253] = 16'b0000000000001110;
    assign weights1[56][254] = 16'b0000000000000101;
    assign weights1[56][255] = 16'b1111111111111111;
    assign weights1[56][256] = 16'b0000000000000111;
    assign weights1[56][257] = 16'b1111111111110010;
    assign weights1[56][258] = 16'b0000000000010010;
    assign weights1[56][259] = 16'b0000000000000001;
    assign weights1[56][260] = 16'b1111111111110101;
    assign weights1[56][261] = 16'b0000000000000101;
    assign weights1[56][262] = 16'b0000000000000010;
    assign weights1[56][263] = 16'b0000000000001011;
    assign weights1[56][264] = 16'b0000000000010001;
    assign weights1[56][265] = 16'b1111111111111011;
    assign weights1[56][266] = 16'b0000000000000010;
    assign weights1[56][267] = 16'b0000000000000101;
    assign weights1[56][268] = 16'b0000000000000000;
    assign weights1[56][269] = 16'b0000000000001011;
    assign weights1[56][270] = 16'b1111111111111001;
    assign weights1[56][271] = 16'b1111111111111100;
    assign weights1[56][272] = 16'b0000000000010010;
    assign weights1[56][273] = 16'b1111111111111110;
    assign weights1[56][274] = 16'b1111111111111110;
    assign weights1[56][275] = 16'b1111111111101101;
    assign weights1[56][276] = 16'b0000000000000011;
    assign weights1[56][277] = 16'b0000000000000101;
    assign weights1[56][278] = 16'b1111111111111010;
    assign weights1[56][279] = 16'b0000000000001001;
    assign weights1[56][280] = 16'b0000000000010110;
    assign weights1[56][281] = 16'b0000000000010011;
    assign weights1[56][282] = 16'b1111111111111110;
    assign weights1[56][283] = 16'b0000000000010100;
    assign weights1[56][284] = 16'b0000000000000110;
    assign weights1[56][285] = 16'b1111111111110001;
    assign weights1[56][286] = 16'b0000000000001001;
    assign weights1[56][287] = 16'b1111111111111001;
    assign weights1[56][288] = 16'b1111111111111001;
    assign weights1[56][289] = 16'b0000000000001111;
    assign weights1[56][290] = 16'b0000000000001000;
    assign weights1[56][291] = 16'b0000000000010001;
    assign weights1[56][292] = 16'b1111111111111011;
    assign weights1[56][293] = 16'b0000000000000011;
    assign weights1[56][294] = 16'b1111111111110111;
    assign weights1[56][295] = 16'b1111111111110111;
    assign weights1[56][296] = 16'b1111111111110101;
    assign weights1[56][297] = 16'b1111111111111111;
    assign weights1[56][298] = 16'b0000000000000010;
    assign weights1[56][299] = 16'b1111111111111011;
    assign weights1[56][300] = 16'b1111111111110011;
    assign weights1[56][301] = 16'b0000000000000001;
    assign weights1[56][302] = 16'b1111111111111100;
    assign weights1[56][303] = 16'b1111111111111111;
    assign weights1[56][304] = 16'b1111111111101000;
    assign weights1[56][305] = 16'b1111111111111101;
    assign weights1[56][306] = 16'b1111111111111001;
    assign weights1[56][307] = 16'b0000000000000000;
    assign weights1[56][308] = 16'b0000000000001000;
    assign weights1[56][309] = 16'b0000000000010010;
    assign weights1[56][310] = 16'b0000000000000001;
    assign weights1[56][311] = 16'b1111111111111101;
    assign weights1[56][312] = 16'b1111111111101100;
    assign weights1[56][313] = 16'b1111111111111110;
    assign weights1[56][314] = 16'b1111111111111000;
    assign weights1[56][315] = 16'b1111111111111011;
    assign weights1[56][316] = 16'b0000000000010001;
    assign weights1[56][317] = 16'b0000000000010010;
    assign weights1[56][318] = 16'b0000000000001000;
    assign weights1[56][319] = 16'b0000000000001110;
    assign weights1[56][320] = 16'b0000000000000000;
    assign weights1[56][321] = 16'b1111111111111010;
    assign weights1[56][322] = 16'b0000000000000111;
    assign weights1[56][323] = 16'b1111111111110000;
    assign weights1[56][324] = 16'b0000000000000110;
    assign weights1[56][325] = 16'b1111111111111101;
    assign weights1[56][326] = 16'b0000000000010010;
    assign weights1[56][327] = 16'b0000000000000101;
    assign weights1[56][328] = 16'b0000000000000100;
    assign weights1[56][329] = 16'b1111111111111011;
    assign weights1[56][330] = 16'b1111111111110101;
    assign weights1[56][331] = 16'b1111111111111111;
    assign weights1[56][332] = 16'b0000000000000010;
    assign weights1[56][333] = 16'b1111111111111001;
    assign weights1[56][334] = 16'b1111111111111001;
    assign weights1[56][335] = 16'b0000000000001110;
    assign weights1[56][336] = 16'b0000000000000000;
    assign weights1[56][337] = 16'b0000000000000100;
    assign weights1[56][338] = 16'b0000000000000100;
    assign weights1[56][339] = 16'b1111111111110010;
    assign weights1[56][340] = 16'b1111111111111110;
    assign weights1[56][341] = 16'b1111111111111100;
    assign weights1[56][342] = 16'b1111111111111011;
    assign weights1[56][343] = 16'b0000000000000001;
    assign weights1[56][344] = 16'b1111111111110000;
    assign weights1[56][345] = 16'b1111111111100001;
    assign weights1[56][346] = 16'b1111111111101100;
    assign weights1[56][347] = 16'b1111111111101101;
    assign weights1[56][348] = 16'b0000000000000101;
    assign weights1[56][349] = 16'b1111111111110101;
    assign weights1[56][350] = 16'b1111111111111000;
    assign weights1[56][351] = 16'b1111111111110111;
    assign weights1[56][352] = 16'b0000000000000000;
    assign weights1[56][353] = 16'b1111111111110010;
    assign weights1[56][354] = 16'b1111111111110011;
    assign weights1[56][355] = 16'b0000000000000001;
    assign weights1[56][356] = 16'b1111111111111110;
    assign weights1[56][357] = 16'b1111111111111011;
    assign weights1[56][358] = 16'b1111111111111010;
    assign weights1[56][359] = 16'b0000000000011000;
    assign weights1[56][360] = 16'b0000000000001100;
    assign weights1[56][361] = 16'b1111111111111111;
    assign weights1[56][362] = 16'b0000000000001110;
    assign weights1[56][363] = 16'b0000000000000011;
    assign weights1[56][364] = 16'b0000000000000011;
    assign weights1[56][365] = 16'b0000000000001000;
    assign weights1[56][366] = 16'b1111111111100100;
    assign weights1[56][367] = 16'b1111111111101111;
    assign weights1[56][368] = 16'b0000000000000100;
    assign weights1[56][369] = 16'b1111111111110111;
    assign weights1[56][370] = 16'b0000000000000100;
    assign weights1[56][371] = 16'b0000000000001110;
    assign weights1[56][372] = 16'b1111111111111100;
    assign weights1[56][373] = 16'b1111111111111111;
    assign weights1[56][374] = 16'b0000000000001110;
    assign weights1[56][375] = 16'b1111111111111001;
    assign weights1[56][376] = 16'b1111111111110010;
    assign weights1[56][377] = 16'b0000000000001001;
    assign weights1[56][378] = 16'b0000000000000100;
    assign weights1[56][379] = 16'b0000000000000000;
    assign weights1[56][380] = 16'b1111111111111000;
    assign weights1[56][381] = 16'b0000000000000101;
    assign weights1[56][382] = 16'b0000000000000110;
    assign weights1[56][383] = 16'b0000000000000000;
    assign weights1[56][384] = 16'b0000000000000001;
    assign weights1[56][385] = 16'b0000000000000011;
    assign weights1[56][386] = 16'b1111111111111111;
    assign weights1[56][387] = 16'b1111111111111100;
    assign weights1[56][388] = 16'b1111111111111110;
    assign weights1[56][389] = 16'b0000000000000001;
    assign weights1[56][390] = 16'b0000000000001011;
    assign weights1[56][391] = 16'b0000000000001011;
    assign weights1[56][392] = 16'b1111111111111110;
    assign weights1[56][393] = 16'b1111111111111011;
    assign weights1[56][394] = 16'b1111111111110010;
    assign weights1[56][395] = 16'b1111111111111011;
    assign weights1[56][396] = 16'b0000000000010101;
    assign weights1[56][397] = 16'b1111111111110001;
    assign weights1[56][398] = 16'b1111111111101111;
    assign weights1[56][399] = 16'b0000000000000000;
    assign weights1[56][400] = 16'b0000000000000001;
    assign weights1[56][401] = 16'b0000000000001101;
    assign weights1[56][402] = 16'b0000000000001100;
    assign weights1[56][403] = 16'b1111111111111001;
    assign weights1[56][404] = 16'b1111111111110111;
    assign weights1[56][405] = 16'b0000000000001101;
    assign weights1[56][406] = 16'b0000000000010100;
    assign weights1[56][407] = 16'b0000000000001111;
    assign weights1[56][408] = 16'b0000000000000111;
    assign weights1[56][409] = 16'b0000000000001011;
    assign weights1[56][410] = 16'b1111111111101110;
    assign weights1[56][411] = 16'b0000000000000101;
    assign weights1[56][412] = 16'b0000000000000001;
    assign weights1[56][413] = 16'b0000000000000010;
    assign weights1[56][414] = 16'b0000000000000100;
    assign weights1[56][415] = 16'b1111111111110100;
    assign weights1[56][416] = 16'b0000000000000111;
    assign weights1[56][417] = 16'b0000000000000100;
    assign weights1[56][418] = 16'b1111111111111101;
    assign weights1[56][419] = 16'b0000000000001111;
    assign weights1[56][420] = 16'b1111111111110001;
    assign weights1[56][421] = 16'b1111111111101111;
    assign weights1[56][422] = 16'b1111111111101010;
    assign weights1[56][423] = 16'b1111111111111101;
    assign weights1[56][424] = 16'b0000000000000010;
    assign weights1[56][425] = 16'b0000000000011011;
    assign weights1[56][426] = 16'b0000000000010101;
    assign weights1[56][427] = 16'b0000000000000010;
    assign weights1[56][428] = 16'b0000000000001111;
    assign weights1[56][429] = 16'b0000000000001100;
    assign weights1[56][430] = 16'b0000000000010011;
    assign weights1[56][431] = 16'b0000000000010010;
    assign weights1[56][432] = 16'b0000000000011101;
    assign weights1[56][433] = 16'b0000000000001100;
    assign weights1[56][434] = 16'b0000000000000111;
    assign weights1[56][435] = 16'b1111111111111001;
    assign weights1[56][436] = 16'b0000000000010001;
    assign weights1[56][437] = 16'b0000000000000010;
    assign weights1[56][438] = 16'b1111111111110110;
    assign weights1[56][439] = 16'b1111111111111110;
    assign weights1[56][440] = 16'b1111111111111010;
    assign weights1[56][441] = 16'b1111111111111110;
    assign weights1[56][442] = 16'b1111111111101010;
    assign weights1[56][443] = 16'b1111111111111011;
    assign weights1[56][444] = 16'b1111111111110100;
    assign weights1[56][445] = 16'b0000000000000000;
    assign weights1[56][446] = 16'b1111111111111100;
    assign weights1[56][447] = 16'b1111111111111100;
    assign weights1[56][448] = 16'b1111111111101000;
    assign weights1[56][449] = 16'b1111111111100001;
    assign weights1[56][450] = 16'b1111111111100001;
    assign weights1[56][451] = 16'b1111111111010101;
    assign weights1[56][452] = 16'b0000000000000100;
    assign weights1[56][453] = 16'b0000000000100101;
    assign weights1[56][454] = 16'b0000000000100000;
    assign weights1[56][455] = 16'b0000000000100110;
    assign weights1[56][456] = 16'b0000000000101011;
    assign weights1[56][457] = 16'b0000000000011011;
    assign weights1[56][458] = 16'b0000000000100101;
    assign weights1[56][459] = 16'b0000000000010101;
    assign weights1[56][460] = 16'b0000000000010011;
    assign weights1[56][461] = 16'b0000000000001101;
    assign weights1[56][462] = 16'b0000000000000011;
    assign weights1[56][463] = 16'b0000000000001111;
    assign weights1[56][464] = 16'b0000000000000100;
    assign weights1[56][465] = 16'b0000000000001010;
    assign weights1[56][466] = 16'b0000000000001001;
    assign weights1[56][467] = 16'b0000000000000110;
    assign weights1[56][468] = 16'b1111111111110100;
    assign weights1[56][469] = 16'b0000000000000001;
    assign weights1[56][470] = 16'b0000000000000100;
    assign weights1[56][471] = 16'b0000000000000111;
    assign weights1[56][472] = 16'b1111111111111001;
    assign weights1[56][473] = 16'b1111111111111101;
    assign weights1[56][474] = 16'b1111111111111011;
    assign weights1[56][475] = 16'b0000000000000010;
    assign weights1[56][476] = 16'b1111111111100000;
    assign weights1[56][477] = 16'b1111111111010010;
    assign weights1[56][478] = 16'b1111111111000001;
    assign weights1[56][479] = 16'b1111111111000000;
    assign weights1[56][480] = 16'b1111111111000101;
    assign weights1[56][481] = 16'b1111111111111111;
    assign weights1[56][482] = 16'b0000000000010011;
    assign weights1[56][483] = 16'b0000000000010110;
    assign weights1[56][484] = 16'b0000000000010101;
    assign weights1[56][485] = 16'b0000000000011101;
    assign weights1[56][486] = 16'b0000000000101001;
    assign weights1[56][487] = 16'b0000000000010110;
    assign weights1[56][488] = 16'b0000000000001100;
    assign weights1[56][489] = 16'b0000000000001001;
    assign weights1[56][490] = 16'b1111111111111101;
    assign weights1[56][491] = 16'b0000000000011010;
    assign weights1[56][492] = 16'b0000000000001111;
    assign weights1[56][493] = 16'b0000000000000100;
    assign weights1[56][494] = 16'b0000000000001000;
    assign weights1[56][495] = 16'b0000000000010001;
    assign weights1[56][496] = 16'b0000000000001001;
    assign weights1[56][497] = 16'b0000000000001100;
    assign weights1[56][498] = 16'b0000000000001011;
    assign weights1[56][499] = 16'b0000000000010100;
    assign weights1[56][500] = 16'b0000000000000111;
    assign weights1[56][501] = 16'b1111111111111001;
    assign weights1[56][502] = 16'b1111111111111100;
    assign weights1[56][503] = 16'b1111111111111001;
    assign weights1[56][504] = 16'b1111111111011011;
    assign weights1[56][505] = 16'b1111111111000000;
    assign weights1[56][506] = 16'b1111111110110101;
    assign weights1[56][507] = 16'b1111111110010101;
    assign weights1[56][508] = 16'b1111111101110110;
    assign weights1[56][509] = 16'b1111111111001011;
    assign weights1[56][510] = 16'b1111111111011011;
    assign weights1[56][511] = 16'b1111111111100111;
    assign weights1[56][512] = 16'b0000000000010011;
    assign weights1[56][513] = 16'b0000000000011000;
    assign weights1[56][514] = 16'b0000000000011100;
    assign weights1[56][515] = 16'b0000000000100111;
    assign weights1[56][516] = 16'b0000000000010011;
    assign weights1[56][517] = 16'b0000000000011000;
    assign weights1[56][518] = 16'b0000000000000111;
    assign weights1[56][519] = 16'b1111111111111110;
    assign weights1[56][520] = 16'b0000000000001101;
    assign weights1[56][521] = 16'b0000000000000110;
    assign weights1[56][522] = 16'b1111111111111110;
    assign weights1[56][523] = 16'b0000000000000100;
    assign weights1[56][524] = 16'b0000000000011000;
    assign weights1[56][525] = 16'b0000000000001000;
    assign weights1[56][526] = 16'b1111111111111001;
    assign weights1[56][527] = 16'b0000000000000010;
    assign weights1[56][528] = 16'b1111111111110010;
    assign weights1[56][529] = 16'b0000000000011000;
    assign weights1[56][530] = 16'b0000000000000010;
    assign weights1[56][531] = 16'b1111111111111111;
    assign weights1[56][532] = 16'b1111111111011110;
    assign weights1[56][533] = 16'b1111111111001001;
    assign weights1[56][534] = 16'b1111111110101101;
    assign weights1[56][535] = 16'b1111111110000000;
    assign weights1[56][536] = 16'b1111111101100011;
    assign weights1[56][537] = 16'b1111111101101010;
    assign weights1[56][538] = 16'b1111111110000011;
    assign weights1[56][539] = 16'b1111111110100000;
    assign weights1[56][540] = 16'b1111111110100010;
    assign weights1[56][541] = 16'b1111111110111110;
    assign weights1[56][542] = 16'b1111111111011110;
    assign weights1[56][543] = 16'b1111111111100111;
    assign weights1[56][544] = 16'b1111111111101101;
    assign weights1[56][545] = 16'b1111111111101010;
    assign weights1[56][546] = 16'b1111111111110001;
    assign weights1[56][547] = 16'b1111111111110101;
    assign weights1[56][548] = 16'b1111111111110010;
    assign weights1[56][549] = 16'b1111111111110000;
    assign weights1[56][550] = 16'b0000000000000001;
    assign weights1[56][551] = 16'b1111111111111100;
    assign weights1[56][552] = 16'b1111111111110100;
    assign weights1[56][553] = 16'b0000000000000100;
    assign weights1[56][554] = 16'b1111111111111000;
    assign weights1[56][555] = 16'b1111111111111011;
    assign weights1[56][556] = 16'b1111111111110000;
    assign weights1[56][557] = 16'b0000000000000101;
    assign weights1[56][558] = 16'b0000000000000001;
    assign weights1[56][559] = 16'b0000000000000011;
    assign weights1[56][560] = 16'b1111111111011111;
    assign weights1[56][561] = 16'b1111111111011010;
    assign weights1[56][562] = 16'b1111111111010001;
    assign weights1[56][563] = 16'b1111111110011111;
    assign weights1[56][564] = 16'b1111111101111101;
    assign weights1[56][565] = 16'b1111111101000000;
    assign weights1[56][566] = 16'b1111111100100000;
    assign weights1[56][567] = 16'b1111111100001100;
    assign weights1[56][568] = 16'b1111111011101101;
    assign weights1[56][569] = 16'b1111111011111111;
    assign weights1[56][570] = 16'b1111111100010000;
    assign weights1[56][571] = 16'b1111111101101000;
    assign weights1[56][572] = 16'b1111111110010011;
    assign weights1[56][573] = 16'b1111111110110110;
    assign weights1[56][574] = 16'b1111111111010101;
    assign weights1[56][575] = 16'b1111111111010000;
    assign weights1[56][576] = 16'b1111111111101111;
    assign weights1[56][577] = 16'b1111111111111100;
    assign weights1[56][578] = 16'b1111111111111101;
    assign weights1[56][579] = 16'b0000000000000011;
    assign weights1[56][580] = 16'b0000000000000000;
    assign weights1[56][581] = 16'b0000000000010000;
    assign weights1[56][582] = 16'b0000000000000110;
    assign weights1[56][583] = 16'b0000000000000000;
    assign weights1[56][584] = 16'b1111111111111011;
    assign weights1[56][585] = 16'b0000000000010010;
    assign weights1[56][586] = 16'b1111111111110101;
    assign weights1[56][587] = 16'b1111111111101001;
    assign weights1[56][588] = 16'b1111111111110000;
    assign weights1[56][589] = 16'b1111111111110101;
    assign weights1[56][590] = 16'b1111111111101101;
    assign weights1[56][591] = 16'b1111111111011101;
    assign weights1[56][592] = 16'b1111111111000110;
    assign weights1[56][593] = 16'b1111111110101001;
    assign weights1[56][594] = 16'b1111111110101100;
    assign weights1[56][595] = 16'b1111111110000111;
    assign weights1[56][596] = 16'b1111111101110111;
    assign weights1[56][597] = 16'b1111111110000010;
    assign weights1[56][598] = 16'b1111111110011110;
    assign weights1[56][599] = 16'b1111111110101010;
    assign weights1[56][600] = 16'b1111111111000000;
    assign weights1[56][601] = 16'b1111111111011001;
    assign weights1[56][602] = 16'b1111111111110001;
    assign weights1[56][603] = 16'b1111111111111001;
    assign weights1[56][604] = 16'b1111111111110010;
    assign weights1[56][605] = 16'b1111111111110111;
    assign weights1[56][606] = 16'b0000000000001111;
    assign weights1[56][607] = 16'b1111111111111110;
    assign weights1[56][608] = 16'b0000000000010001;
    assign weights1[56][609] = 16'b0000000000000010;
    assign weights1[56][610] = 16'b0000000000001000;
    assign weights1[56][611] = 16'b0000000000001101;
    assign weights1[56][612] = 16'b1111111111111111;
    assign weights1[56][613] = 16'b0000000000000110;
    assign weights1[56][614] = 16'b1111111111111100;
    assign weights1[56][615] = 16'b1111111111100111;
    assign weights1[56][616] = 16'b1111111111101011;
    assign weights1[56][617] = 16'b1111111111110101;
    assign weights1[56][618] = 16'b0000000000001100;
    assign weights1[56][619] = 16'b0000000000010011;
    assign weights1[56][620] = 16'b0000000000001000;
    assign weights1[56][621] = 16'b0000000000000000;
    assign weights1[56][622] = 16'b0000000000001101;
    assign weights1[56][623] = 16'b0000000000001011;
    assign weights1[56][624] = 16'b0000000001000000;
    assign weights1[56][625] = 16'b0000000000100010;
    assign weights1[56][626] = 16'b0000000000111000;
    assign weights1[56][627] = 16'b0000000000101101;
    assign weights1[56][628] = 16'b0000000000011101;
    assign weights1[56][629] = 16'b0000000000010001;
    assign weights1[56][630] = 16'b0000000000000110;
    assign weights1[56][631] = 16'b0000000000000100;
    assign weights1[56][632] = 16'b0000000000000010;
    assign weights1[56][633] = 16'b0000000000000000;
    assign weights1[56][634] = 16'b1111111111101110;
    assign weights1[56][635] = 16'b1111111111101111;
    assign weights1[56][636] = 16'b0000000000001111;
    assign weights1[56][637] = 16'b1111111111111101;
    assign weights1[56][638] = 16'b0000000000000110;
    assign weights1[56][639] = 16'b0000000000000101;
    assign weights1[56][640] = 16'b0000000000000010;
    assign weights1[56][641] = 16'b0000000000000011;
    assign weights1[56][642] = 16'b1111111111110011;
    assign weights1[56][643] = 16'b1111111111101101;
    assign weights1[56][644] = 16'b1111111111110110;
    assign weights1[56][645] = 16'b1111111111110110;
    assign weights1[56][646] = 16'b0000000000001100;
    assign weights1[56][647] = 16'b0000000000011111;
    assign weights1[56][648] = 16'b0000000000101000;
    assign weights1[56][649] = 16'b0000000000110111;
    assign weights1[56][650] = 16'b0000000001000101;
    assign weights1[56][651] = 16'b0000000001001100;
    assign weights1[56][652] = 16'b0000000000111100;
    assign weights1[56][653] = 16'b0000000001010001;
    assign weights1[56][654] = 16'b0000000001000010;
    assign weights1[56][655] = 16'b0000000000101101;
    assign weights1[56][656] = 16'b0000000000011010;
    assign weights1[56][657] = 16'b0000000000010110;
    assign weights1[56][658] = 16'b0000000000000111;
    assign weights1[56][659] = 16'b0000000000000000;
    assign weights1[56][660] = 16'b1111111111110001;
    assign weights1[56][661] = 16'b0000000000000010;
    assign weights1[56][662] = 16'b1111111111110011;
    assign weights1[56][663] = 16'b0000000000000001;
    assign weights1[56][664] = 16'b1111111111111110;
    assign weights1[56][665] = 16'b1111111111111100;
    assign weights1[56][666] = 16'b0000000000000010;
    assign weights1[56][667] = 16'b0000000000000101;
    assign weights1[56][668] = 16'b1111111111111111;
    assign weights1[56][669] = 16'b0000000000000011;
    assign weights1[56][670] = 16'b1111111111111110;
    assign weights1[56][671] = 16'b1111111111101101;
    assign weights1[56][672] = 16'b1111111111111111;
    assign weights1[56][673] = 16'b0000000000000000;
    assign weights1[56][674] = 16'b1111111111111111;
    assign weights1[56][675] = 16'b0000000000010101;
    assign weights1[56][676] = 16'b0000000000100101;
    assign weights1[56][677] = 16'b0000000000101110;
    assign weights1[56][678] = 16'b0000000000110111;
    assign weights1[56][679] = 16'b0000000000101011;
    assign weights1[56][680] = 16'b0000000000100000;
    assign weights1[56][681] = 16'b0000000000100001;
    assign weights1[56][682] = 16'b0000000000011110;
    assign weights1[56][683] = 16'b0000000000000101;
    assign weights1[56][684] = 16'b0000000000010101;
    assign weights1[56][685] = 16'b0000000000000011;
    assign weights1[56][686] = 16'b0000000000010000;
    assign weights1[56][687] = 16'b1111111111111001;
    assign weights1[56][688] = 16'b1111111111111000;
    assign weights1[56][689] = 16'b0000000000000011;
    assign weights1[56][690] = 16'b1111111111111001;
    assign weights1[56][691] = 16'b1111111111101010;
    assign weights1[56][692] = 16'b1111111111111011;
    assign weights1[56][693] = 16'b0000000000001010;
    assign weights1[56][694] = 16'b0000000000001110;
    assign weights1[56][695] = 16'b0000000000010010;
    assign weights1[56][696] = 16'b0000000000000000;
    assign weights1[56][697] = 16'b1111111111100100;
    assign weights1[56][698] = 16'b1111111111111100;
    assign weights1[56][699] = 16'b1111111111110010;
    assign weights1[56][700] = 16'b0000000000000101;
    assign weights1[56][701] = 16'b0000000000000110;
    assign weights1[56][702] = 16'b0000000000010011;
    assign weights1[56][703] = 16'b0000000000100000;
    assign weights1[56][704] = 16'b0000000000011101;
    assign weights1[56][705] = 16'b0000000000111111;
    assign weights1[56][706] = 16'b0000000000011110;
    assign weights1[56][707] = 16'b0000000000001110;
    assign weights1[56][708] = 16'b0000000000001110;
    assign weights1[56][709] = 16'b0000000000011001;
    assign weights1[56][710] = 16'b0000000000000100;
    assign weights1[56][711] = 16'b0000000000010010;
    assign weights1[56][712] = 16'b0000000000000011;
    assign weights1[56][713] = 16'b1111111111111100;
    assign weights1[56][714] = 16'b0000000000000100;
    assign weights1[56][715] = 16'b0000000000000011;
    assign weights1[56][716] = 16'b0000000000000110;
    assign weights1[56][717] = 16'b0000000000000011;
    assign weights1[56][718] = 16'b1111111111111111;
    assign weights1[56][719] = 16'b1111111111111111;
    assign weights1[56][720] = 16'b0000000000000000;
    assign weights1[56][721] = 16'b1111111111110100;
    assign weights1[56][722] = 16'b1111111111111110;
    assign weights1[56][723] = 16'b0000000000001111;
    assign weights1[56][724] = 16'b0000000000001101;
    assign weights1[56][725] = 16'b0000000000000100;
    assign weights1[56][726] = 16'b1111111111111000;
    assign weights1[56][727] = 16'b1111111111111100;
    assign weights1[56][728] = 16'b0000000000000011;
    assign weights1[56][729] = 16'b0000000000001001;
    assign weights1[56][730] = 16'b0000000000001111;
    assign weights1[56][731] = 16'b0000000000011010;
    assign weights1[56][732] = 16'b0000000000001000;
    assign weights1[56][733] = 16'b0000000000011111;
    assign weights1[56][734] = 16'b0000000000010101;
    assign weights1[56][735] = 16'b0000000000000101;
    assign weights1[56][736] = 16'b0000000000011011;
    assign weights1[56][737] = 16'b0000000000001110;
    assign weights1[56][738] = 16'b0000000000000111;
    assign weights1[56][739] = 16'b0000000000000110;
    assign weights1[56][740] = 16'b0000000000001001;
    assign weights1[56][741] = 16'b0000000000010000;
    assign weights1[56][742] = 16'b0000000000000110;
    assign weights1[56][743] = 16'b1111111111111000;
    assign weights1[56][744] = 16'b0000000000000000;
    assign weights1[56][745] = 16'b1111111111101110;
    assign weights1[56][746] = 16'b0000000000000000;
    assign weights1[56][747] = 16'b1111111111111010;
    assign weights1[56][748] = 16'b1111111111111011;
    assign weights1[56][749] = 16'b0000000000000010;
    assign weights1[56][750] = 16'b1111111111111000;
    assign weights1[56][751] = 16'b1111111111110111;
    assign weights1[56][752] = 16'b1111111111111111;
    assign weights1[56][753] = 16'b0000000000000011;
    assign weights1[56][754] = 16'b1111111111111001;
    assign weights1[56][755] = 16'b0000000000000010;
    assign weights1[56][756] = 16'b0000000000001010;
    assign weights1[56][757] = 16'b0000000000010100;
    assign weights1[56][758] = 16'b0000000000010100;
    assign weights1[56][759] = 16'b0000000000001001;
    assign weights1[56][760] = 16'b0000000000011010;
    assign weights1[56][761] = 16'b0000000000011011;
    assign weights1[56][762] = 16'b0000000000010000;
    assign weights1[56][763] = 16'b0000000000000011;
    assign weights1[56][764] = 16'b0000000000001100;
    assign weights1[56][765] = 16'b0000000000000101;
    assign weights1[56][766] = 16'b0000000000000011;
    assign weights1[56][767] = 16'b0000000000000000;
    assign weights1[56][768] = 16'b1111111111111010;
    assign weights1[56][769] = 16'b1111111111110011;
    assign weights1[56][770] = 16'b1111111111110111;
    assign weights1[56][771] = 16'b1111111111110100;
    assign weights1[56][772] = 16'b0000000000000100;
    assign weights1[56][773] = 16'b1111111111111110;
    assign weights1[56][774] = 16'b1111111111111001;
    assign weights1[56][775] = 16'b1111111111110011;
    assign weights1[56][776] = 16'b1111111111110111;
    assign weights1[56][777] = 16'b1111111111110110;
    assign weights1[56][778] = 16'b0000000000000001;
    assign weights1[56][779] = 16'b1111111111111011;
    assign weights1[56][780] = 16'b1111111111110110;
    assign weights1[56][781] = 16'b0000000000000001;
    assign weights1[56][782] = 16'b1111111111111011;
    assign weights1[56][783] = 16'b0000000000000000;
    assign weights1[57][0] = 16'b1111111111111111;
    assign weights1[57][1] = 16'b0000000000000000;
    assign weights1[57][2] = 16'b0000000000000000;
    assign weights1[57][3] = 16'b0000000000000001;
    assign weights1[57][4] = 16'b0000000000000011;
    assign weights1[57][5] = 16'b0000000000001111;
    assign weights1[57][6] = 16'b0000000000011111;
    assign weights1[57][7] = 16'b0000000000101000;
    assign weights1[57][8] = 16'b0000000000100010;
    assign weights1[57][9] = 16'b0000000000011110;
    assign weights1[57][10] = 16'b0000000000001000;
    assign weights1[57][11] = 16'b1111111111001110;
    assign weights1[57][12] = 16'b1111111110100111;
    assign weights1[57][13] = 16'b1111111110011001;
    assign weights1[57][14] = 16'b1111111110011111;
    assign weights1[57][15] = 16'b1111111110111111;
    assign weights1[57][16] = 16'b1111111111010011;
    assign weights1[57][17] = 16'b1111111111110110;
    assign weights1[57][18] = 16'b0000000000000011;
    assign weights1[57][19] = 16'b0000000000001101;
    assign weights1[57][20] = 16'b0000000000001110;
    assign weights1[57][21] = 16'b0000000000010010;
    assign weights1[57][22] = 16'b0000000000000001;
    assign weights1[57][23] = 16'b1111111111111010;
    assign weights1[57][24] = 16'b1111111111110100;
    assign weights1[57][25] = 16'b1111111111111000;
    assign weights1[57][26] = 16'b1111111111111001;
    assign weights1[57][27] = 16'b0000000000000001;
    assign weights1[57][28] = 16'b1111111111111111;
    assign weights1[57][29] = 16'b0000000000000011;
    assign weights1[57][30] = 16'b0000000000000111;
    assign weights1[57][31] = 16'b0000000000000100;
    assign weights1[57][32] = 16'b0000000000001011;
    assign weights1[57][33] = 16'b0000000000001110;
    assign weights1[57][34] = 16'b0000000000100100;
    assign weights1[57][35] = 16'b0000000000101111;
    assign weights1[57][36] = 16'b0000000000011011;
    assign weights1[57][37] = 16'b0000000000010100;
    assign weights1[57][38] = 16'b1111111111110101;
    assign weights1[57][39] = 16'b1111111111001010;
    assign weights1[57][40] = 16'b1111111110001000;
    assign weights1[57][41] = 16'b1111111110000001;
    assign weights1[57][42] = 16'b1111111110101011;
    assign weights1[57][43] = 16'b1111111111100100;
    assign weights1[57][44] = 16'b1111111111101011;
    assign weights1[57][45] = 16'b1111111111111101;
    assign weights1[57][46] = 16'b0000000000001111;
    assign weights1[57][47] = 16'b0000000000010101;
    assign weights1[57][48] = 16'b0000000000010110;
    assign weights1[57][49] = 16'b0000000000010001;
    assign weights1[57][50] = 16'b0000000000000111;
    assign weights1[57][51] = 16'b1111111111111011;
    assign weights1[57][52] = 16'b1111111111101111;
    assign weights1[57][53] = 16'b1111111111100101;
    assign weights1[57][54] = 16'b1111111111110011;
    assign weights1[57][55] = 16'b1111111111111010;
    assign weights1[57][56] = 16'b1111111111111111;
    assign weights1[57][57] = 16'b0000000000000011;
    assign weights1[57][58] = 16'b0000000000000000;
    assign weights1[57][59] = 16'b1111111111111111;
    assign weights1[57][60] = 16'b0000000000000001;
    assign weights1[57][61] = 16'b0000000000010100;
    assign weights1[57][62] = 16'b0000000000100010;
    assign weights1[57][63] = 16'b0000000000110110;
    assign weights1[57][64] = 16'b0000000000011011;
    assign weights1[57][65] = 16'b0000000000001110;
    assign weights1[57][66] = 16'b1111111111100010;
    assign weights1[57][67] = 16'b1111111110011011;
    assign weights1[57][68] = 16'b1111111101101101;
    assign weights1[57][69] = 16'b1111111110001100;
    assign weights1[57][70] = 16'b1111111110111100;
    assign weights1[57][71] = 16'b1111111111110010;
    assign weights1[57][72] = 16'b0000000000011011;
    assign weights1[57][73] = 16'b0000000000001111;
    assign weights1[57][74] = 16'b0000000000011111;
    assign weights1[57][75] = 16'b0000000000010101;
    assign weights1[57][76] = 16'b0000000000010001;
    assign weights1[57][77] = 16'b1111111111111110;
    assign weights1[57][78] = 16'b1111111111111000;
    assign weights1[57][79] = 16'b1111111111011101;
    assign weights1[57][80] = 16'b1111111111010011;
    assign weights1[57][81] = 16'b1111111111100010;
    assign weights1[57][82] = 16'b1111111111100110;
    assign weights1[57][83] = 16'b1111111111101111;
    assign weights1[57][84] = 16'b0000000000000011;
    assign weights1[57][85] = 16'b0000000000000011;
    assign weights1[57][86] = 16'b1111111111111001;
    assign weights1[57][87] = 16'b0000000000000001;
    assign weights1[57][88] = 16'b0000000000000110;
    assign weights1[57][89] = 16'b0000000000011110;
    assign weights1[57][90] = 16'b0000000000011101;
    assign weights1[57][91] = 16'b0000000000101010;
    assign weights1[57][92] = 16'b0000000000010101;
    assign weights1[57][93] = 16'b0000000000010101;
    assign weights1[57][94] = 16'b1111111111110000;
    assign weights1[57][95] = 16'b1111111110000011;
    assign weights1[57][96] = 16'b1111111101010011;
    assign weights1[57][97] = 16'b1111111101100110;
    assign weights1[57][98] = 16'b1111111110110001;
    assign weights1[57][99] = 16'b1111111111110111;
    assign weights1[57][100] = 16'b1111111111101011;
    assign weights1[57][101] = 16'b0000000000000011;
    assign weights1[57][102] = 16'b0000000000110100;
    assign weights1[57][103] = 16'b0000000000101010;
    assign weights1[57][104] = 16'b0000000000011001;
    assign weights1[57][105] = 16'b0000000000001101;
    assign weights1[57][106] = 16'b1111111111101111;
    assign weights1[57][107] = 16'b1111111111000111;
    assign weights1[57][108] = 16'b1111111111000011;
    assign weights1[57][109] = 16'b1111111111011000;
    assign weights1[57][110] = 16'b1111111111100101;
    assign weights1[57][111] = 16'b1111111111110110;
    assign weights1[57][112] = 16'b0000000000000001;
    assign weights1[57][113] = 16'b1111111111111100;
    assign weights1[57][114] = 16'b1111111111111110;
    assign weights1[57][115] = 16'b0000000000000110;
    assign weights1[57][116] = 16'b0000000000001110;
    assign weights1[57][117] = 16'b0000000000101010;
    assign weights1[57][118] = 16'b0000000000010010;
    assign weights1[57][119] = 16'b0000000000100001;
    assign weights1[57][120] = 16'b0000000000100000;
    assign weights1[57][121] = 16'b0000000000100000;
    assign weights1[57][122] = 16'b1111111111100011;
    assign weights1[57][123] = 16'b1111111101100101;
    assign weights1[57][124] = 16'b1111111100111110;
    assign weights1[57][125] = 16'b1111111101001101;
    assign weights1[57][126] = 16'b1111111111001111;
    assign weights1[57][127] = 16'b0000000000001111;
    assign weights1[57][128] = 16'b0000000000001011;
    assign weights1[57][129] = 16'b0000000000011111;
    assign weights1[57][130] = 16'b0000000000010010;
    assign weights1[57][131] = 16'b0000000000001100;
    assign weights1[57][132] = 16'b0000000000001111;
    assign weights1[57][133] = 16'b1111111111011110;
    assign weights1[57][134] = 16'b1111111111001110;
    assign weights1[57][135] = 16'b1111111110111001;
    assign weights1[57][136] = 16'b1111111110111000;
    assign weights1[57][137] = 16'b1111111111011001;
    assign weights1[57][138] = 16'b1111111111101101;
    assign weights1[57][139] = 16'b1111111111111100;
    assign weights1[57][140] = 16'b1111111111111100;
    assign weights1[57][141] = 16'b1111111111111001;
    assign weights1[57][142] = 16'b1111111111110111;
    assign weights1[57][143] = 16'b1111111111110101;
    assign weights1[57][144] = 16'b0000000000000011;
    assign weights1[57][145] = 16'b0000000000011110;
    assign weights1[57][146] = 16'b0000000000100011;
    assign weights1[57][147] = 16'b0000000000111000;
    assign weights1[57][148] = 16'b0000000000100100;
    assign weights1[57][149] = 16'b0000000000011111;
    assign weights1[57][150] = 16'b1111111111010011;
    assign weights1[57][151] = 16'b1111111101001000;
    assign weights1[57][152] = 16'b1111111100101000;
    assign weights1[57][153] = 16'b1111111101110101;
    assign weights1[57][154] = 16'b0000000000111111;
    assign weights1[57][155] = 16'b0000000000111100;
    assign weights1[57][156] = 16'b0000000000011001;
    assign weights1[57][157] = 16'b0000000000110101;
    assign weights1[57][158] = 16'b0000000000101101;
    assign weights1[57][159] = 16'b0000000000011000;
    assign weights1[57][160] = 16'b1111111111110010;
    assign weights1[57][161] = 16'b1111111111001000;
    assign weights1[57][162] = 16'b1111111110110010;
    assign weights1[57][163] = 16'b1111111110101111;
    assign weights1[57][164] = 16'b1111111111000110;
    assign weights1[57][165] = 16'b1111111111011101;
    assign weights1[57][166] = 16'b1111111111101011;
    assign weights1[57][167] = 16'b1111111111110011;
    assign weights1[57][168] = 16'b1111111111110100;
    assign weights1[57][169] = 16'b1111111111110010;
    assign weights1[57][170] = 16'b1111111111101000;
    assign weights1[57][171] = 16'b1111111111110111;
    assign weights1[57][172] = 16'b1111111111111011;
    assign weights1[57][173] = 16'b0000000000000010;
    assign weights1[57][174] = 16'b0000000000011101;
    assign weights1[57][175] = 16'b0000000000100011;
    assign weights1[57][176] = 16'b0000000000101100;
    assign weights1[57][177] = 16'b0000000000111011;
    assign weights1[57][178] = 16'b1111111110110001;
    assign weights1[57][179] = 16'b1111111101001111;
    assign weights1[57][180] = 16'b1111111100111001;
    assign weights1[57][181] = 16'b1111111111000000;
    assign weights1[57][182] = 16'b0000000000100000;
    assign weights1[57][183] = 16'b0000000000111010;
    assign weights1[57][184] = 16'b0000000000011111;
    assign weights1[57][185] = 16'b0000000000010111;
    assign weights1[57][186] = 16'b0000000000001101;
    assign weights1[57][187] = 16'b0000000000010011;
    assign weights1[57][188] = 16'b1111111111001110;
    assign weights1[57][189] = 16'b1111111110101100;
    assign weights1[57][190] = 16'b1111111110010001;
    assign weights1[57][191] = 16'b1111111110010110;
    assign weights1[57][192] = 16'b1111111111001011;
    assign weights1[57][193] = 16'b1111111111100001;
    assign weights1[57][194] = 16'b1111111111111010;
    assign weights1[57][195] = 16'b0000000000000100;
    assign weights1[57][196] = 16'b1111111111110010;
    assign weights1[57][197] = 16'b1111111111011111;
    assign weights1[57][198] = 16'b1111111111011101;
    assign weights1[57][199] = 16'b1111111111110111;
    assign weights1[57][200] = 16'b1111111111100101;
    assign weights1[57][201] = 16'b1111111111111111;
    assign weights1[57][202] = 16'b0000000000010101;
    assign weights1[57][203] = 16'b0000000000011001;
    assign weights1[57][204] = 16'b0000000000101101;
    assign weights1[57][205] = 16'b0000000000111110;
    assign weights1[57][206] = 16'b1111111111000100;
    assign weights1[57][207] = 16'b1111111100100101;
    assign weights1[57][208] = 16'b1111111101100110;
    assign weights1[57][209] = 16'b1111111111110101;
    assign weights1[57][210] = 16'b0000000000100101;
    assign weights1[57][211] = 16'b0000000000101101;
    assign weights1[57][212] = 16'b0000000000011111;
    assign weights1[57][213] = 16'b0000000000101011;
    assign weights1[57][214] = 16'b0000000000001001;
    assign weights1[57][215] = 16'b1111111111111101;
    assign weights1[57][216] = 16'b1111111111011001;
    assign weights1[57][217] = 16'b1111111110010111;
    assign weights1[57][218] = 16'b1111111110011010;
    assign weights1[57][219] = 16'b1111111111000101;
    assign weights1[57][220] = 16'b1111111111111100;
    assign weights1[57][221] = 16'b1111111111111101;
    assign weights1[57][222] = 16'b0000000000010000;
    assign weights1[57][223] = 16'b0000000000001111;
    assign weights1[57][224] = 16'b1111111111110110;
    assign weights1[57][225] = 16'b1111111111101011;
    assign weights1[57][226] = 16'b1111111111101011;
    assign weights1[57][227] = 16'b1111111111111000;
    assign weights1[57][228] = 16'b0000000000001100;
    assign weights1[57][229] = 16'b0000000000001000;
    assign weights1[57][230] = 16'b0000000000010000;
    assign weights1[57][231] = 16'b0000000000011110;
    assign weights1[57][232] = 16'b0000000000111000;
    assign weights1[57][233] = 16'b0000000000101100;
    assign weights1[57][234] = 16'b1111111111000110;
    assign weights1[57][235] = 16'b1111111101001000;
    assign weights1[57][236] = 16'b1111111110111100;
    assign weights1[57][237] = 16'b1111111111110000;
    assign weights1[57][238] = 16'b0000000000001101;
    assign weights1[57][239] = 16'b0000000000111010;
    assign weights1[57][240] = 16'b0000000000011101;
    assign weights1[57][241] = 16'b0000000000010010;
    assign weights1[57][242] = 16'b0000000000000010;
    assign weights1[57][243] = 16'b1111111111011110;
    assign weights1[57][244] = 16'b1111111110111001;
    assign weights1[57][245] = 16'b1111111110010011;
    assign weights1[57][246] = 16'b1111111111001110;
    assign weights1[57][247] = 16'b0000000000001101;
    assign weights1[57][248] = 16'b0000000000010100;
    assign weights1[57][249] = 16'b0000000000010001;
    assign weights1[57][250] = 16'b0000000000100010;
    assign weights1[57][251] = 16'b0000000000011111;
    assign weights1[57][252] = 16'b1111111111110111;
    assign weights1[57][253] = 16'b1111111111101100;
    assign weights1[57][254] = 16'b1111111111110100;
    assign weights1[57][255] = 16'b1111111111101001;
    assign weights1[57][256] = 16'b0000000000000010;
    assign weights1[57][257] = 16'b0000000000000001;
    assign weights1[57][258] = 16'b0000000000000100;
    assign weights1[57][259] = 16'b0000000000010101;
    assign weights1[57][260] = 16'b0000000000001110;
    assign weights1[57][261] = 16'b0000000000110110;
    assign weights1[57][262] = 16'b1111111111001001;
    assign weights1[57][263] = 16'b1111111110100100;
    assign weights1[57][264] = 16'b1111111111000100;
    assign weights1[57][265] = 16'b1111111111111100;
    assign weights1[57][266] = 16'b0000000000011011;
    assign weights1[57][267] = 16'b0000000000011011;
    assign weights1[57][268] = 16'b0000000000010011;
    assign weights1[57][269] = 16'b0000000000011111;
    assign weights1[57][270] = 16'b1111111111101011;
    assign weights1[57][271] = 16'b1111111111011110;
    assign weights1[57][272] = 16'b1111111110101110;
    assign weights1[57][273] = 16'b1111111110110001;
    assign weights1[57][274] = 16'b0000000000001001;
    assign weights1[57][275] = 16'b0000000000100100;
    assign weights1[57][276] = 16'b0000000000011110;
    assign weights1[57][277] = 16'b0000000000010000;
    assign weights1[57][278] = 16'b0000000000011110;
    assign weights1[57][279] = 16'b0000000000001110;
    assign weights1[57][280] = 16'b1111111111110111;
    assign weights1[57][281] = 16'b1111111111110010;
    assign weights1[57][282] = 16'b1111111111111011;
    assign weights1[57][283] = 16'b0000000000001001;
    assign weights1[57][284] = 16'b0000000000001100;
    assign weights1[57][285] = 16'b1111111111111100;
    assign weights1[57][286] = 16'b1111111111111100;
    assign weights1[57][287] = 16'b0000000000010010;
    assign weights1[57][288] = 16'b0000000000010011;
    assign weights1[57][289] = 16'b0000000000100000;
    assign weights1[57][290] = 16'b1111111111011011;
    assign weights1[57][291] = 16'b1111111111000100;
    assign weights1[57][292] = 16'b1111111111100101;
    assign weights1[57][293] = 16'b0000000000000001;
    assign weights1[57][294] = 16'b0000000000000100;
    assign weights1[57][295] = 16'b0000000000100001;
    assign weights1[57][296] = 16'b0000000000001111;
    assign weights1[57][297] = 16'b0000000000000010;
    assign weights1[57][298] = 16'b1111111111101101;
    assign weights1[57][299] = 16'b1111111111010100;
    assign weights1[57][300] = 16'b1111111111001011;
    assign weights1[57][301] = 16'b1111111111101000;
    assign weights1[57][302] = 16'b0000000000100101;
    assign weights1[57][303] = 16'b0000000000010111;
    assign weights1[57][304] = 16'b0000000000011111;
    assign weights1[57][305] = 16'b0000000000101000;
    assign weights1[57][306] = 16'b0000000000001111;
    assign weights1[57][307] = 16'b0000000000001001;
    assign weights1[57][308] = 16'b1111111111110111;
    assign weights1[57][309] = 16'b1111111111110110;
    assign weights1[57][310] = 16'b1111111111101001;
    assign weights1[57][311] = 16'b1111111111111001;
    assign weights1[57][312] = 16'b1111111111110100;
    assign weights1[57][313] = 16'b1111111111110100;
    assign weights1[57][314] = 16'b0000000000010001;
    assign weights1[57][315] = 16'b1111111111110001;
    assign weights1[57][316] = 16'b0000000000001101;
    assign weights1[57][317] = 16'b0000000000010110;
    assign weights1[57][318] = 16'b1111111111101111;
    assign weights1[57][319] = 16'b1111111111100001;
    assign weights1[57][320] = 16'b1111111111100010;
    assign weights1[57][321] = 16'b0000000000001000;
    assign weights1[57][322] = 16'b0000000000001000;
    assign weights1[57][323] = 16'b1111111111111011;
    assign weights1[57][324] = 16'b1111111111111011;
    assign weights1[57][325] = 16'b1111111111111010;
    assign weights1[57][326] = 16'b1111111111111110;
    assign weights1[57][327] = 16'b1111111111000010;
    assign weights1[57][328] = 16'b1111111111101100;
    assign weights1[57][329] = 16'b1111111111111101;
    assign weights1[57][330] = 16'b0000000000010010;
    assign weights1[57][331] = 16'b0000000000010010;
    assign weights1[57][332] = 16'b0000000000000111;
    assign weights1[57][333] = 16'b0000000000001100;
    assign weights1[57][334] = 16'b1111111111111111;
    assign weights1[57][335] = 16'b0000000000001001;
    assign weights1[57][336] = 16'b1111111111110100;
    assign weights1[57][337] = 16'b1111111111110010;
    assign weights1[57][338] = 16'b0000000000000111;
    assign weights1[57][339] = 16'b0000000000000000;
    assign weights1[57][340] = 16'b1111111111111100;
    assign weights1[57][341] = 16'b0000000000000100;
    assign weights1[57][342] = 16'b0000000000001010;
    assign weights1[57][343] = 16'b0000000000000101;
    assign weights1[57][344] = 16'b0000000000010101;
    assign weights1[57][345] = 16'b0000000000001010;
    assign weights1[57][346] = 16'b1111111111111100;
    assign weights1[57][347] = 16'b1111111111100100;
    assign weights1[57][348] = 16'b1111111111110001;
    assign weights1[57][349] = 16'b0000000000001111;
    assign weights1[57][350] = 16'b0000000000000000;
    assign weights1[57][351] = 16'b0000000000000011;
    assign weights1[57][352] = 16'b0000000000010010;
    assign weights1[57][353] = 16'b1111111111110001;
    assign weights1[57][354] = 16'b1111111111101111;
    assign weights1[57][355] = 16'b1111111111010001;
    assign weights1[57][356] = 16'b1111111111110100;
    assign weights1[57][357] = 16'b0000000000010101;
    assign weights1[57][358] = 16'b0000000000010111;
    assign weights1[57][359] = 16'b0000000000000011;
    assign weights1[57][360] = 16'b0000000000001010;
    assign weights1[57][361] = 16'b0000000000001000;
    assign weights1[57][362] = 16'b0000000000000110;
    assign weights1[57][363] = 16'b0000000000001111;
    assign weights1[57][364] = 16'b1111111111110011;
    assign weights1[57][365] = 16'b1111111111111100;
    assign weights1[57][366] = 16'b1111111111111010;
    assign weights1[57][367] = 16'b1111111111110010;
    assign weights1[57][368] = 16'b0000000000000001;
    assign weights1[57][369] = 16'b0000000000001000;
    assign weights1[57][370] = 16'b0000000000000000;
    assign weights1[57][371] = 16'b0000000000000100;
    assign weights1[57][372] = 16'b0000000000000010;
    assign weights1[57][373] = 16'b0000000000010000;
    assign weights1[57][374] = 16'b0000000000001001;
    assign weights1[57][375] = 16'b0000000000000001;
    assign weights1[57][376] = 16'b0000000000000011;
    assign weights1[57][377] = 16'b1111111111111100;
    assign weights1[57][378] = 16'b1111111111110010;
    assign weights1[57][379] = 16'b0000000000000000;
    assign weights1[57][380] = 16'b1111111111110011;
    assign weights1[57][381] = 16'b1111111111100010;
    assign weights1[57][382] = 16'b0000000000000000;
    assign weights1[57][383] = 16'b1111111111101110;
    assign weights1[57][384] = 16'b0000000000000111;
    assign weights1[57][385] = 16'b0000000000001001;
    assign weights1[57][386] = 16'b0000000000010111;
    assign weights1[57][387] = 16'b0000000000001100;
    assign weights1[57][388] = 16'b1111111111110010;
    assign weights1[57][389] = 16'b0000000000000000;
    assign weights1[57][390] = 16'b0000000000001000;
    assign weights1[57][391] = 16'b0000000000010001;
    assign weights1[57][392] = 16'b1111111111111011;
    assign weights1[57][393] = 16'b1111111111110011;
    assign weights1[57][394] = 16'b1111111111101010;
    assign weights1[57][395] = 16'b1111111111111100;
    assign weights1[57][396] = 16'b1111111111101101;
    assign weights1[57][397] = 16'b0000000000001111;
    assign weights1[57][398] = 16'b1111111111111011;
    assign weights1[57][399] = 16'b0000000000001010;
    assign weights1[57][400] = 16'b0000000000001110;
    assign weights1[57][401] = 16'b0000000000000111;
    assign weights1[57][402] = 16'b0000000000000011;
    assign weights1[57][403] = 16'b0000000000001111;
    assign weights1[57][404] = 16'b1111111111111101;
    assign weights1[57][405] = 16'b0000000000000100;
    assign weights1[57][406] = 16'b0000000000000101;
    assign weights1[57][407] = 16'b1111111111110110;
    assign weights1[57][408] = 16'b1111111111111010;
    assign weights1[57][409] = 16'b0000000000010000;
    assign weights1[57][410] = 16'b0000000000000001;
    assign weights1[57][411] = 16'b0000000000001101;
    assign weights1[57][412] = 16'b0000000000001010;
    assign weights1[57][413] = 16'b0000000000000110;
    assign weights1[57][414] = 16'b0000000000000101;
    assign weights1[57][415] = 16'b1111111111111000;
    assign weights1[57][416] = 16'b0000000000001110;
    assign weights1[57][417] = 16'b0000000000000101;
    assign weights1[57][418] = 16'b0000000000000101;
    assign weights1[57][419] = 16'b1111111111111110;
    assign weights1[57][420] = 16'b1111111111110100;
    assign weights1[57][421] = 16'b1111111111110011;
    assign weights1[57][422] = 16'b1111111111111101;
    assign weights1[57][423] = 16'b1111111111110010;
    assign weights1[57][424] = 16'b1111111111111011;
    assign weights1[57][425] = 16'b0000000000001010;
    assign weights1[57][426] = 16'b0000000000000000;
    assign weights1[57][427] = 16'b0000000000010110;
    assign weights1[57][428] = 16'b0000000000010010;
    assign weights1[57][429] = 16'b0000000000010100;
    assign weights1[57][430] = 16'b1111111111111101;
    assign weights1[57][431] = 16'b0000000000010101;
    assign weights1[57][432] = 16'b1111111111110110;
    assign weights1[57][433] = 16'b1111111111110000;
    assign weights1[57][434] = 16'b0000000000000001;
    assign weights1[57][435] = 16'b1111111111111010;
    assign weights1[57][436] = 16'b1111111111100010;
    assign weights1[57][437] = 16'b0000000000001011;
    assign weights1[57][438] = 16'b1111111111111101;
    assign weights1[57][439] = 16'b0000000000001000;
    assign weights1[57][440] = 16'b0000000000010011;
    assign weights1[57][441] = 16'b0000000000010001;
    assign weights1[57][442] = 16'b0000000000000110;
    assign weights1[57][443] = 16'b0000000000001010;
    assign weights1[57][444] = 16'b0000000000000111;
    assign weights1[57][445] = 16'b1111111111111011;
    assign weights1[57][446] = 16'b0000000000000100;
    assign weights1[57][447] = 16'b1111111111111110;
    assign weights1[57][448] = 16'b1111111111111000;
    assign weights1[57][449] = 16'b1111111111111011;
    assign weights1[57][450] = 16'b0000000000000101;
    assign weights1[57][451] = 16'b1111111111111111;
    assign weights1[57][452] = 16'b0000000000000111;
    assign weights1[57][453] = 16'b0000000000001101;
    assign weights1[57][454] = 16'b0000000000001110;
    assign weights1[57][455] = 16'b0000000000000010;
    assign weights1[57][456] = 16'b1111111111111010;
    assign weights1[57][457] = 16'b0000000000001001;
    assign weights1[57][458] = 16'b0000000000001000;
    assign weights1[57][459] = 16'b1111111111110101;
    assign weights1[57][460] = 16'b0000000000010110;
    assign weights1[57][461] = 16'b0000000000001001;
    assign weights1[57][462] = 16'b0000000000000000;
    assign weights1[57][463] = 16'b1111111111110011;
    assign weights1[57][464] = 16'b0000000000000001;
    assign weights1[57][465] = 16'b0000000000000110;
    assign weights1[57][466] = 16'b1111111111111001;
    assign weights1[57][467] = 16'b0000000000001000;
    assign weights1[57][468] = 16'b0000000000001000;
    assign weights1[57][469] = 16'b0000000000001100;
    assign weights1[57][470] = 16'b0000000000000000;
    assign weights1[57][471] = 16'b0000000000000101;
    assign weights1[57][472] = 16'b1111111111111111;
    assign weights1[57][473] = 16'b0000000000001001;
    assign weights1[57][474] = 16'b0000000000010100;
    assign weights1[57][475] = 16'b1111111111111011;
    assign weights1[57][476] = 16'b1111111111111101;
    assign weights1[57][477] = 16'b0000000000001111;
    assign weights1[57][478] = 16'b0000000000011010;
    assign weights1[57][479] = 16'b0000000000010011;
    assign weights1[57][480] = 16'b0000000000011011;
    assign weights1[57][481] = 16'b0000000000001000;
    assign weights1[57][482] = 16'b0000000000000101;
    assign weights1[57][483] = 16'b0000000000000100;
    assign weights1[57][484] = 16'b0000000000001011;
    assign weights1[57][485] = 16'b1111111111111110;
    assign weights1[57][486] = 16'b1111111111111001;
    assign weights1[57][487] = 16'b0000000000001000;
    assign weights1[57][488] = 16'b1111111111101101;
    assign weights1[57][489] = 16'b0000000000000000;
    assign weights1[57][490] = 16'b0000000000000000;
    assign weights1[57][491] = 16'b1111111111110000;
    assign weights1[57][492] = 16'b0000000000000000;
    assign weights1[57][493] = 16'b1111111111110010;
    assign weights1[57][494] = 16'b0000000000000011;
    assign weights1[57][495] = 16'b0000000000001000;
    assign weights1[57][496] = 16'b0000000000000111;
    assign weights1[57][497] = 16'b1111111111110101;
    assign weights1[57][498] = 16'b0000000000000011;
    assign weights1[57][499] = 16'b0000000000001000;
    assign weights1[57][500] = 16'b1111111111110101;
    assign weights1[57][501] = 16'b0000000000001000;
    assign weights1[57][502] = 16'b0000000000010011;
    assign weights1[57][503] = 16'b0000000000010110;
    assign weights1[57][504] = 16'b0000000000000110;
    assign weights1[57][505] = 16'b0000000000001110;
    assign weights1[57][506] = 16'b0000000000000101;
    assign weights1[57][507] = 16'b0000000000010100;
    assign weights1[57][508] = 16'b1111111111111111;
    assign weights1[57][509] = 16'b1111111111101100;
    assign weights1[57][510] = 16'b0000000000000101;
    assign weights1[57][511] = 16'b1111111111111101;
    assign weights1[57][512] = 16'b1111111111111000;
    assign weights1[57][513] = 16'b0000000000011000;
    assign weights1[57][514] = 16'b1111111111111111;
    assign weights1[57][515] = 16'b0000000000000001;
    assign weights1[57][516] = 16'b0000000000000011;
    assign weights1[57][517] = 16'b1111111111111101;
    assign weights1[57][518] = 16'b1111111111110110;
    assign weights1[57][519] = 16'b0000000000000100;
    assign weights1[57][520] = 16'b1111111111111111;
    assign weights1[57][521] = 16'b0000000000000000;
    assign weights1[57][522] = 16'b0000000000001001;
    assign weights1[57][523] = 16'b0000000000000000;
    assign weights1[57][524] = 16'b0000000000000011;
    assign weights1[57][525] = 16'b0000000000011000;
    assign weights1[57][526] = 16'b1111111111110101;
    assign weights1[57][527] = 16'b0000000000010010;
    assign weights1[57][528] = 16'b1111111111110010;
    assign weights1[57][529] = 16'b0000000000001001;
    assign weights1[57][530] = 16'b0000000000001110;
    assign weights1[57][531] = 16'b0000000000010100;
    assign weights1[57][532] = 16'b0000000000000100;
    assign weights1[57][533] = 16'b0000000000001011;
    assign weights1[57][534] = 16'b0000000000001001;
    assign weights1[57][535] = 16'b1111111111110001;
    assign weights1[57][536] = 16'b0000000000010000;
    assign weights1[57][537] = 16'b0000000000010101;
    assign weights1[57][538] = 16'b0000000000000100;
    assign weights1[57][539] = 16'b1111111111110100;
    assign weights1[57][540] = 16'b1111111111110000;
    assign weights1[57][541] = 16'b0000000000000110;
    assign weights1[57][542] = 16'b1111111111101011;
    assign weights1[57][543] = 16'b0000000000000010;
    assign weights1[57][544] = 16'b0000000000001001;
    assign weights1[57][545] = 16'b0000000000000010;
    assign weights1[57][546] = 16'b1111111111110010;
    assign weights1[57][547] = 16'b0000000000010111;
    assign weights1[57][548] = 16'b1111111111111101;
    assign weights1[57][549] = 16'b1111111111110100;
    assign weights1[57][550] = 16'b0000000000001110;
    assign weights1[57][551] = 16'b1111111111110110;
    assign weights1[57][552] = 16'b0000000000000111;
    assign weights1[57][553] = 16'b1111111111111001;
    assign weights1[57][554] = 16'b1111111111110001;
    assign weights1[57][555] = 16'b0000000000010110;
    assign weights1[57][556] = 16'b0000000000000000;
    assign weights1[57][557] = 16'b0000000000001011;
    assign weights1[57][558] = 16'b0000000000001010;
    assign weights1[57][559] = 16'b0000000000001101;
    assign weights1[57][560] = 16'b0000000000001010;
    assign weights1[57][561] = 16'b1111111111110001;
    assign weights1[57][562] = 16'b0000000000000111;
    assign weights1[57][563] = 16'b1111111111111100;
    assign weights1[57][564] = 16'b1111111111111111;
    assign weights1[57][565] = 16'b1111111111111010;
    assign weights1[57][566] = 16'b1111111111111100;
    assign weights1[57][567] = 16'b1111111111100111;
    assign weights1[57][568] = 16'b0000000000001110;
    assign weights1[57][569] = 16'b1111111111111000;
    assign weights1[57][570] = 16'b1111111111110001;
    assign weights1[57][571] = 16'b0000000000001110;
    assign weights1[57][572] = 16'b1111111111111010;
    assign weights1[57][573] = 16'b1111111111101001;
    assign weights1[57][574] = 16'b1111111111111111;
    assign weights1[57][575] = 16'b1111111111111110;
    assign weights1[57][576] = 16'b1111111111111111;
    assign weights1[57][577] = 16'b0000000000001101;
    assign weights1[57][578] = 16'b0000000000001101;
    assign weights1[57][579] = 16'b1111111111111010;
    assign weights1[57][580] = 16'b0000000000010100;
    assign weights1[57][581] = 16'b0000000000001111;
    assign weights1[57][582] = 16'b1111111111110100;
    assign weights1[57][583] = 16'b1111111111111111;
    assign weights1[57][584] = 16'b1111111111111111;
    assign weights1[57][585] = 16'b0000000000010100;
    assign weights1[57][586] = 16'b0000000000001001;
    assign weights1[57][587] = 16'b0000000000000101;
    assign weights1[57][588] = 16'b0000000000010011;
    assign weights1[57][589] = 16'b0000000000000100;
    assign weights1[57][590] = 16'b0000000000000101;
    assign weights1[57][591] = 16'b0000000000000000;
    assign weights1[57][592] = 16'b0000000000001110;
    assign weights1[57][593] = 16'b0000000000000010;
    assign weights1[57][594] = 16'b1111111111101100;
    assign weights1[57][595] = 16'b0000000000001001;
    assign weights1[57][596] = 16'b1111111111111000;
    assign weights1[57][597] = 16'b1111111111110111;
    assign weights1[57][598] = 16'b1111111111110011;
    assign weights1[57][599] = 16'b0000000000001110;
    assign weights1[57][600] = 16'b0000000000001010;
    assign weights1[57][601] = 16'b0000000000000100;
    assign weights1[57][602] = 16'b1111111111111110;
    assign weights1[57][603] = 16'b0000000000000101;
    assign weights1[57][604] = 16'b1111111111111111;
    assign weights1[57][605] = 16'b1111111111110111;
    assign weights1[57][606] = 16'b1111111111111110;
    assign weights1[57][607] = 16'b1111111111111101;
    assign weights1[57][608] = 16'b1111111111110110;
    assign weights1[57][609] = 16'b0000000000000010;
    assign weights1[57][610] = 16'b0000000000001101;
    assign weights1[57][611] = 16'b0000000000000100;
    assign weights1[57][612] = 16'b0000000000001111;
    assign weights1[57][613] = 16'b0000000000000100;
    assign weights1[57][614] = 16'b0000000000000000;
    assign weights1[57][615] = 16'b1111111111111011;
    assign weights1[57][616] = 16'b0000000000000111;
    assign weights1[57][617] = 16'b0000000000000100;
    assign weights1[57][618] = 16'b0000000000000101;
    assign weights1[57][619] = 16'b1111111111110011;
    assign weights1[57][620] = 16'b1111111111111110;
    assign weights1[57][621] = 16'b1111111111110110;
    assign weights1[57][622] = 16'b1111111111111010;
    assign weights1[57][623] = 16'b0000000000000111;
    assign weights1[57][624] = 16'b1111111111101010;
    assign weights1[57][625] = 16'b1111111111110010;
    assign weights1[57][626] = 16'b0000000000000100;
    assign weights1[57][627] = 16'b1111111111100101;
    assign weights1[57][628] = 16'b1111111111111010;
    assign weights1[57][629] = 16'b0000000000001100;
    assign weights1[57][630] = 16'b0000000000001001;
    assign weights1[57][631] = 16'b0000000000000101;
    assign weights1[57][632] = 16'b0000000000000000;
    assign weights1[57][633] = 16'b1111111111111110;
    assign weights1[57][634] = 16'b1111111111111011;
    assign weights1[57][635] = 16'b0000000000000011;
    assign weights1[57][636] = 16'b1111111111111100;
    assign weights1[57][637] = 16'b0000000000001110;
    assign weights1[57][638] = 16'b0000000000000000;
    assign weights1[57][639] = 16'b0000000000000011;
    assign weights1[57][640] = 16'b0000000000000111;
    assign weights1[57][641] = 16'b1111111111111011;
    assign weights1[57][642] = 16'b1111111111110101;
    assign weights1[57][643] = 16'b1111111111110110;
    assign weights1[57][644] = 16'b1111111111111010;
    assign weights1[57][645] = 16'b1111111111111011;
    assign weights1[57][646] = 16'b1111111111110011;
    assign weights1[57][647] = 16'b0000000000000010;
    assign weights1[57][648] = 16'b1111111111111010;
    assign weights1[57][649] = 16'b0000000000010001;
    assign weights1[57][650] = 16'b1111111111110101;
    assign weights1[57][651] = 16'b1111111111111101;
    assign weights1[57][652] = 16'b1111111111101100;
    assign weights1[57][653] = 16'b0000000000000001;
    assign weights1[57][654] = 16'b1111111111111001;
    assign weights1[57][655] = 16'b0000000000000010;
    assign weights1[57][656] = 16'b1111111111110011;
    assign weights1[57][657] = 16'b1111111111111001;
    assign weights1[57][658] = 16'b0000000000001111;
    assign weights1[57][659] = 16'b1111111111111100;
    assign weights1[57][660] = 16'b0000000000001001;
    assign weights1[57][661] = 16'b0000000000001001;
    assign weights1[57][662] = 16'b0000000000001101;
    assign weights1[57][663] = 16'b0000000000001100;
    assign weights1[57][664] = 16'b0000000000000011;
    assign weights1[57][665] = 16'b1111111111111001;
    assign weights1[57][666] = 16'b1111111111111110;
    assign weights1[57][667] = 16'b1111111111110110;
    assign weights1[57][668] = 16'b1111111111111011;
    assign weights1[57][669] = 16'b1111111111110101;
    assign weights1[57][670] = 16'b1111111111111010;
    assign weights1[57][671] = 16'b1111111111110000;
    assign weights1[57][672] = 16'b0000000000000000;
    assign weights1[57][673] = 16'b0000000000000011;
    assign weights1[57][674] = 16'b0000000000000101;
    assign weights1[57][675] = 16'b1111111111110101;
    assign weights1[57][676] = 16'b0000000000000100;
    assign weights1[57][677] = 16'b1111111111111011;
    assign weights1[57][678] = 16'b0000000000000001;
    assign weights1[57][679] = 16'b0000000000000100;
    assign weights1[57][680] = 16'b0000000000000011;
    assign weights1[57][681] = 16'b1111111111111010;
    assign weights1[57][682] = 16'b0000000000001101;
    assign weights1[57][683] = 16'b0000000000000010;
    assign weights1[57][684] = 16'b0000000000001000;
    assign weights1[57][685] = 16'b1111111111011110;
    assign weights1[57][686] = 16'b1111111111110000;
    assign weights1[57][687] = 16'b0000000000000110;
    assign weights1[57][688] = 16'b1111111111110000;
    assign weights1[57][689] = 16'b1111111111111111;
    assign weights1[57][690] = 16'b0000000000001000;
    assign weights1[57][691] = 16'b1111111111110010;
    assign weights1[57][692] = 16'b0000000000000000;
    assign weights1[57][693] = 16'b0000000000010101;
    assign weights1[57][694] = 16'b1111111111101111;
    assign weights1[57][695] = 16'b1111111111110011;
    assign weights1[57][696] = 16'b1111111111101011;
    assign weights1[57][697] = 16'b1111111111110001;
    assign weights1[57][698] = 16'b1111111111111000;
    assign weights1[57][699] = 16'b1111111111101011;
    assign weights1[57][700] = 16'b0000000000000000;
    assign weights1[57][701] = 16'b0000000000000000;
    assign weights1[57][702] = 16'b0000000000001000;
    assign weights1[57][703] = 16'b0000000000000010;
    assign weights1[57][704] = 16'b0000000000000000;
    assign weights1[57][705] = 16'b1111111111110000;
    assign weights1[57][706] = 16'b1111111111111111;
    assign weights1[57][707] = 16'b0000000000001101;
    assign weights1[57][708] = 16'b1111111111110010;
    assign weights1[57][709] = 16'b0000000000001010;
    assign weights1[57][710] = 16'b1111111111110000;
    assign weights1[57][711] = 16'b1111111111101111;
    assign weights1[57][712] = 16'b0000000000000110;
    assign weights1[57][713] = 16'b1111111111111011;
    assign weights1[57][714] = 16'b0000000000001010;
    assign weights1[57][715] = 16'b1111111111110100;
    assign weights1[57][716] = 16'b1111111111110100;
    assign weights1[57][717] = 16'b0000000000000001;
    assign weights1[57][718] = 16'b1111111111111100;
    assign weights1[57][719] = 16'b1111111111011010;
    assign weights1[57][720] = 16'b1111111111100110;
    assign weights1[57][721] = 16'b1111111111100010;
    assign weights1[57][722] = 16'b1111111111101001;
    assign weights1[57][723] = 16'b1111111111100100;
    assign weights1[57][724] = 16'b1111111111101100;
    assign weights1[57][725] = 16'b1111111111101100;
    assign weights1[57][726] = 16'b1111111111110111;
    assign weights1[57][727] = 16'b1111111111110101;
    assign weights1[57][728] = 16'b0000000000000010;
    assign weights1[57][729] = 16'b1111111111111010;
    assign weights1[57][730] = 16'b1111111111111101;
    assign weights1[57][731] = 16'b1111111111111110;
    assign weights1[57][732] = 16'b0000000000001100;
    assign weights1[57][733] = 16'b0000000000000000;
    assign weights1[57][734] = 16'b1111111111111100;
    assign weights1[57][735] = 16'b1111111111111111;
    assign weights1[57][736] = 16'b1111111111111010;
    assign weights1[57][737] = 16'b1111111111111001;
    assign weights1[57][738] = 16'b1111111111110110;
    assign weights1[57][739] = 16'b0000000000000100;
    assign weights1[57][740] = 16'b1111111111110100;
    assign weights1[57][741] = 16'b1111111111111011;
    assign weights1[57][742] = 16'b1111111111101101;
    assign weights1[57][743] = 16'b0000000000001000;
    assign weights1[57][744] = 16'b1111111111111001;
    assign weights1[57][745] = 16'b1111111111101010;
    assign weights1[57][746] = 16'b1111111111110100;
    assign weights1[57][747] = 16'b1111111111110001;
    assign weights1[57][748] = 16'b1111111111110010;
    assign weights1[57][749] = 16'b1111111111110000;
    assign weights1[57][750] = 16'b1111111111101011;
    assign weights1[57][751] = 16'b1111111111101110;
    assign weights1[57][752] = 16'b1111111111101001;
    assign weights1[57][753] = 16'b1111111111101000;
    assign weights1[57][754] = 16'b1111111111110010;
    assign weights1[57][755] = 16'b1111111111111001;
    assign weights1[57][756] = 16'b1111111111111110;
    assign weights1[57][757] = 16'b1111111111111110;
    assign weights1[57][758] = 16'b1111111111111001;
    assign weights1[57][759] = 16'b1111111111111110;
    assign weights1[57][760] = 16'b1111111111110100;
    assign weights1[57][761] = 16'b0000000000000011;
    assign weights1[57][762] = 16'b0000000000000000;
    assign weights1[57][763] = 16'b1111111111101010;
    assign weights1[57][764] = 16'b1111111111101111;
    assign weights1[57][765] = 16'b1111111111100000;
    assign weights1[57][766] = 16'b1111111111111011;
    assign weights1[57][767] = 16'b1111111111110100;
    assign weights1[57][768] = 16'b1111111111111001;
    assign weights1[57][769] = 16'b1111111111111011;
    assign weights1[57][770] = 16'b1111111111110001;
    assign weights1[57][771] = 16'b1111111111101001;
    assign weights1[57][772] = 16'b1111111111111010;
    assign weights1[57][773] = 16'b1111111111101101;
    assign weights1[57][774] = 16'b1111111111101101;
    assign weights1[57][775] = 16'b1111111111101101;
    assign weights1[57][776] = 16'b1111111111100011;
    assign weights1[57][777] = 16'b1111111111101010;
    assign weights1[57][778] = 16'b1111111111011101;
    assign weights1[57][779] = 16'b1111111111110000;
    assign weights1[57][780] = 16'b1111111111101101;
    assign weights1[57][781] = 16'b1111111111110010;
    assign weights1[57][782] = 16'b1111111111110111;
    assign weights1[57][783] = 16'b1111111111111110;
    assign weights1[58][0] = 16'b0000000000000000;
    assign weights1[58][1] = 16'b0000000000000000;
    assign weights1[58][2] = 16'b0000000000000011;
    assign weights1[58][3] = 16'b0000000000000011;
    assign weights1[58][4] = 16'b1111111111111101;
    assign weights1[58][5] = 16'b0000000000000000;
    assign weights1[58][6] = 16'b0000000000000000;
    assign weights1[58][7] = 16'b0000000000010100;
    assign weights1[58][8] = 16'b0000000000011111;
    assign weights1[58][9] = 16'b0000000000011100;
    assign weights1[58][10] = 16'b0000000000011111;
    assign weights1[58][11] = 16'b0000000000010110;
    assign weights1[58][12] = 16'b1111111111111101;
    assign weights1[58][13] = 16'b1111111111111001;
    assign weights1[58][14] = 16'b0000000000010110;
    assign weights1[58][15] = 16'b0000000000001111;
    assign weights1[58][16] = 16'b1111111111111111;
    assign weights1[58][17] = 16'b1111111111101001;
    assign weights1[58][18] = 16'b0000000000001010;
    assign weights1[58][19] = 16'b1111111111111110;
    assign weights1[58][20] = 16'b0000000000000101;
    assign weights1[58][21] = 16'b1111111111111110;
    assign weights1[58][22] = 16'b1111111111111001;
    assign weights1[58][23] = 16'b1111111111111100;
    assign weights1[58][24] = 16'b0000000000000001;
    assign weights1[58][25] = 16'b0000000000000010;
    assign weights1[58][26] = 16'b0000000000000000;
    assign weights1[58][27] = 16'b0000000000000000;
    assign weights1[58][28] = 16'b0000000000000001;
    assign weights1[58][29] = 16'b0000000000000001;
    assign weights1[58][30] = 16'b0000000000000000;
    assign weights1[58][31] = 16'b0000000000000101;
    assign weights1[58][32] = 16'b0000000000000011;
    assign weights1[58][33] = 16'b1111111111111010;
    assign weights1[58][34] = 16'b0000000000010000;
    assign weights1[58][35] = 16'b0000000000001110;
    assign weights1[58][36] = 16'b0000000000011110;
    assign weights1[58][37] = 16'b0000000000100000;
    assign weights1[58][38] = 16'b0000000000010111;
    assign weights1[58][39] = 16'b0000000000100111;
    assign weights1[58][40] = 16'b0000000000010001;
    assign weights1[58][41] = 16'b0000000000000100;
    assign weights1[58][42] = 16'b0000000000010000;
    assign weights1[58][43] = 16'b0000000000000011;
    assign weights1[58][44] = 16'b1111111111110100;
    assign weights1[58][45] = 16'b1111111111111111;
    assign weights1[58][46] = 16'b0000000000001011;
    assign weights1[58][47] = 16'b1111111111111110;
    assign weights1[58][48] = 16'b0000000000001011;
    assign weights1[58][49] = 16'b0000000000000010;
    assign weights1[58][50] = 16'b0000000000000011;
    assign weights1[58][51] = 16'b0000000000000100;
    assign weights1[58][52] = 16'b0000000000000110;
    assign weights1[58][53] = 16'b0000000000000010;
    assign weights1[58][54] = 16'b0000000000000010;
    assign weights1[58][55] = 16'b0000000000000001;
    assign weights1[58][56] = 16'b0000000000000011;
    assign weights1[58][57] = 16'b0000000000000011;
    assign weights1[58][58] = 16'b0000000000000101;
    assign weights1[58][59] = 16'b0000000000000011;
    assign weights1[58][60] = 16'b1111111111111111;
    assign weights1[58][61] = 16'b0000000000000100;
    assign weights1[58][62] = 16'b0000000000001110;
    assign weights1[58][63] = 16'b0000000000010111;
    assign weights1[58][64] = 16'b0000000000010000;
    assign weights1[58][65] = 16'b0000000000001110;
    assign weights1[58][66] = 16'b0000000000011010;
    assign weights1[58][67] = 16'b0000000000001011;
    assign weights1[58][68] = 16'b0000000000001001;
    assign weights1[58][69] = 16'b0000000000001010;
    assign weights1[58][70] = 16'b0000000000000000;
    assign weights1[58][71] = 16'b0000000000001111;
    assign weights1[58][72] = 16'b0000000000001100;
    assign weights1[58][73] = 16'b1111111111111100;
    assign weights1[58][74] = 16'b1111111111101111;
    assign weights1[58][75] = 16'b0000000000001101;
    assign weights1[58][76] = 16'b0000000000010000;
    assign weights1[58][77] = 16'b0000000000000001;
    assign weights1[58][78] = 16'b0000000000001100;
    assign weights1[58][79] = 16'b1111111111111111;
    assign weights1[58][80] = 16'b0000000000010001;
    assign weights1[58][81] = 16'b0000000000000010;
    assign weights1[58][82] = 16'b0000000000000011;
    assign weights1[58][83] = 16'b0000000000000010;
    assign weights1[58][84] = 16'b0000000000000111;
    assign weights1[58][85] = 16'b0000000000000010;
    assign weights1[58][86] = 16'b0000000000001000;
    assign weights1[58][87] = 16'b0000000000001000;
    assign weights1[58][88] = 16'b1111111111111100;
    assign weights1[58][89] = 16'b0000000000000100;
    assign weights1[58][90] = 16'b0000000000010100;
    assign weights1[58][91] = 16'b0000000000010110;
    assign weights1[58][92] = 16'b0000000000011001;
    assign weights1[58][93] = 16'b0000000000010111;
    assign weights1[58][94] = 16'b0000000000011000;
    assign weights1[58][95] = 16'b0000000000010101;
    assign weights1[58][96] = 16'b0000000000011000;
    assign weights1[58][97] = 16'b0000000000000100;
    assign weights1[58][98] = 16'b0000000000001100;
    assign weights1[58][99] = 16'b0000000000010111;
    assign weights1[58][100] = 16'b0000000000001000;
    assign weights1[58][101] = 16'b0000000000011011;
    assign weights1[58][102] = 16'b0000000000010011;
    assign weights1[58][103] = 16'b0000000000010000;
    assign weights1[58][104] = 16'b0000000000010111;
    assign weights1[58][105] = 16'b0000000000001111;
    assign weights1[58][106] = 16'b0000000000011110;
    assign weights1[58][107] = 16'b0000000000011111;
    assign weights1[58][108] = 16'b0000000000100000;
    assign weights1[58][109] = 16'b0000000000010010;
    assign weights1[58][110] = 16'b0000000000010000;
    assign weights1[58][111] = 16'b1111111111111110;
    assign weights1[58][112] = 16'b0000000000001001;
    assign weights1[58][113] = 16'b0000000000000111;
    assign weights1[58][114] = 16'b0000000000001001;
    assign weights1[58][115] = 16'b0000000000000000;
    assign weights1[58][116] = 16'b0000000000010001;
    assign weights1[58][117] = 16'b0000000000000001;
    assign weights1[58][118] = 16'b0000000000001111;
    assign weights1[58][119] = 16'b0000000000100011;
    assign weights1[58][120] = 16'b0000000000100001;
    assign weights1[58][121] = 16'b1111111111111100;
    assign weights1[58][122] = 16'b0000000000010100;
    assign weights1[58][123] = 16'b0000000000010010;
    assign weights1[58][124] = 16'b0000000000001000;
    assign weights1[58][125] = 16'b0000000000011001;
    assign weights1[58][126] = 16'b0000000000010010;
    assign weights1[58][127] = 16'b0000000000000001;
    assign weights1[58][128] = 16'b0000000000010100;
    assign weights1[58][129] = 16'b0000000000011010;
    assign weights1[58][130] = 16'b0000000000010011;
    assign weights1[58][131] = 16'b0000000000001011;
    assign weights1[58][132] = 16'b0000000000000010;
    assign weights1[58][133] = 16'b1111111111111001;
    assign weights1[58][134] = 16'b0000000000000100;
    assign weights1[58][135] = 16'b0000000000000110;
    assign weights1[58][136] = 16'b0000000000011000;
    assign weights1[58][137] = 16'b0000000000010100;
    assign weights1[58][138] = 16'b0000000000010000;
    assign weights1[58][139] = 16'b0000000000001010;
    assign weights1[58][140] = 16'b0000000000000110;
    assign weights1[58][141] = 16'b0000000000001101;
    assign weights1[58][142] = 16'b0000000000001011;
    assign weights1[58][143] = 16'b0000000000000100;
    assign weights1[58][144] = 16'b0000000000000000;
    assign weights1[58][145] = 16'b0000000000001110;
    assign weights1[58][146] = 16'b0000000000011010;
    assign weights1[58][147] = 16'b0000000000011100;
    assign weights1[58][148] = 16'b1111111111111011;
    assign weights1[58][149] = 16'b0000000000100110;
    assign weights1[58][150] = 16'b0000000000000100;
    assign weights1[58][151] = 16'b0000000000000001;
    assign weights1[58][152] = 16'b0000000000001001;
    assign weights1[58][153] = 16'b0000000000001110;
    assign weights1[58][154] = 16'b0000000000001111;
    assign weights1[58][155] = 16'b0000000000000011;
    assign weights1[58][156] = 16'b0000000000101010;
    assign weights1[58][157] = 16'b0000000000010101;
    assign weights1[58][158] = 16'b0000000000001101;
    assign weights1[58][159] = 16'b0000000000000100;
    assign weights1[58][160] = 16'b0000000000100100;
    assign weights1[58][161] = 16'b0000000000010000;
    assign weights1[58][162] = 16'b0000000000011010;
    assign weights1[58][163] = 16'b0000000000011100;
    assign weights1[58][164] = 16'b0000000000101011;
    assign weights1[58][165] = 16'b0000000000100100;
    assign weights1[58][166] = 16'b0000000000001010;
    assign weights1[58][167] = 16'b0000000000001101;
    assign weights1[58][168] = 16'b0000000000000101;
    assign weights1[58][169] = 16'b1111111111111111;
    assign weights1[58][170] = 16'b0000000000000000;
    assign weights1[58][171] = 16'b1111111111111010;
    assign weights1[58][172] = 16'b1111111111101101;
    assign weights1[58][173] = 16'b0000000000010011;
    assign weights1[58][174] = 16'b0000000000010011;
    assign weights1[58][175] = 16'b0000000000001100;
    assign weights1[58][176] = 16'b0000000000010011;
    assign weights1[58][177] = 16'b1111111111111001;
    assign weights1[58][178] = 16'b0000000000001001;
    assign weights1[58][179] = 16'b0000000000011100;
    assign weights1[58][180] = 16'b0000000000100001;
    assign weights1[58][181] = 16'b0000000000000011;
    assign weights1[58][182] = 16'b0000000000000111;
    assign weights1[58][183] = 16'b0000000000011110;
    assign weights1[58][184] = 16'b0000000000010100;
    assign weights1[58][185] = 16'b0000000000001011;
    assign weights1[58][186] = 16'b0000000000101000;
    assign weights1[58][187] = 16'b0000000000011111;
    assign weights1[58][188] = 16'b0000000000100111;
    assign weights1[58][189] = 16'b0000000000011111;
    assign weights1[58][190] = 16'b0000000000101110;
    assign weights1[58][191] = 16'b0000000000011101;
    assign weights1[58][192] = 16'b0000000000101100;
    assign weights1[58][193] = 16'b0000000000011111;
    assign weights1[58][194] = 16'b0000000000001010;
    assign weights1[58][195] = 16'b0000000000000100;
    assign weights1[58][196] = 16'b1111111111111111;
    assign weights1[58][197] = 16'b1111111111110111;
    assign weights1[58][198] = 16'b1111111111101011;
    assign weights1[58][199] = 16'b1111111111101110;
    assign weights1[58][200] = 16'b1111111111110101;
    assign weights1[58][201] = 16'b0000000000000011;
    assign weights1[58][202] = 16'b0000000000011110;
    assign weights1[58][203] = 16'b0000000000011111;
    assign weights1[58][204] = 16'b0000000000011000;
    assign weights1[58][205] = 16'b0000000000010000;
    assign weights1[58][206] = 16'b0000000000100111;
    assign weights1[58][207] = 16'b0000000000001111;
    assign weights1[58][208] = 16'b0000000000100010;
    assign weights1[58][209] = 16'b1111111111110101;
    assign weights1[58][210] = 16'b0000000000011010;
    assign weights1[58][211] = 16'b0000000000000000;
    assign weights1[58][212] = 16'b0000000000000100;
    assign weights1[58][213] = 16'b0000000000010101;
    assign weights1[58][214] = 16'b0000000000011010;
    assign weights1[58][215] = 16'b0000000000001101;
    assign weights1[58][216] = 16'b0000000000011011;
    assign weights1[58][217] = 16'b0000000000000110;
    assign weights1[58][218] = 16'b0000000000000101;
    assign weights1[58][219] = 16'b0000000001000011;
    assign weights1[58][220] = 16'b0000000000011001;
    assign weights1[58][221] = 16'b0000000000100000;
    assign weights1[58][222] = 16'b0000000000000110;
    assign weights1[58][223] = 16'b0000000000000111;
    assign weights1[58][224] = 16'b1111111111111000;
    assign weights1[58][225] = 16'b1111111111101101;
    assign weights1[58][226] = 16'b1111111111100101;
    assign weights1[58][227] = 16'b1111111111011101;
    assign weights1[58][228] = 16'b1111111111010110;
    assign weights1[58][229] = 16'b1111111111111110;
    assign weights1[58][230] = 16'b0000000000101101;
    assign weights1[58][231] = 16'b0000000000100010;
    assign weights1[58][232] = 16'b0000000000100110;
    assign weights1[58][233] = 16'b0000000000010001;
    assign weights1[58][234] = 16'b0000000000011001;
    assign weights1[58][235] = 16'b0000000000011110;
    assign weights1[58][236] = 16'b0000000000001101;
    assign weights1[58][237] = 16'b0000000000001011;
    assign weights1[58][238] = 16'b0000000000011001;
    assign weights1[58][239] = 16'b0000000000010110;
    assign weights1[58][240] = 16'b0000000000010000;
    assign weights1[58][241] = 16'b0000000000000111;
    assign weights1[58][242] = 16'b0000000000001111;
    assign weights1[58][243] = 16'b0000000000011111;
    assign weights1[58][244] = 16'b0000000000011111;
    assign weights1[58][245] = 16'b0000000000011111;
    assign weights1[58][246] = 16'b0000000000100011;
    assign weights1[58][247] = 16'b0000000000101000;
    assign weights1[58][248] = 16'b0000000000100011;
    assign weights1[58][249] = 16'b0000000000000001;
    assign weights1[58][250] = 16'b1111111111111000;
    assign weights1[58][251] = 16'b1111111111111111;
    assign weights1[58][252] = 16'b1111111111110010;
    assign weights1[58][253] = 16'b1111111111100010;
    assign weights1[58][254] = 16'b1111111111011110;
    assign weights1[58][255] = 16'b1111111111000110;
    assign weights1[58][256] = 16'b1111111111000100;
    assign weights1[58][257] = 16'b1111111111011001;
    assign weights1[58][258] = 16'b0000000000001101;
    assign weights1[58][259] = 16'b0000000000011001;
    assign weights1[58][260] = 16'b0000000000010001;
    assign weights1[58][261] = 16'b0000000000110011;
    assign weights1[58][262] = 16'b0000000000101100;
    assign weights1[58][263] = 16'b0000000000111011;
    assign weights1[58][264] = 16'b0000000000010010;
    assign weights1[58][265] = 16'b0000000000111000;
    assign weights1[58][266] = 16'b0000000000101100;
    assign weights1[58][267] = 16'b0000000000001100;
    assign weights1[58][268] = 16'b0000000000001101;
    assign weights1[58][269] = 16'b0000000000001111;
    assign weights1[58][270] = 16'b0000000000000101;
    assign weights1[58][271] = 16'b0000000000000110;
    assign weights1[58][272] = 16'b0000000000000101;
    assign weights1[58][273] = 16'b0000000000101011;
    assign weights1[58][274] = 16'b0000000000100001;
    assign weights1[58][275] = 16'b0000000000001001;
    assign weights1[58][276] = 16'b1111111111110011;
    assign weights1[58][277] = 16'b1111111111101100;
    assign weights1[58][278] = 16'b1111111111110001;
    assign weights1[58][279] = 16'b1111111111110011;
    assign weights1[58][280] = 16'b1111111111101010;
    assign weights1[58][281] = 16'b1111111111011101;
    assign weights1[58][282] = 16'b1111111111010100;
    assign weights1[58][283] = 16'b1111111111000010;
    assign weights1[58][284] = 16'b1111111110111010;
    assign weights1[58][285] = 16'b1111111110100010;
    assign weights1[58][286] = 16'b1111111111001111;
    assign weights1[58][287] = 16'b1111111111111111;
    assign weights1[58][288] = 16'b0000000000011000;
    assign weights1[58][289] = 16'b0000000000010100;
    assign weights1[58][290] = 16'b0000000000011011;
    assign weights1[58][291] = 16'b0000000000110001;
    assign weights1[58][292] = 16'b0000000000110000;
    assign weights1[58][293] = 16'b0000000000010010;
    assign weights1[58][294] = 16'b0000000000011100;
    assign weights1[58][295] = 16'b0000000000100010;
    assign weights1[58][296] = 16'b0000000000101001;
    assign weights1[58][297] = 16'b1111111111111101;
    assign weights1[58][298] = 16'b0000000000001110;
    assign weights1[58][299] = 16'b0000000000001001;
    assign weights1[58][300] = 16'b0000000000111011;
    assign weights1[58][301] = 16'b0000000001000000;
    assign weights1[58][302] = 16'b0000000000110010;
    assign weights1[58][303] = 16'b1111111111110010;
    assign weights1[58][304] = 16'b1111111111011000;
    assign weights1[58][305] = 16'b1111111111100110;
    assign weights1[58][306] = 16'b1111111111100000;
    assign weights1[58][307] = 16'b1111111111100101;
    assign weights1[58][308] = 16'b1111111111100111;
    assign weights1[58][309] = 16'b1111111111011100;
    assign weights1[58][310] = 16'b1111111111001111;
    assign weights1[58][311] = 16'b1111111111001110;
    assign weights1[58][312] = 16'b1111111110111001;
    assign weights1[58][313] = 16'b1111111110001010;
    assign weights1[58][314] = 16'b1111111110010001;
    assign weights1[58][315] = 16'b1111111111011000;
    assign weights1[58][316] = 16'b1111111111101010;
    assign weights1[58][317] = 16'b0000000000000110;
    assign weights1[58][318] = 16'b0000000000011111;
    assign weights1[58][319] = 16'b0000000000101110;
    assign weights1[58][320] = 16'b0000000000111101;
    assign weights1[58][321] = 16'b0000000000011100;
    assign weights1[58][322] = 16'b0000000000110000;
    assign weights1[58][323] = 16'b0000000000100101;
    assign weights1[58][324] = 16'b0000000000100101;
    assign weights1[58][325] = 16'b0000000000100001;
    assign weights1[58][326] = 16'b0000000000101000;
    assign weights1[58][327] = 16'b0000000000010000;
    assign weights1[58][328] = 16'b0000000000000010;
    assign weights1[58][329] = 16'b0000000000000001;
    assign weights1[58][330] = 16'b1111111111011100;
    assign weights1[58][331] = 16'b1111111111010000;
    assign weights1[58][332] = 16'b1111111111001000;
    assign weights1[58][333] = 16'b1111111111011110;
    assign weights1[58][334] = 16'b1111111111100111;
    assign weights1[58][335] = 16'b1111111111100011;
    assign weights1[58][336] = 16'b1111111111100111;
    assign weights1[58][337] = 16'b1111111111100100;
    assign weights1[58][338] = 16'b1111111111100001;
    assign weights1[58][339] = 16'b1111111111011010;
    assign weights1[58][340] = 16'b1111111111010100;
    assign weights1[58][341] = 16'b1111111110110011;
    assign weights1[58][342] = 16'b1111111110010100;
    assign weights1[58][343] = 16'b1111111110010110;
    assign weights1[58][344] = 16'b1111111110110001;
    assign weights1[58][345] = 16'b1111111111111100;
    assign weights1[58][346] = 16'b1111111111111111;
    assign weights1[58][347] = 16'b0000000000101010;
    assign weights1[58][348] = 16'b0000000000111000;
    assign weights1[58][349] = 16'b0000000000101111;
    assign weights1[58][350] = 16'b0000000000011111;
    assign weights1[58][351] = 16'b0000000000011001;
    assign weights1[58][352] = 16'b0000000000011001;
    assign weights1[58][353] = 16'b0000000000011010;
    assign weights1[58][354] = 16'b0000000000000111;
    assign weights1[58][355] = 16'b1111111111110010;
    assign weights1[58][356] = 16'b1111111111100000;
    assign weights1[58][357] = 16'b1111111111000010;
    assign weights1[58][358] = 16'b1111111110010111;
    assign weights1[58][359] = 16'b1111111110100011;
    assign weights1[58][360] = 16'b1111111110111001;
    assign weights1[58][361] = 16'b1111111111010110;
    assign weights1[58][362] = 16'b1111111111010111;
    assign weights1[58][363] = 16'b1111111111100000;
    assign weights1[58][364] = 16'b1111111111110011;
    assign weights1[58][365] = 16'b1111111111101111;
    assign weights1[58][366] = 16'b1111111111110110;
    assign weights1[58][367] = 16'b1111111111111001;
    assign weights1[58][368] = 16'b1111111111100001;
    assign weights1[58][369] = 16'b1111111111011110;
    assign weights1[58][370] = 16'b1111111110111110;
    assign weights1[58][371] = 16'b1111111110101110;
    assign weights1[58][372] = 16'b1111111110100001;
    assign weights1[58][373] = 16'b1111111110101111;
    assign weights1[58][374] = 16'b1111111111001010;
    assign weights1[58][375] = 16'b1111111111100100;
    assign weights1[58][376] = 16'b0000000000110001;
    assign weights1[58][377] = 16'b0000000000110101;
    assign weights1[58][378] = 16'b0000000000100111;
    assign weights1[58][379] = 16'b0000000000101010;
    assign weights1[58][380] = 16'b0000000000001000;
    assign weights1[58][381] = 16'b1111111111110110;
    assign weights1[58][382] = 16'b1111111111101110;
    assign weights1[58][383] = 16'b1111111111100100;
    assign weights1[58][384] = 16'b1111111110010110;
    assign weights1[58][385] = 16'b1111111101111011;
    assign weights1[58][386] = 16'b1111111110010101;
    assign weights1[58][387] = 16'b1111111110110100;
    assign weights1[58][388] = 16'b1111111111001100;
    assign weights1[58][389] = 16'b1111111111011100;
    assign weights1[58][390] = 16'b1111111111101000;
    assign weights1[58][391] = 16'b1111111111101100;
    assign weights1[58][392] = 16'b0000000000000011;
    assign weights1[58][393] = 16'b0000000000000000;
    assign weights1[58][394] = 16'b1111111111111110;
    assign weights1[58][395] = 16'b1111111111111000;
    assign weights1[58][396] = 16'b0000000000001001;
    assign weights1[58][397] = 16'b1111111111110001;
    assign weights1[58][398] = 16'b1111111111111001;
    assign weights1[58][399] = 16'b1111111111000010;
    assign weights1[58][400] = 16'b1111111110111110;
    assign weights1[58][401] = 16'b1111111110110101;
    assign weights1[58][402] = 16'b1111111111000001;
    assign weights1[58][403] = 16'b1111111110111111;
    assign weights1[58][404] = 16'b1111111111011100;
    assign weights1[58][405] = 16'b0000000000001011;
    assign weights1[58][406] = 16'b0000000000000000;
    assign weights1[58][407] = 16'b0000000000000000;
    assign weights1[58][408] = 16'b1111111111111101;
    assign weights1[58][409] = 16'b1111111111101110;
    assign weights1[58][410] = 16'b1111111111010011;
    assign weights1[58][411] = 16'b1111111111010011;
    assign weights1[58][412] = 16'b1111111110111010;
    assign weights1[58][413] = 16'b1111111110101001;
    assign weights1[58][414] = 16'b1111111111000001;
    assign weights1[58][415] = 16'b1111111110111101;
    assign weights1[58][416] = 16'b1111111111001100;
    assign weights1[58][417] = 16'b1111111111100111;
    assign weights1[58][418] = 16'b1111111111110010;
    assign weights1[58][419] = 16'b1111111111110001;
    assign weights1[58][420] = 16'b0000000000000000;
    assign weights1[58][421] = 16'b1111111111111000;
    assign weights1[58][422] = 16'b1111111111110011;
    assign weights1[58][423] = 16'b1111111111111010;
    assign weights1[58][424] = 16'b0000000000001110;
    assign weights1[58][425] = 16'b0000000000001110;
    assign weights1[58][426] = 16'b1111111111110101;
    assign weights1[58][427] = 16'b1111111111111110;
    assign weights1[58][428] = 16'b1111111111011111;
    assign weights1[58][429] = 16'b1111111111001010;
    assign weights1[58][430] = 16'b1111111110110110;
    assign weights1[58][431] = 16'b1111111110101110;
    assign weights1[58][432] = 16'b1111111111000111;
    assign weights1[58][433] = 16'b1111111111110101;
    assign weights1[58][434] = 16'b1111111111101001;
    assign weights1[58][435] = 16'b1111111111011111;
    assign weights1[58][436] = 16'b1111111111101000;
    assign weights1[58][437] = 16'b1111111111010100;
    assign weights1[58][438] = 16'b1111111111101100;
    assign weights1[58][439] = 16'b1111111111011110;
    assign weights1[58][440] = 16'b1111111111110101;
    assign weights1[58][441] = 16'b0000000000000010;
    assign weights1[58][442] = 16'b1111111111010010;
    assign weights1[58][443] = 16'b1111111111000111;
    assign weights1[58][444] = 16'b1111111111001110;
    assign weights1[58][445] = 16'b1111111111101100;
    assign weights1[58][446] = 16'b1111111111101111;
    assign weights1[58][447] = 16'b1111111111101111;
    assign weights1[58][448] = 16'b0000000000000101;
    assign weights1[58][449] = 16'b1111111111110101;
    assign weights1[58][450] = 16'b0000000000000010;
    assign weights1[58][451] = 16'b1111111111111001;
    assign weights1[58][452] = 16'b0000000000000100;
    assign weights1[58][453] = 16'b0000000000010011;
    assign weights1[58][454] = 16'b0000000000000111;
    assign weights1[58][455] = 16'b0000000000010001;
    assign weights1[58][456] = 16'b1111111111110110;
    assign weights1[58][457] = 16'b1111111111110010;
    assign weights1[58][458] = 16'b1111111111011110;
    assign weights1[58][459] = 16'b1111111111100011;
    assign weights1[58][460] = 16'b1111111110111100;
    assign weights1[58][461] = 16'b1111111110111101;
    assign weights1[58][462] = 16'b1111111111101000;
    assign weights1[58][463] = 16'b1111111111101110;
    assign weights1[58][464] = 16'b1111111111011100;
    assign weights1[58][465] = 16'b1111111111100110;
    assign weights1[58][466] = 16'b1111111111011100;
    assign weights1[58][467] = 16'b1111111111111100;
    assign weights1[58][468] = 16'b0000000000011000;
    assign weights1[58][469] = 16'b1111111111111000;
    assign weights1[58][470] = 16'b1111111110111101;
    assign weights1[58][471] = 16'b1111111110111010;
    assign weights1[58][472] = 16'b1111111111010100;
    assign weights1[58][473] = 16'b1111111111100111;
    assign weights1[58][474] = 16'b1111111111110010;
    assign weights1[58][475] = 16'b1111111111110110;
    assign weights1[58][476] = 16'b0000000000000000;
    assign weights1[58][477] = 16'b0000000000000011;
    assign weights1[58][478] = 16'b0000000000001101;
    assign weights1[58][479] = 16'b0000000000001100;
    assign weights1[58][480] = 16'b0000000000000000;
    assign weights1[58][481] = 16'b1111111111110111;
    assign weights1[58][482] = 16'b0000000000001101;
    assign weights1[58][483] = 16'b0000000000000010;
    assign weights1[58][484] = 16'b0000000000000011;
    assign weights1[58][485] = 16'b0000000000001010;
    assign weights1[58][486] = 16'b1111111111100101;
    assign weights1[58][487] = 16'b1111111111111001;
    assign weights1[58][488] = 16'b1111111111011101;
    assign weights1[58][489] = 16'b1111111111010000;
    assign weights1[58][490] = 16'b1111111111101100;
    assign weights1[58][491] = 16'b1111111111101000;
    assign weights1[58][492] = 16'b0000000000000110;
    assign weights1[58][493] = 16'b0000000000000101;
    assign weights1[58][494] = 16'b1111111111111100;
    assign weights1[58][495] = 16'b1111111111111010;
    assign weights1[58][496] = 16'b0000000000000001;
    assign weights1[58][497] = 16'b0000000000000111;
    assign weights1[58][498] = 16'b1111111111001110;
    assign weights1[58][499] = 16'b1111111111001001;
    assign weights1[58][500] = 16'b1111111111011011;
    assign weights1[58][501] = 16'b1111111111100010;
    assign weights1[58][502] = 16'b1111111111111000;
    assign weights1[58][503] = 16'b1111111111110101;
    assign weights1[58][504] = 16'b1111111111111110;
    assign weights1[58][505] = 16'b1111111111111011;
    assign weights1[58][506] = 16'b1111111111111101;
    assign weights1[58][507] = 16'b1111111111111010;
    assign weights1[58][508] = 16'b1111111111110111;
    assign weights1[58][509] = 16'b1111111111111000;
    assign weights1[58][510] = 16'b1111111111110111;
    assign weights1[58][511] = 16'b0000000000010000;
    assign weights1[58][512] = 16'b0000000000000101;
    assign weights1[58][513] = 16'b1111111111101101;
    assign weights1[58][514] = 16'b1111111111111101;
    assign weights1[58][515] = 16'b1111111111111011;
    assign weights1[58][516] = 16'b1111111111010001;
    assign weights1[58][517] = 16'b1111111111110000;
    assign weights1[58][518] = 16'b1111111111100111;
    assign weights1[58][519] = 16'b1111111111101011;
    assign weights1[58][520] = 16'b1111111111111001;
    assign weights1[58][521] = 16'b1111111111110111;
    assign weights1[58][522] = 16'b0000000000001000;
    assign weights1[58][523] = 16'b0000000000010111;
    assign weights1[58][524] = 16'b0000000000010110;
    assign weights1[58][525] = 16'b0000000000001111;
    assign weights1[58][526] = 16'b1111111111000110;
    assign weights1[58][527] = 16'b1111111111001111;
    assign weights1[58][528] = 16'b1111111111010100;
    assign weights1[58][529] = 16'b1111111111100010;
    assign weights1[58][530] = 16'b1111111111111001;
    assign weights1[58][531] = 16'b1111111111110111;
    assign weights1[58][532] = 16'b1111111111110111;
    assign weights1[58][533] = 16'b1111111111110001;
    assign weights1[58][534] = 16'b1111111111101101;
    assign weights1[58][535] = 16'b1111111111100101;
    assign weights1[58][536] = 16'b0000000000001101;
    assign weights1[58][537] = 16'b1111111111110110;
    assign weights1[58][538] = 16'b0000000000010101;
    assign weights1[58][539] = 16'b0000000000000011;
    assign weights1[58][540] = 16'b0000000000010001;
    assign weights1[58][541] = 16'b1111111111101100;
    assign weights1[58][542] = 16'b1111111111101000;
    assign weights1[58][543] = 16'b1111111111111000;
    assign weights1[58][544] = 16'b0000000000000011;
    assign weights1[58][545] = 16'b0000000000000100;
    assign weights1[58][546] = 16'b1111111111111111;
    assign weights1[58][547] = 16'b1111111111101000;
    assign weights1[58][548] = 16'b1111111111110100;
    assign weights1[58][549] = 16'b1111111111111011;
    assign weights1[58][550] = 16'b1111111111111001;
    assign weights1[58][551] = 16'b0000000000001010;
    assign weights1[58][552] = 16'b0000000000011100;
    assign weights1[58][553] = 16'b1111111111101000;
    assign weights1[58][554] = 16'b1111111111001101;
    assign weights1[58][555] = 16'b1111111111000111;
    assign weights1[58][556] = 16'b1111111111101000;
    assign weights1[58][557] = 16'b1111111111101011;
    assign weights1[58][558] = 16'b1111111111110100;
    assign weights1[58][559] = 16'b1111111111111000;
    assign weights1[58][560] = 16'b1111111111111011;
    assign weights1[58][561] = 16'b1111111111110101;
    assign weights1[58][562] = 16'b1111111111110110;
    assign weights1[58][563] = 16'b1111111111100000;
    assign weights1[58][564] = 16'b1111111111110101;
    assign weights1[58][565] = 16'b1111111111101101;
    assign weights1[58][566] = 16'b0000000000000010;
    assign weights1[58][567] = 16'b1111111111110100;
    assign weights1[58][568] = 16'b1111111111111110;
    assign weights1[58][569] = 16'b1111111111111001;
    assign weights1[58][570] = 16'b0000000000000101;
    assign weights1[58][571] = 16'b1111111111111111;
    assign weights1[58][572] = 16'b1111111111011000;
    assign weights1[58][573] = 16'b1111111111110110;
    assign weights1[58][574] = 16'b1111111111111001;
    assign weights1[58][575] = 16'b1111111111101101;
    assign weights1[58][576] = 16'b1111111111101010;
    assign weights1[58][577] = 16'b0000000000001000;
    assign weights1[58][578] = 16'b1111111111110100;
    assign weights1[58][579] = 16'b1111111111111001;
    assign weights1[58][580] = 16'b0000000000000101;
    assign weights1[58][581] = 16'b1111111111110000;
    assign weights1[58][582] = 16'b1111111110111110;
    assign weights1[58][583] = 16'b1111111111011010;
    assign weights1[58][584] = 16'b1111111111101111;
    assign weights1[58][585] = 16'b1111111111110110;
    assign weights1[58][586] = 16'b1111111111111000;
    assign weights1[58][587] = 16'b1111111111110110;
    assign weights1[58][588] = 16'b0000000000000010;
    assign weights1[58][589] = 16'b1111111111111100;
    assign weights1[58][590] = 16'b1111111111111010;
    assign weights1[58][591] = 16'b1111111111100001;
    assign weights1[58][592] = 16'b1111111111111010;
    assign weights1[58][593] = 16'b1111111111100110;
    assign weights1[58][594] = 16'b1111111111111000;
    assign weights1[58][595] = 16'b1111111111101010;
    assign weights1[58][596] = 16'b0000000000000111;
    assign weights1[58][597] = 16'b1111111111110110;
    assign weights1[58][598] = 16'b1111111111111101;
    assign weights1[58][599] = 16'b0000000000000000;
    assign weights1[58][600] = 16'b1111111111111000;
    assign weights1[58][601] = 16'b1111111111110111;
    assign weights1[58][602] = 16'b1111111111110100;
    assign weights1[58][603] = 16'b0000000000000001;
    assign weights1[58][604] = 16'b1111111111101001;
    assign weights1[58][605] = 16'b1111111111111001;
    assign weights1[58][606] = 16'b0000000000000001;
    assign weights1[58][607] = 16'b1111111111100011;
    assign weights1[58][608] = 16'b0000000000000100;
    assign weights1[58][609] = 16'b1111111111000111;
    assign weights1[58][610] = 16'b1111111110111110;
    assign weights1[58][611] = 16'b1111111111010110;
    assign weights1[58][612] = 16'b1111111111110011;
    assign weights1[58][613] = 16'b1111111111110100;
    assign weights1[58][614] = 16'b1111111111111101;
    assign weights1[58][615] = 16'b1111111111111011;
    assign weights1[58][616] = 16'b1111111111111100;
    assign weights1[58][617] = 16'b1111111111111100;
    assign weights1[58][618] = 16'b1111111111110010;
    assign weights1[58][619] = 16'b1111111111101111;
    assign weights1[58][620] = 16'b1111111111100011;
    assign weights1[58][621] = 16'b1111111111111010;
    assign weights1[58][622] = 16'b1111111111101000;
    assign weights1[58][623] = 16'b1111111111110111;
    assign weights1[58][624] = 16'b1111111111101111;
    assign weights1[58][625] = 16'b1111111111100110;
    assign weights1[58][626] = 16'b1111111111111011;
    assign weights1[58][627] = 16'b1111111111111111;
    assign weights1[58][628] = 16'b1111111111101011;
    assign weights1[58][629] = 16'b0000000000000000;
    assign weights1[58][630] = 16'b1111111111101110;
    assign weights1[58][631] = 16'b0000000000000001;
    assign weights1[58][632] = 16'b1111111111110000;
    assign weights1[58][633] = 16'b0000000000010101;
    assign weights1[58][634] = 16'b1111111111101010;
    assign weights1[58][635] = 16'b1111111111010111;
    assign weights1[58][636] = 16'b1111111111000111;
    assign weights1[58][637] = 16'b1111111111001100;
    assign weights1[58][638] = 16'b1111111111100001;
    assign weights1[58][639] = 16'b1111111111101111;
    assign weights1[58][640] = 16'b1111111111110101;
    assign weights1[58][641] = 16'b1111111111111011;
    assign weights1[58][642] = 16'b1111111111111111;
    assign weights1[58][643] = 16'b1111111111111111;
    assign weights1[58][644] = 16'b1111111111111100;
    assign weights1[58][645] = 16'b1111111111111110;
    assign weights1[58][646] = 16'b1111111111110011;
    assign weights1[58][647] = 16'b1111111111111101;
    assign weights1[58][648] = 16'b1111111111100010;
    assign weights1[58][649] = 16'b1111111111100111;
    assign weights1[58][650] = 16'b1111111111100010;
    assign weights1[58][651] = 16'b1111111111101111;
    assign weights1[58][652] = 16'b0000000000000010;
    assign weights1[58][653] = 16'b1111111111110011;
    assign weights1[58][654] = 16'b1111111111111000;
    assign weights1[58][655] = 16'b1111111111111110;
    assign weights1[58][656] = 16'b0000000000001001;
    assign weights1[58][657] = 16'b0000000000000111;
    assign weights1[58][658] = 16'b1111111111110000;
    assign weights1[58][659] = 16'b1111111111111000;
    assign weights1[58][660] = 16'b1111111111110011;
    assign weights1[58][661] = 16'b0000000000000110;
    assign weights1[58][662] = 16'b1111111111101010;
    assign weights1[58][663] = 16'b1111111111100101;
    assign weights1[58][664] = 16'b1111111111011110;
    assign weights1[58][665] = 16'b1111111111010010;
    assign weights1[58][666] = 16'b1111111111100111;
    assign weights1[58][667] = 16'b1111111111111011;
    assign weights1[58][668] = 16'b1111111111110110;
    assign weights1[58][669] = 16'b1111111111111100;
    assign weights1[58][670] = 16'b1111111111111101;
    assign weights1[58][671] = 16'b0000000000000000;
    assign weights1[58][672] = 16'b0000000000000000;
    assign weights1[58][673] = 16'b1111111111111111;
    assign weights1[58][674] = 16'b1111111111111101;
    assign weights1[58][675] = 16'b1111111111111110;
    assign weights1[58][676] = 16'b0000000000000011;
    assign weights1[58][677] = 16'b1111111111110000;
    assign weights1[58][678] = 16'b1111111111010111;
    assign weights1[58][679] = 16'b0000000000010101;
    assign weights1[58][680] = 16'b1111111111111010;
    assign weights1[58][681] = 16'b1111111111111001;
    assign weights1[58][682] = 16'b1111111111111101;
    assign weights1[58][683] = 16'b1111111111100111;
    assign weights1[58][684] = 16'b1111111111111110;
    assign weights1[58][685] = 16'b0000000000010001;
    assign weights1[58][686] = 16'b1111111111010010;
    assign weights1[58][687] = 16'b0000000000010100;
    assign weights1[58][688] = 16'b0000000000001001;
    assign weights1[58][689] = 16'b1111111111101000;
    assign weights1[58][690] = 16'b1111111111010101;
    assign weights1[58][691] = 16'b1111111111100000;
    assign weights1[58][692] = 16'b1111111111011001;
    assign weights1[58][693] = 16'b1111111111100001;
    assign weights1[58][694] = 16'b1111111111101101;
    assign weights1[58][695] = 16'b0000000000000000;
    assign weights1[58][696] = 16'b0000000000000010;
    assign weights1[58][697] = 16'b0000000000000011;
    assign weights1[58][698] = 16'b1111111111111111;
    assign weights1[58][699] = 16'b1111111111111111;
    assign weights1[58][700] = 16'b0000000000000000;
    assign weights1[58][701] = 16'b1111111111111110;
    assign weights1[58][702] = 16'b0000000000000011;
    assign weights1[58][703] = 16'b0000000000000000;
    assign weights1[58][704] = 16'b0000000000000011;
    assign weights1[58][705] = 16'b1111111111110100;
    assign weights1[58][706] = 16'b1111111111110101;
    assign weights1[58][707] = 16'b1111111111101111;
    assign weights1[58][708] = 16'b1111111111100000;
    assign weights1[58][709] = 16'b1111111111101001;
    assign weights1[58][710] = 16'b1111111111011100;
    assign weights1[58][711] = 16'b1111111111010111;
    assign weights1[58][712] = 16'b1111111111110001;
    assign weights1[58][713] = 16'b1111111111111110;
    assign weights1[58][714] = 16'b1111111111101011;
    assign weights1[58][715] = 16'b1111111111101111;
    assign weights1[58][716] = 16'b1111111111100001;
    assign weights1[58][717] = 16'b1111111111100111;
    assign weights1[58][718] = 16'b1111111111110001;
    assign weights1[58][719] = 16'b1111111111101100;
    assign weights1[58][720] = 16'b1111111111110011;
    assign weights1[58][721] = 16'b1111111111111000;
    assign weights1[58][722] = 16'b1111111111111110;
    assign weights1[58][723] = 16'b0000000000000000;
    assign weights1[58][724] = 16'b0000000000000001;
    assign weights1[58][725] = 16'b0000000000000000;
    assign weights1[58][726] = 16'b1111111111111101;
    assign weights1[58][727] = 16'b1111111111111111;
    assign weights1[58][728] = 16'b0000000000000000;
    assign weights1[58][729] = 16'b1111111111111111;
    assign weights1[58][730] = 16'b0000000000000100;
    assign weights1[58][731] = 16'b0000000000001000;
    assign weights1[58][732] = 16'b0000000000000110;
    assign weights1[58][733] = 16'b0000000000000000;
    assign weights1[58][734] = 16'b0000000000000000;
    assign weights1[58][735] = 16'b1111111111111000;
    assign weights1[58][736] = 16'b1111111111111010;
    assign weights1[58][737] = 16'b1111111111101111;
    assign weights1[58][738] = 16'b1111111111110101;
    assign weights1[58][739] = 16'b1111111111100001;
    assign weights1[58][740] = 16'b1111111111110101;
    assign weights1[58][741] = 16'b1111111111111001;
    assign weights1[58][742] = 16'b1111111111110000;
    assign weights1[58][743] = 16'b1111111111110100;
    assign weights1[58][744] = 16'b1111111111111111;
    assign weights1[58][745] = 16'b1111111111110010;
    assign weights1[58][746] = 16'b1111111111110101;
    assign weights1[58][747] = 16'b1111111111111011;
    assign weights1[58][748] = 16'b1111111111111101;
    assign weights1[58][749] = 16'b1111111111111001;
    assign weights1[58][750] = 16'b1111111111111000;
    assign weights1[58][751] = 16'b1111111111111100;
    assign weights1[58][752] = 16'b1111111111111011;
    assign weights1[58][753] = 16'b1111111111111101;
    assign weights1[58][754] = 16'b0000000000000000;
    assign weights1[58][755] = 16'b0000000000000000;
    assign weights1[58][756] = 16'b0000000000000000;
    assign weights1[58][757] = 16'b0000000000000001;
    assign weights1[58][758] = 16'b0000000000000011;
    assign weights1[58][759] = 16'b0000000000000110;
    assign weights1[58][760] = 16'b0000000000001001;
    assign weights1[58][761] = 16'b0000000000000000;
    assign weights1[58][762] = 16'b0000000000000110;
    assign weights1[58][763] = 16'b0000000000001010;
    assign weights1[58][764] = 16'b0000000000000000;
    assign weights1[58][765] = 16'b0000000000000100;
    assign weights1[58][766] = 16'b1111111111110110;
    assign weights1[58][767] = 16'b1111111111111011;
    assign weights1[58][768] = 16'b0000000000000100;
    assign weights1[58][769] = 16'b1111111111110101;
    assign weights1[58][770] = 16'b1111111111110110;
    assign weights1[58][771] = 16'b1111111111111010;
    assign weights1[58][772] = 16'b1111111111101111;
    assign weights1[58][773] = 16'b1111111111101001;
    assign weights1[58][774] = 16'b1111111111111010;
    assign weights1[58][775] = 16'b1111111111111100;
    assign weights1[58][776] = 16'b1111111111111010;
    assign weights1[58][777] = 16'b1111111111111001;
    assign weights1[58][778] = 16'b1111111111111111;
    assign weights1[58][779] = 16'b1111111111111110;
    assign weights1[58][780] = 16'b1111111111111100;
    assign weights1[58][781] = 16'b1111111111111101;
    assign weights1[58][782] = 16'b1111111111111110;
    assign weights1[58][783] = 16'b0000000000000000;
    assign weights1[59][0] = 16'b0000000000000001;
    assign weights1[59][1] = 16'b0000000000000000;
    assign weights1[59][2] = 16'b1111111111111111;
    assign weights1[59][3] = 16'b1111111111111100;
    assign weights1[59][4] = 16'b1111111111111101;
    assign weights1[59][5] = 16'b1111111111111000;
    assign weights1[59][6] = 16'b1111111111110111;
    assign weights1[59][7] = 16'b1111111111110011;
    assign weights1[59][8] = 16'b1111111111111001;
    assign weights1[59][9] = 16'b1111111111111100;
    assign weights1[59][10] = 16'b1111111111111011;
    assign weights1[59][11] = 16'b1111111111110100;
    assign weights1[59][12] = 16'b0000000000000000;
    assign weights1[59][13] = 16'b1111111111111110;
    assign weights1[59][14] = 16'b1111111111111001;
    assign weights1[59][15] = 16'b0000000000000001;
    assign weights1[59][16] = 16'b1111111111110001;
    assign weights1[59][17] = 16'b0000000000001101;
    assign weights1[59][18] = 16'b0000000000001110;
    assign weights1[59][19] = 16'b0000000000010000;
    assign weights1[59][20] = 16'b0000000000011110;
    assign weights1[59][21] = 16'b0000000000001101;
    assign weights1[59][22] = 16'b0000000000010011;
    assign weights1[59][23] = 16'b0000000000001000;
    assign weights1[59][24] = 16'b0000000000000011;
    assign weights1[59][25] = 16'b0000000000000010;
    assign weights1[59][26] = 16'b0000000000000001;
    assign weights1[59][27] = 16'b0000000000000110;
    assign weights1[59][28] = 16'b0000000000000000;
    assign weights1[59][29] = 16'b1111111111111111;
    assign weights1[59][30] = 16'b1111111111111010;
    assign weights1[59][31] = 16'b1111111111111100;
    assign weights1[59][32] = 16'b1111111111111001;
    assign weights1[59][33] = 16'b0000000000001000;
    assign weights1[59][34] = 16'b1111111111110110;
    assign weights1[59][35] = 16'b1111111111111101;
    assign weights1[59][36] = 16'b0000000000000010;
    assign weights1[59][37] = 16'b1111111111111011;
    assign weights1[59][38] = 16'b1111111111100010;
    assign weights1[59][39] = 16'b0000000000000110;
    assign weights1[59][40] = 16'b0000000000001100;
    assign weights1[59][41] = 16'b0000000000010000;
    assign weights1[59][42] = 16'b0000000000001101;
    assign weights1[59][43] = 16'b0000000000000111;
    assign weights1[59][44] = 16'b1111111111110111;
    assign weights1[59][45] = 16'b0000000000010001;
    assign weights1[59][46] = 16'b0000000000010110;
    assign weights1[59][47] = 16'b0000000000001100;
    assign weights1[59][48] = 16'b0000000000001101;
    assign weights1[59][49] = 16'b0000000000011001;
    assign weights1[59][50] = 16'b0000000000011100;
    assign weights1[59][51] = 16'b0000000000001000;
    assign weights1[59][52] = 16'b0000000000000010;
    assign weights1[59][53] = 16'b0000000000001010;
    assign weights1[59][54] = 16'b0000000000001111;
    assign weights1[59][55] = 16'b0000000000000110;
    assign weights1[59][56] = 16'b0000000000000000;
    assign weights1[59][57] = 16'b1111111111111100;
    assign weights1[59][58] = 16'b1111111111111110;
    assign weights1[59][59] = 16'b0000000000000100;
    assign weights1[59][60] = 16'b0000000000001001;
    assign weights1[59][61] = 16'b0000000000001100;
    assign weights1[59][62] = 16'b0000000000001000;
    assign weights1[59][63] = 16'b1111111111111000;
    assign weights1[59][64] = 16'b0000000000000101;
    assign weights1[59][65] = 16'b0000000000000110;
    assign weights1[59][66] = 16'b0000000000000000;
    assign weights1[59][67] = 16'b0000000000000110;
    assign weights1[59][68] = 16'b0000000000001010;
    assign weights1[59][69] = 16'b0000000000000110;
    assign weights1[59][70] = 16'b1111111111110110;
    assign weights1[59][71] = 16'b1111111111110110;
    assign weights1[59][72] = 16'b0000000000010000;
    assign weights1[59][73] = 16'b0000000000010010;
    assign weights1[59][74] = 16'b0000000000010010;
    assign weights1[59][75] = 16'b0000000000011010;
    assign weights1[59][76] = 16'b0000000000001111;
    assign weights1[59][77] = 16'b0000000000010100;
    assign weights1[59][78] = 16'b0000000000011100;
    assign weights1[59][79] = 16'b0000000000100001;
    assign weights1[59][80] = 16'b0000000000011001;
    assign weights1[59][81] = 16'b0000000000100111;
    assign weights1[59][82] = 16'b0000000000011100;
    assign weights1[59][83] = 16'b0000000000001011;
    assign weights1[59][84] = 16'b1111111111111101;
    assign weights1[59][85] = 16'b1111111111110110;
    assign weights1[59][86] = 16'b1111111111111111;
    assign weights1[59][87] = 16'b0000000000001101;
    assign weights1[59][88] = 16'b0000000000010101;
    assign weights1[59][89] = 16'b0000000000011011;
    assign weights1[59][90] = 16'b0000000000100100;
    assign weights1[59][91] = 16'b0000000000010110;
    assign weights1[59][92] = 16'b0000000000011111;
    assign weights1[59][93] = 16'b0000000000011001;
    assign weights1[59][94] = 16'b0000000000010010;
    assign weights1[59][95] = 16'b0000000000010010;
    assign weights1[59][96] = 16'b0000000000010010;
    assign weights1[59][97] = 16'b0000000000010100;
    assign weights1[59][98] = 16'b0000000000010010;
    assign weights1[59][99] = 16'b0000000000010111;
    assign weights1[59][100] = 16'b0000000000010111;
    assign weights1[59][101] = 16'b0000000000011101;
    assign weights1[59][102] = 16'b0000000000101110;
    assign weights1[59][103] = 16'b0000000000001010;
    assign weights1[59][104] = 16'b0000000000010011;
    assign weights1[59][105] = 16'b0000000000101001;
    assign weights1[59][106] = 16'b0000000000100000;
    assign weights1[59][107] = 16'b0000000000011011;
    assign weights1[59][108] = 16'b0000000000101010;
    assign weights1[59][109] = 16'b0000000000100100;
    assign weights1[59][110] = 16'b0000000000010111;
    assign weights1[59][111] = 16'b0000000000010001;
    assign weights1[59][112] = 16'b1111111111111110;
    assign weights1[59][113] = 16'b1111111111111001;
    assign weights1[59][114] = 16'b0000000000000100;
    assign weights1[59][115] = 16'b0000000000010001;
    assign weights1[59][116] = 16'b0000000000100010;
    assign weights1[59][117] = 16'b0000000000100001;
    assign weights1[59][118] = 16'b0000000000100001;
    assign weights1[59][119] = 16'b0000000000100111;
    assign weights1[59][120] = 16'b0000000000110001;
    assign weights1[59][121] = 16'b0000000000111011;
    assign weights1[59][122] = 16'b0000000000101000;
    assign weights1[59][123] = 16'b0000000000100001;
    assign weights1[59][124] = 16'b0000000000101010;
    assign weights1[59][125] = 16'b0000000000100001;
    assign weights1[59][126] = 16'b0000000000011001;
    assign weights1[59][127] = 16'b0000000000001110;
    assign weights1[59][128] = 16'b0000000000111001;
    assign weights1[59][129] = 16'b0000000000010011;
    assign weights1[59][130] = 16'b0000000000010101;
    assign weights1[59][131] = 16'b0000000000101000;
    assign weights1[59][132] = 16'b0000000000101000;
    assign weights1[59][133] = 16'b0000000000100101;
    assign weights1[59][134] = 16'b0000000000110001;
    assign weights1[59][135] = 16'b0000000000100101;
    assign weights1[59][136] = 16'b0000000000100011;
    assign weights1[59][137] = 16'b0000000000010101;
    assign weights1[59][138] = 16'b0000000000010100;
    assign weights1[59][139] = 16'b0000000000010110;
    assign weights1[59][140] = 16'b0000000000001001;
    assign weights1[59][141] = 16'b0000000000001001;
    assign weights1[59][142] = 16'b0000000000010110;
    assign weights1[59][143] = 16'b0000000000010010;
    assign weights1[59][144] = 16'b0000000000101010;
    assign weights1[59][145] = 16'b0000000001000010;
    assign weights1[59][146] = 16'b0000000000100110;
    assign weights1[59][147] = 16'b0000000000101101;
    assign weights1[59][148] = 16'b0000000001000001;
    assign weights1[59][149] = 16'b0000000001000011;
    assign weights1[59][150] = 16'b0000000000111001;
    assign weights1[59][151] = 16'b0000000000110001;
    assign weights1[59][152] = 16'b0000000000100110;
    assign weights1[59][153] = 16'b0000000000001010;
    assign weights1[59][154] = 16'b0000000000101111;
    assign weights1[59][155] = 16'b0000000000100100;
    assign weights1[59][156] = 16'b0000000000011101;
    assign weights1[59][157] = 16'b0000000000010010;
    assign weights1[59][158] = 16'b0000000000101010;
    assign weights1[59][159] = 16'b0000000000100111;
    assign weights1[59][160] = 16'b0000000000100001;
    assign weights1[59][161] = 16'b0000000000011100;
    assign weights1[59][162] = 16'b0000000000110110;
    assign weights1[59][163] = 16'b0000000000010001;
    assign weights1[59][164] = 16'b0000000000001110;
    assign weights1[59][165] = 16'b0000000000001001;
    assign weights1[59][166] = 16'b0000000000011001;
    assign weights1[59][167] = 16'b0000000000001110;
    assign weights1[59][168] = 16'b0000000000010010;
    assign weights1[59][169] = 16'b0000000000011010;
    assign weights1[59][170] = 16'b0000000000011000;
    assign weights1[59][171] = 16'b0000000000101011;
    assign weights1[59][172] = 16'b0000000000101001;
    assign weights1[59][173] = 16'b0000000000110010;
    assign weights1[59][174] = 16'b0000000000101110;
    assign weights1[59][175] = 16'b0000000001000111;
    assign weights1[59][176] = 16'b0000000000101100;
    assign weights1[59][177] = 16'b0000000000111011;
    assign weights1[59][178] = 16'b0000000000111110;
    assign weights1[59][179] = 16'b0000000001000001;
    assign weights1[59][180] = 16'b0000000000100011;
    assign weights1[59][181] = 16'b0000000000100010;
    assign weights1[59][182] = 16'b0000000000111011;
    assign weights1[59][183] = 16'b0000000000011100;
    assign weights1[59][184] = 16'b0000000001000000;
    assign weights1[59][185] = 16'b0000000000011010;
    assign weights1[59][186] = 16'b0000000000011100;
    assign weights1[59][187] = 16'b0000000000011110;
    assign weights1[59][188] = 16'b0000000000010001;
    assign weights1[59][189] = 16'b0000000000110111;
    assign weights1[59][190] = 16'b0000000000011011;
    assign weights1[59][191] = 16'b0000000000101100;
    assign weights1[59][192] = 16'b0000000000010101;
    assign weights1[59][193] = 16'b0000000000000011;
    assign weights1[59][194] = 16'b0000000000011010;
    assign weights1[59][195] = 16'b0000000000010111;
    assign weights1[59][196] = 16'b0000000000011011;
    assign weights1[59][197] = 16'b0000000000101101;
    assign weights1[59][198] = 16'b0000000000011101;
    assign weights1[59][199] = 16'b0000000000100010;
    assign weights1[59][200] = 16'b0000000000100011;
    assign weights1[59][201] = 16'b0000000000011111;
    assign weights1[59][202] = 16'b0000000000100000;
    assign weights1[59][203] = 16'b0000000000100011;
    assign weights1[59][204] = 16'b0000000000011010;
    assign weights1[59][205] = 16'b0000000001010010;
    assign weights1[59][206] = 16'b0000000001010101;
    assign weights1[59][207] = 16'b0000000001000101;
    assign weights1[59][208] = 16'b0000000001000010;
    assign weights1[59][209] = 16'b0000000000111011;
    assign weights1[59][210] = 16'b0000000001001101;
    assign weights1[59][211] = 16'b0000000000110000;
    assign weights1[59][212] = 16'b0000000000100101;
    assign weights1[59][213] = 16'b0000000000110110;
    assign weights1[59][214] = 16'b0000000000100000;
    assign weights1[59][215] = 16'b0000000000010010;
    assign weights1[59][216] = 16'b0000000000001110;
    assign weights1[59][217] = 16'b0000000000001110;
    assign weights1[59][218] = 16'b0000000000101100;
    assign weights1[59][219] = 16'b0000000001000011;
    assign weights1[59][220] = 16'b0000000000110011;
    assign weights1[59][221] = 16'b0000000000010110;
    assign weights1[59][222] = 16'b0000000000010000;
    assign weights1[59][223] = 16'b0000000000010101;
    assign weights1[59][224] = 16'b0000000000100110;
    assign weights1[59][225] = 16'b0000000000101111;
    assign weights1[59][226] = 16'b0000000000011111;
    assign weights1[59][227] = 16'b0000000000011011;
    assign weights1[59][228] = 16'b0000000000010001;
    assign weights1[59][229] = 16'b0000000000101110;
    assign weights1[59][230] = 16'b0000000000100111;
    assign weights1[59][231] = 16'b0000000000011011;
    assign weights1[59][232] = 16'b0000000000101110;
    assign weights1[59][233] = 16'b0000000000110011;
    assign weights1[59][234] = 16'b0000000000101001;
    assign weights1[59][235] = 16'b0000000000011101;
    assign weights1[59][236] = 16'b0000000000011000;
    assign weights1[59][237] = 16'b0000000000101101;
    assign weights1[59][238] = 16'b0000000000101111;
    assign weights1[59][239] = 16'b0000000000100001;
    assign weights1[59][240] = 16'b0000000000100111;
    assign weights1[59][241] = 16'b0000000000010110;
    assign weights1[59][242] = 16'b0000000000010110;
    assign weights1[59][243] = 16'b0000000000100001;
    assign weights1[59][244] = 16'b0000000000001001;
    assign weights1[59][245] = 16'b0000000000001101;
    assign weights1[59][246] = 16'b0000000000011001;
    assign weights1[59][247] = 16'b0000000000101110;
    assign weights1[59][248] = 16'b0000000000110100;
    assign weights1[59][249] = 16'b0000000000101001;
    assign weights1[59][250] = 16'b0000000000010000;
    assign weights1[59][251] = 16'b0000000000011010;
    assign weights1[59][252] = 16'b0000000000100110;
    assign weights1[59][253] = 16'b0000000000101011;
    assign weights1[59][254] = 16'b0000000000100000;
    assign weights1[59][255] = 16'b0000000000010101;
    assign weights1[59][256] = 16'b0000000000001011;
    assign weights1[59][257] = 16'b0000000000010011;
    assign weights1[59][258] = 16'b0000000000010001;
    assign weights1[59][259] = 16'b0000000000001100;
    assign weights1[59][260] = 16'b0000000000010101;
    assign weights1[59][261] = 16'b0000000000111101;
    assign weights1[59][262] = 16'b0000000000000111;
    assign weights1[59][263] = 16'b1111111111010100;
    assign weights1[59][264] = 16'b1111111111010111;
    assign weights1[59][265] = 16'b0000000000000010;
    assign weights1[59][266] = 16'b1111111111111010;
    assign weights1[59][267] = 16'b1111111111100000;
    assign weights1[59][268] = 16'b1111111111101010;
    assign weights1[59][269] = 16'b1111111111110110;
    assign weights1[59][270] = 16'b1111111111011101;
    assign weights1[59][271] = 16'b1111111111111010;
    assign weights1[59][272] = 16'b1111111111110010;
    assign weights1[59][273] = 16'b0000000000000101;
    assign weights1[59][274] = 16'b0000000000010001;
    assign weights1[59][275] = 16'b0000000000101101;
    assign weights1[59][276] = 16'b0000000000101001;
    assign weights1[59][277] = 16'b0000000000100011;
    assign weights1[59][278] = 16'b0000000000100111;
    assign weights1[59][279] = 16'b0000000000010000;
    assign weights1[59][280] = 16'b0000000000100111;
    assign weights1[59][281] = 16'b0000000000101011;
    assign weights1[59][282] = 16'b0000000000010010;
    assign weights1[59][283] = 16'b0000000000010101;
    assign weights1[59][284] = 16'b0000000000001001;
    assign weights1[59][285] = 16'b0000000000010010;
    assign weights1[59][286] = 16'b1111111111110110;
    assign weights1[59][287] = 16'b0000000000010101;
    assign weights1[59][288] = 16'b0000000000010010;
    assign weights1[59][289] = 16'b0000000000001101;
    assign weights1[59][290] = 16'b1111111110111100;
    assign weights1[59][291] = 16'b1111111101111101;
    assign weights1[59][292] = 16'b1111111110101011;
    assign weights1[59][293] = 16'b1111111110111011;
    assign weights1[59][294] = 16'b1111111110111011;
    assign weights1[59][295] = 16'b1111111110111011;
    assign weights1[59][296] = 16'b1111111111010111;
    assign weights1[59][297] = 16'b1111111111010001;
    assign weights1[59][298] = 16'b1111111111111000;
    assign weights1[59][299] = 16'b1111111111111110;
    assign weights1[59][300] = 16'b1111111111110010;
    assign weights1[59][301] = 16'b0000000000000000;
    assign weights1[59][302] = 16'b0000000000011010;
    assign weights1[59][303] = 16'b0000000000101010;
    assign weights1[59][304] = 16'b0000000000011110;
    assign weights1[59][305] = 16'b0000000000101110;
    assign weights1[59][306] = 16'b0000000000101001;
    assign weights1[59][307] = 16'b0000000000001110;
    assign weights1[59][308] = 16'b0000000000100011;
    assign weights1[59][309] = 16'b0000000000101001;
    assign weights1[59][310] = 16'b0000000000011111;
    assign weights1[59][311] = 16'b0000000000001111;
    assign weights1[59][312] = 16'b0000000000000110;
    assign weights1[59][313] = 16'b0000000000000010;
    assign weights1[59][314] = 16'b0000000000000101;
    assign weights1[59][315] = 16'b0000000000010000;
    assign weights1[59][316] = 16'b0000000000001101;
    assign weights1[59][317] = 16'b1111111111100100;
    assign weights1[59][318] = 16'b1111111101111101;
    assign weights1[59][319] = 16'b1111111101111110;
    assign weights1[59][320] = 16'b1111111110111001;
    assign weights1[59][321] = 16'b1111111111010111;
    assign weights1[59][322] = 16'b1111111111100001;
    assign weights1[59][323] = 16'b1111111111010010;
    assign weights1[59][324] = 16'b1111111111001111;
    assign weights1[59][325] = 16'b1111111111001110;
    assign weights1[59][326] = 16'b1111111111000100;
    assign weights1[59][327] = 16'b1111111111011010;
    assign weights1[59][328] = 16'b1111111111101010;
    assign weights1[59][329] = 16'b1111111111101011;
    assign weights1[59][330] = 16'b1111111111111101;
    assign weights1[59][331] = 16'b0000000000101000;
    assign weights1[59][332] = 16'b0000000000100000;
    assign weights1[59][333] = 16'b0000000000100100;
    assign weights1[59][334] = 16'b0000000000110101;
    assign weights1[59][335] = 16'b0000000000010011;
    assign weights1[59][336] = 16'b0000000000011110;
    assign weights1[59][337] = 16'b0000000000100011;
    assign weights1[59][338] = 16'b0000000000011011;
    assign weights1[59][339] = 16'b0000000000000111;
    assign weights1[59][340] = 16'b1111111111111110;
    assign weights1[59][341] = 16'b1111111111111011;
    assign weights1[59][342] = 16'b0000000000010001;
    assign weights1[59][343] = 16'b1111111111101001;
    assign weights1[59][344] = 16'b1111111111111000;
    assign weights1[59][345] = 16'b1111111110110101;
    assign weights1[59][346] = 16'b1111111110011100;
    assign weights1[59][347] = 16'b1111111110111110;
    assign weights1[59][348] = 16'b1111111111101011;
    assign weights1[59][349] = 16'b1111111111101001;
    assign weights1[59][350] = 16'b1111111111001110;
    assign weights1[59][351] = 16'b1111111111010010;
    assign weights1[59][352] = 16'b1111111111100100;
    assign weights1[59][353] = 16'b1111111111001101;
    assign weights1[59][354] = 16'b1111111111011010;
    assign weights1[59][355] = 16'b1111111111010100;
    assign weights1[59][356] = 16'b1111111111101001;
    assign weights1[59][357] = 16'b1111111111101011;
    assign weights1[59][358] = 16'b1111111111100111;
    assign weights1[59][359] = 16'b0000000000010110;
    assign weights1[59][360] = 16'b0000000000010010;
    assign weights1[59][361] = 16'b0000000000010001;
    assign weights1[59][362] = 16'b0000000000010001;
    assign weights1[59][363] = 16'b0000000000001100;
    assign weights1[59][364] = 16'b0000000000010010;
    assign weights1[59][365] = 16'b0000000000011110;
    assign weights1[59][366] = 16'b0000000000011100;
    assign weights1[59][367] = 16'b0000000000001010;
    assign weights1[59][368] = 16'b1111111111111101;
    assign weights1[59][369] = 16'b1111111111111001;
    assign weights1[59][370] = 16'b1111111111111001;
    assign weights1[59][371] = 16'b1111111111101101;
    assign weights1[59][372] = 16'b1111111111011001;
    assign weights1[59][373] = 16'b1111111110111011;
    assign weights1[59][374] = 16'b1111111110011101;
    assign weights1[59][375] = 16'b1111111111010101;
    assign weights1[59][376] = 16'b1111111111110101;
    assign weights1[59][377] = 16'b1111111111011001;
    assign weights1[59][378] = 16'b1111111111001010;
    assign weights1[59][379] = 16'b1111111111101101;
    assign weights1[59][380] = 16'b1111111111011111;
    assign weights1[59][381] = 16'b1111111111001101;
    assign weights1[59][382] = 16'b1111111111101010;
    assign weights1[59][383] = 16'b1111111111001101;
    assign weights1[59][384] = 16'b1111111111011011;
    assign weights1[59][385] = 16'b1111111111010000;
    assign weights1[59][386] = 16'b1111111111110001;
    assign weights1[59][387] = 16'b0000000000000010;
    assign weights1[59][388] = 16'b0000000000000011;
    assign weights1[59][389] = 16'b0000000000000111;
    assign weights1[59][390] = 16'b0000000000000110;
    assign weights1[59][391] = 16'b0000000000000010;
    assign weights1[59][392] = 16'b0000000000001101;
    assign weights1[59][393] = 16'b0000000000001001;
    assign weights1[59][394] = 16'b0000000000010100;
    assign weights1[59][395] = 16'b0000000000001000;
    assign weights1[59][396] = 16'b1111111111111110;
    assign weights1[59][397] = 16'b0000000000001000;
    assign weights1[59][398] = 16'b1111111111101000;
    assign weights1[59][399] = 16'b1111111111111001;
    assign weights1[59][400] = 16'b1111111111100011;
    assign weights1[59][401] = 16'b1111111111011101;
    assign weights1[59][402] = 16'b1111111110111111;
    assign weights1[59][403] = 16'b1111111111101101;
    assign weights1[59][404] = 16'b1111111111111011;
    assign weights1[59][405] = 16'b1111111111101100;
    assign weights1[59][406] = 16'b1111111111111001;
    assign weights1[59][407] = 16'b0000000000010000;
    assign weights1[59][408] = 16'b1111111111011001;
    assign weights1[59][409] = 16'b1111111111111000;
    assign weights1[59][410] = 16'b1111111111110110;
    assign weights1[59][411] = 16'b1111111111011111;
    assign weights1[59][412] = 16'b1111111111100100;
    assign weights1[59][413] = 16'b1111111111110011;
    assign weights1[59][414] = 16'b0000000000000111;
    assign weights1[59][415] = 16'b1111111111110110;
    assign weights1[59][416] = 16'b1111111111111001;
    assign weights1[59][417] = 16'b1111111111111100;
    assign weights1[59][418] = 16'b1111111111111111;
    assign weights1[59][419] = 16'b0000000000000100;
    assign weights1[59][420] = 16'b1111111111111000;
    assign weights1[59][421] = 16'b0000000000000010;
    assign weights1[59][422] = 16'b0000000000000010;
    assign weights1[59][423] = 16'b0000000000001110;
    assign weights1[59][424] = 16'b1111111111111101;
    assign weights1[59][425] = 16'b1111111111111011;
    assign weights1[59][426] = 16'b0000000000000011;
    assign weights1[59][427] = 16'b1111111111101101;
    assign weights1[59][428] = 16'b1111111111110001;
    assign weights1[59][429] = 16'b1111111111010000;
    assign weights1[59][430] = 16'b1111111111100000;
    assign weights1[59][431] = 16'b1111111111011111;
    assign weights1[59][432] = 16'b1111111111101101;
    assign weights1[59][433] = 16'b1111111111100101;
    assign weights1[59][434] = 16'b1111111111101111;
    assign weights1[59][435] = 16'b1111111111101001;
    assign weights1[59][436] = 16'b1111111111110111;
    assign weights1[59][437] = 16'b1111111111011110;
    assign weights1[59][438] = 16'b1111111111100101;
    assign weights1[59][439] = 16'b1111111111111001;
    assign weights1[59][440] = 16'b1111111111110000;
    assign weights1[59][441] = 16'b1111111111111010;
    assign weights1[59][442] = 16'b1111111111101011;
    assign weights1[59][443] = 16'b1111111111110111;
    assign weights1[59][444] = 16'b1111111111100010;
    assign weights1[59][445] = 16'b1111111111111100;
    assign weights1[59][446] = 16'b1111111111111100;
    assign weights1[59][447] = 16'b1111111111110110;
    assign weights1[59][448] = 16'b1111111111101101;
    assign weights1[59][449] = 16'b1111111111111011;
    assign weights1[59][450] = 16'b1111111111101111;
    assign weights1[59][451] = 16'b1111111111111110;
    assign weights1[59][452] = 16'b0000000000000001;
    assign weights1[59][453] = 16'b0000000000000000;
    assign weights1[59][454] = 16'b1111111111101101;
    assign weights1[59][455] = 16'b1111111111110110;
    assign weights1[59][456] = 16'b1111111111011111;
    assign weights1[59][457] = 16'b1111111111100000;
    assign weights1[59][458] = 16'b1111111111010100;
    assign weights1[59][459] = 16'b1111111111110001;
    assign weights1[59][460] = 16'b1111111111110011;
    assign weights1[59][461] = 16'b0000000000001000;
    assign weights1[59][462] = 16'b1111111111110100;
    assign weights1[59][463] = 16'b0000000000000101;
    assign weights1[59][464] = 16'b1111111111111110;
    assign weights1[59][465] = 16'b1111111111101010;
    assign weights1[59][466] = 16'b0000000000001000;
    assign weights1[59][467] = 16'b1111111111101011;
    assign weights1[59][468] = 16'b1111111111001110;
    assign weights1[59][469] = 16'b1111111111110111;
    assign weights1[59][470] = 16'b1111111111101010;
    assign weights1[59][471] = 16'b1111111111111001;
    assign weights1[59][472] = 16'b1111111111101010;
    assign weights1[59][473] = 16'b1111111111101001;
    assign weights1[59][474] = 16'b1111111111100110;
    assign weights1[59][475] = 16'b1111111111100111;
    assign weights1[59][476] = 16'b1111111111110000;
    assign weights1[59][477] = 16'b1111111111101101;
    assign weights1[59][478] = 16'b1111111111110000;
    assign weights1[59][479] = 16'b1111111111110000;
    assign weights1[59][480] = 16'b1111111111101110;
    assign weights1[59][481] = 16'b1111111111111000;
    assign weights1[59][482] = 16'b1111111111101010;
    assign weights1[59][483] = 16'b1111111111111100;
    assign weights1[59][484] = 16'b1111111111110000;
    assign weights1[59][485] = 16'b1111111111110100;
    assign weights1[59][486] = 16'b1111111111100111;
    assign weights1[59][487] = 16'b0000000000000111;
    assign weights1[59][488] = 16'b0000000000000100;
    assign weights1[59][489] = 16'b1111111111110111;
    assign weights1[59][490] = 16'b1111111111111111;
    assign weights1[59][491] = 16'b0000000000000001;
    assign weights1[59][492] = 16'b1111111111110011;
    assign weights1[59][493] = 16'b1111111111011000;
    assign weights1[59][494] = 16'b1111111111100101;
    assign weights1[59][495] = 16'b1111111111011111;
    assign weights1[59][496] = 16'b1111111111110000;
    assign weights1[59][497] = 16'b1111111111111000;
    assign weights1[59][498] = 16'b1111111111101111;
    assign weights1[59][499] = 16'b1111111111110001;
    assign weights1[59][500] = 16'b1111111111010110;
    assign weights1[59][501] = 16'b1111111111100011;
    assign weights1[59][502] = 16'b1111111111011111;
    assign weights1[59][503] = 16'b1111111111100101;
    assign weights1[59][504] = 16'b1111111111111011;
    assign weights1[59][505] = 16'b1111111111111010;
    assign weights1[59][506] = 16'b1111111111110111;
    assign weights1[59][507] = 16'b1111111111111010;
    assign weights1[59][508] = 16'b1111111111011111;
    assign weights1[59][509] = 16'b1111111111111101;
    assign weights1[59][510] = 16'b1111111111110100;
    assign weights1[59][511] = 16'b1111111111110101;
    assign weights1[59][512] = 16'b1111111111100000;
    assign weights1[59][513] = 16'b1111111111110111;
    assign weights1[59][514] = 16'b1111111111100000;
    assign weights1[59][515] = 16'b1111111111100001;
    assign weights1[59][516] = 16'b0000000000000111;
    assign weights1[59][517] = 16'b0000000000000011;
    assign weights1[59][518] = 16'b1111111111110001;
    assign weights1[59][519] = 16'b0000000000000110;
    assign weights1[59][520] = 16'b1111111111101001;
    assign weights1[59][521] = 16'b1111111111100100;
    assign weights1[59][522] = 16'b1111111111011010;
    assign weights1[59][523] = 16'b1111111111101110;
    assign weights1[59][524] = 16'b1111111111110110;
    assign weights1[59][525] = 16'b1111111111100100;
    assign weights1[59][526] = 16'b1111111111111001;
    assign weights1[59][527] = 16'b1111111111101001;
    assign weights1[59][528] = 16'b1111111111110000;
    assign weights1[59][529] = 16'b1111111111100100;
    assign weights1[59][530] = 16'b1111111111100001;
    assign weights1[59][531] = 16'b1111111111101000;
    assign weights1[59][532] = 16'b1111111111111010;
    assign weights1[59][533] = 16'b1111111111111111;
    assign weights1[59][534] = 16'b0000000000000011;
    assign weights1[59][535] = 16'b1111111111110010;
    assign weights1[59][536] = 16'b1111111111110010;
    assign weights1[59][537] = 16'b1111111111100111;
    assign weights1[59][538] = 16'b1111111111100010;
    assign weights1[59][539] = 16'b1111111111111000;
    assign weights1[59][540] = 16'b1111111111101100;
    assign weights1[59][541] = 16'b1111111111110110;
    assign weights1[59][542] = 16'b0000000000000001;
    assign weights1[59][543] = 16'b1111111111100011;
    assign weights1[59][544] = 16'b1111111111110110;
    assign weights1[59][545] = 16'b1111111111101111;
    assign weights1[59][546] = 16'b1111111111101111;
    assign weights1[59][547] = 16'b1111111111111010;
    assign weights1[59][548] = 16'b1111111111100101;
    assign weights1[59][549] = 16'b1111111111101001;
    assign weights1[59][550] = 16'b1111111111101100;
    assign weights1[59][551] = 16'b1111111111100101;
    assign weights1[59][552] = 16'b1111111111101111;
    assign weights1[59][553] = 16'b1111111111111000;
    assign weights1[59][554] = 16'b1111111111110110;
    assign weights1[59][555] = 16'b1111111111101101;
    assign weights1[59][556] = 16'b1111111111100000;
    assign weights1[59][557] = 16'b1111111111101010;
    assign weights1[59][558] = 16'b1111111111101110;
    assign weights1[59][559] = 16'b1111111111110010;
    assign weights1[59][560] = 16'b1111111111111000;
    assign weights1[59][561] = 16'b1111111111111000;
    assign weights1[59][562] = 16'b1111111111110101;
    assign weights1[59][563] = 16'b0000000000001000;
    assign weights1[59][564] = 16'b1111111111100000;
    assign weights1[59][565] = 16'b0000000000000011;
    assign weights1[59][566] = 16'b0000000000001011;
    assign weights1[59][567] = 16'b1111111111110100;
    assign weights1[59][568] = 16'b1111111111111101;
    assign weights1[59][569] = 16'b1111111111111010;
    assign weights1[59][570] = 16'b1111111111011001;
    assign weights1[59][571] = 16'b1111111111111111;
    assign weights1[59][572] = 16'b1111111111110010;
    assign weights1[59][573] = 16'b0000000000000111;
    assign weights1[59][574] = 16'b1111111111110100;
    assign weights1[59][575] = 16'b1111111111100101;
    assign weights1[59][576] = 16'b1111111111101111;
    assign weights1[59][577] = 16'b1111111111111010;
    assign weights1[59][578] = 16'b1111111111100101;
    assign weights1[59][579] = 16'b1111111111100111;
    assign weights1[59][580] = 16'b1111111111111011;
    assign weights1[59][581] = 16'b1111111111111000;
    assign weights1[59][582] = 16'b1111111111101111;
    assign weights1[59][583] = 16'b1111111111011001;
    assign weights1[59][584] = 16'b1111111111001011;
    assign weights1[59][585] = 16'b1111111111100010;
    assign weights1[59][586] = 16'b1111111111101111;
    assign weights1[59][587] = 16'b1111111111111001;
    assign weights1[59][588] = 16'b1111111111111011;
    assign weights1[59][589] = 16'b0000000000000000;
    assign weights1[59][590] = 16'b1111111111111011;
    assign weights1[59][591] = 16'b1111111111111011;
    assign weights1[59][592] = 16'b1111111111101111;
    assign weights1[59][593] = 16'b1111111111101000;
    assign weights1[59][594] = 16'b1111111111111001;
    assign weights1[59][595] = 16'b1111111111110100;
    assign weights1[59][596] = 16'b1111111111011111;
    assign weights1[59][597] = 16'b1111111111111001;
    assign weights1[59][598] = 16'b0000000000000001;
    assign weights1[59][599] = 16'b0000000000000111;
    assign weights1[59][600] = 16'b0000000000000010;
    assign weights1[59][601] = 16'b0000000000001110;
    assign weights1[59][602] = 16'b1111111111100100;
    assign weights1[59][603] = 16'b1111111111001111;
    assign weights1[59][604] = 16'b1111111111011111;
    assign weights1[59][605] = 16'b1111111111100110;
    assign weights1[59][606] = 16'b1111111111010100;
    assign weights1[59][607] = 16'b0000000000000010;
    assign weights1[59][608] = 16'b1111111111111100;
    assign weights1[59][609] = 16'b1111111111100000;
    assign weights1[59][610] = 16'b1111111111011011;
    assign weights1[59][611] = 16'b1111111111010000;
    assign weights1[59][612] = 16'b1111111111100001;
    assign weights1[59][613] = 16'b1111111111101100;
    assign weights1[59][614] = 16'b1111111111110101;
    assign weights1[59][615] = 16'b1111111111111000;
    assign weights1[59][616] = 16'b1111111111111110;
    assign weights1[59][617] = 16'b1111111111111011;
    assign weights1[59][618] = 16'b1111111111111110;
    assign weights1[59][619] = 16'b1111111111101110;
    assign weights1[59][620] = 16'b1111111111110001;
    assign weights1[59][621] = 16'b1111111111110101;
    assign weights1[59][622] = 16'b1111111111100010;
    assign weights1[59][623] = 16'b1111111111101010;
    assign weights1[59][624] = 16'b1111111111111011;
    assign weights1[59][625] = 16'b1111111111110001;
    assign weights1[59][626] = 16'b1111111111110011;
    assign weights1[59][627] = 16'b1111111111111010;
    assign weights1[59][628] = 16'b0000000000000010;
    assign weights1[59][629] = 16'b0000000000001001;
    assign weights1[59][630] = 16'b1111111111101011;
    assign weights1[59][631] = 16'b1111111111101101;
    assign weights1[59][632] = 16'b1111111111111010;
    assign weights1[59][633] = 16'b1111111111100111;
    assign weights1[59][634] = 16'b1111111111110101;
    assign weights1[59][635] = 16'b1111111111110001;
    assign weights1[59][636] = 16'b1111111111100100;
    assign weights1[59][637] = 16'b1111111111010100;
    assign weights1[59][638] = 16'b1111111111010101;
    assign weights1[59][639] = 16'b1111111111011110;
    assign weights1[59][640] = 16'b1111111111100010;
    assign weights1[59][641] = 16'b1111111111101110;
    assign weights1[59][642] = 16'b1111111111111001;
    assign weights1[59][643] = 16'b1111111111111011;
    assign weights1[59][644] = 16'b1111111111111011;
    assign weights1[59][645] = 16'b1111111111111011;
    assign weights1[59][646] = 16'b1111111111110101;
    assign weights1[59][647] = 16'b1111111111111001;
    assign weights1[59][648] = 16'b1111111111110000;
    assign weights1[59][649] = 16'b1111111111100110;
    assign weights1[59][650] = 16'b0000000000001001;
    assign weights1[59][651] = 16'b1111111111101110;
    assign weights1[59][652] = 16'b1111111111110010;
    assign weights1[59][653] = 16'b1111111111110100;
    assign weights1[59][654] = 16'b0000000000001001;
    assign weights1[59][655] = 16'b1111111111001101;
    assign weights1[59][656] = 16'b1111111111101111;
    assign weights1[59][657] = 16'b1111111111101110;
    assign weights1[59][658] = 16'b1111111111101101;
    assign weights1[59][659] = 16'b1111111111010001;
    assign weights1[59][660] = 16'b1111111111101001;
    assign weights1[59][661] = 16'b1111111111011000;
    assign weights1[59][662] = 16'b1111111111010101;
    assign weights1[59][663] = 16'b1111111111010100;
    assign weights1[59][664] = 16'b1111111111001111;
    assign weights1[59][665] = 16'b1111111111010111;
    assign weights1[59][666] = 16'b1111111111011111;
    assign weights1[59][667] = 16'b1111111111011011;
    assign weights1[59][668] = 16'b1111111111100100;
    assign weights1[59][669] = 16'b1111111111110101;
    assign weights1[59][670] = 16'b1111111111111101;
    assign weights1[59][671] = 16'b1111111111111110;
    assign weights1[59][672] = 16'b1111111111111101;
    assign weights1[59][673] = 16'b0000000000000010;
    assign weights1[59][674] = 16'b1111111111111100;
    assign weights1[59][675] = 16'b1111111111110100;
    assign weights1[59][676] = 16'b1111111111101001;
    assign weights1[59][677] = 16'b1111111111110100;
    assign weights1[59][678] = 16'b1111111111110001;
    assign weights1[59][679] = 16'b1111111111110100;
    assign weights1[59][680] = 16'b0000000000000010;
    assign weights1[59][681] = 16'b1111111111110111;
    assign weights1[59][682] = 16'b1111111111111101;
    assign weights1[59][683] = 16'b1111111111111010;
    assign weights1[59][684] = 16'b1111111111101011;
    assign weights1[59][685] = 16'b1111111111111100;
    assign weights1[59][686] = 16'b1111111111010110;
    assign weights1[59][687] = 16'b1111111111100110;
    assign weights1[59][688] = 16'b1111111111001001;
    assign weights1[59][689] = 16'b1111111111001011;
    assign weights1[59][690] = 16'b1111111110111011;
    assign weights1[59][691] = 16'b1111111111000101;
    assign weights1[59][692] = 16'b1111111111010100;
    assign weights1[59][693] = 16'b1111111111010011;
    assign weights1[59][694] = 16'b1111111111011111;
    assign weights1[59][695] = 16'b1111111111101110;
    assign weights1[59][696] = 16'b1111111111110010;
    assign weights1[59][697] = 16'b1111111111111010;
    assign weights1[59][698] = 16'b1111111111111111;
    assign weights1[59][699] = 16'b1111111111111111;
    assign weights1[59][700] = 16'b1111111111111110;
    assign weights1[59][701] = 16'b1111111111111111;
    assign weights1[59][702] = 16'b1111111111111111;
    assign weights1[59][703] = 16'b1111111111111001;
    assign weights1[59][704] = 16'b1111111111110110;
    assign weights1[59][705] = 16'b1111111111110011;
    assign weights1[59][706] = 16'b0000000000000011;
    assign weights1[59][707] = 16'b1111111111111111;
    assign weights1[59][708] = 16'b0000000000000100;
    assign weights1[59][709] = 16'b0000000000010100;
    assign weights1[59][710] = 16'b0000000000001010;
    assign weights1[59][711] = 16'b1111111111111101;
    assign weights1[59][712] = 16'b1111111111101110;
    assign weights1[59][713] = 16'b1111111111111001;
    assign weights1[59][714] = 16'b1111111111101001;
    assign weights1[59][715] = 16'b1111111111101101;
    assign weights1[59][716] = 16'b1111111111010101;
    assign weights1[59][717] = 16'b1111111110111100;
    assign weights1[59][718] = 16'b1111111111010110;
    assign weights1[59][719] = 16'b1111111111010100;
    assign weights1[59][720] = 16'b1111111111100110;
    assign weights1[59][721] = 16'b1111111111110000;
    assign weights1[59][722] = 16'b1111111111101110;
    assign weights1[59][723] = 16'b1111111111110100;
    assign weights1[59][724] = 16'b1111111111110111;
    assign weights1[59][725] = 16'b1111111111111010;
    assign weights1[59][726] = 16'b1111111111111100;
    assign weights1[59][727] = 16'b0000000000000000;
    assign weights1[59][728] = 16'b0000000000000000;
    assign weights1[59][729] = 16'b1111111111111110;
    assign weights1[59][730] = 16'b0000000000000001;
    assign weights1[59][731] = 16'b1111111111111110;
    assign weights1[59][732] = 16'b1111111111111101;
    assign weights1[59][733] = 16'b1111111111110000;
    assign weights1[59][734] = 16'b1111111111111001;
    assign weights1[59][735] = 16'b1111111111111111;
    assign weights1[59][736] = 16'b1111111111111001;
    assign weights1[59][737] = 16'b1111111111111010;
    assign weights1[59][738] = 16'b1111111111111111;
    assign weights1[59][739] = 16'b0000000000000100;
    assign weights1[59][740] = 16'b1111111111111111;
    assign weights1[59][741] = 16'b0000000000000100;
    assign weights1[59][742] = 16'b1111111111111001;
    assign weights1[59][743] = 16'b1111111111111011;
    assign weights1[59][744] = 16'b1111111111110011;
    assign weights1[59][745] = 16'b1111111111101011;
    assign weights1[59][746] = 16'b1111111111100101;
    assign weights1[59][747] = 16'b1111111111110000;
    assign weights1[59][748] = 16'b1111111111110100;
    assign weights1[59][749] = 16'b1111111111110101;
    assign weights1[59][750] = 16'b1111111111110011;
    assign weights1[59][751] = 16'b1111111111110111;
    assign weights1[59][752] = 16'b1111111111111001;
    assign weights1[59][753] = 16'b1111111111111101;
    assign weights1[59][754] = 16'b1111111111111111;
    assign weights1[59][755] = 16'b0000000000000000;
    assign weights1[59][756] = 16'b0000000000000000;
    assign weights1[59][757] = 16'b0000000000000000;
    assign weights1[59][758] = 16'b0000000000000000;
    assign weights1[59][759] = 16'b1111111111111110;
    assign weights1[59][760] = 16'b1111111111111100;
    assign weights1[59][761] = 16'b1111111111111001;
    assign weights1[59][762] = 16'b1111111111111110;
    assign weights1[59][763] = 16'b0000000000001000;
    assign weights1[59][764] = 16'b1111111111111100;
    assign weights1[59][765] = 16'b0000000000000010;
    assign weights1[59][766] = 16'b1111111111111101;
    assign weights1[59][767] = 16'b1111111111111110;
    assign weights1[59][768] = 16'b1111111111111110;
    assign weights1[59][769] = 16'b0000000000000100;
    assign weights1[59][770] = 16'b1111111111111101;
    assign weights1[59][771] = 16'b1111111111110111;
    assign weights1[59][772] = 16'b1111111111110011;
    assign weights1[59][773] = 16'b1111111111110111;
    assign weights1[59][774] = 16'b1111111111110111;
    assign weights1[59][775] = 16'b1111111111110111;
    assign weights1[59][776] = 16'b1111111111110111;
    assign weights1[59][777] = 16'b1111111111110110;
    assign weights1[59][778] = 16'b1111111111111000;
    assign weights1[59][779] = 16'b1111111111111101;
    assign weights1[59][780] = 16'b1111111111111110;
    assign weights1[59][781] = 16'b1111111111111110;
    assign weights1[59][782] = 16'b1111111111111110;
    assign weights1[59][783] = 16'b1111111111111111;
    assign weights1[60][0] = 16'b0000000000000000;
    assign weights1[60][1] = 16'b0000000000000000;
    assign weights1[60][2] = 16'b1111111111111110;
    assign weights1[60][3] = 16'b1111111111111011;
    assign weights1[60][4] = 16'b1111111111111000;
    assign weights1[60][5] = 16'b1111111111110110;
    assign weights1[60][6] = 16'b1111111111110010;
    assign weights1[60][7] = 16'b1111111111110000;
    assign weights1[60][8] = 16'b1111111111101111;
    assign weights1[60][9] = 16'b1111111111101100;
    assign weights1[60][10] = 16'b1111111111101011;
    assign weights1[60][11] = 16'b1111111111110111;
    assign weights1[60][12] = 16'b1111111111110111;
    assign weights1[60][13] = 16'b1111111111110101;
    assign weights1[60][14] = 16'b1111111111110111;
    assign weights1[60][15] = 16'b1111111111110111;
    assign weights1[60][16] = 16'b1111111111110110;
    assign weights1[60][17] = 16'b1111111111110110;
    assign weights1[60][18] = 16'b1111111111110101;
    assign weights1[60][19] = 16'b1111111111110111;
    assign weights1[60][20] = 16'b1111111111111001;
    assign weights1[60][21] = 16'b1111111111111101;
    assign weights1[60][22] = 16'b0000000000000010;
    assign weights1[60][23] = 16'b1111111111111111;
    assign weights1[60][24] = 16'b0000000000000001;
    assign weights1[60][25] = 16'b1111111111111111;
    assign weights1[60][26] = 16'b1111111111111111;
    assign weights1[60][27] = 16'b0000000000000000;
    assign weights1[60][28] = 16'b0000000000000000;
    assign weights1[60][29] = 16'b0000000000000000;
    assign weights1[60][30] = 16'b1111111111111100;
    assign weights1[60][31] = 16'b1111111111111001;
    assign weights1[60][32] = 16'b1111111111110010;
    assign weights1[60][33] = 16'b1111111111101101;
    assign weights1[60][34] = 16'b1111111111101001;
    assign weights1[60][35] = 16'b1111111111100100;
    assign weights1[60][36] = 16'b1111111111100111;
    assign weights1[60][37] = 16'b1111111111100000;
    assign weights1[60][38] = 16'b1111111111100001;
    assign weights1[60][39] = 16'b1111111111101110;
    assign weights1[60][40] = 16'b1111111111100110;
    assign weights1[60][41] = 16'b1111111111100101;
    assign weights1[60][42] = 16'b1111111111101001;
    assign weights1[60][43] = 16'b1111111111101110;
    assign weights1[60][44] = 16'b1111111111110100;
    assign weights1[60][45] = 16'b1111111111100110;
    assign weights1[60][46] = 16'b1111111111110000;
    assign weights1[60][47] = 16'b1111111111110100;
    assign weights1[60][48] = 16'b1111111111111001;
    assign weights1[60][49] = 16'b1111111111110110;
    assign weights1[60][50] = 16'b1111111111111001;
    assign weights1[60][51] = 16'b1111111111111010;
    assign weights1[60][52] = 16'b1111111111111100;
    assign weights1[60][53] = 16'b1111111111111101;
    assign weights1[60][54] = 16'b1111111111111101;
    assign weights1[60][55] = 16'b0000000000000000;
    assign weights1[60][56] = 16'b1111111111111110;
    assign weights1[60][57] = 16'b1111111111111110;
    assign weights1[60][58] = 16'b1111111111111001;
    assign weights1[60][59] = 16'b1111111111110000;
    assign weights1[60][60] = 16'b1111111111100101;
    assign weights1[60][61] = 16'b1111111111100011;
    assign weights1[60][62] = 16'b1111111111011010;
    assign weights1[60][63] = 16'b1111111111010111;
    assign weights1[60][64] = 16'b1111111111011100;
    assign weights1[60][65] = 16'b1111111111001110;
    assign weights1[60][66] = 16'b1111111111010011;
    assign weights1[60][67] = 16'b1111111111001110;
    assign weights1[60][68] = 16'b1111111111010101;
    assign weights1[60][69] = 16'b1111111111011001;
    assign weights1[60][70] = 16'b1111111111011010;
    assign weights1[60][71] = 16'b1111111111011011;
    assign weights1[60][72] = 16'b1111111111100001;
    assign weights1[60][73] = 16'b1111111111011111;
    assign weights1[60][74] = 16'b1111111111010111;
    assign weights1[60][75] = 16'b1111111111101001;
    assign weights1[60][76] = 16'b1111111111101001;
    assign weights1[60][77] = 16'b1111111111101010;
    assign weights1[60][78] = 16'b1111111111110011;
    assign weights1[60][79] = 16'b1111111111110111;
    assign weights1[60][80] = 16'b1111111111110110;
    assign weights1[60][81] = 16'b1111111111111000;
    assign weights1[60][82] = 16'b1111111111111100;
    assign weights1[60][83] = 16'b1111111111111101;
    assign weights1[60][84] = 16'b1111111111111111;
    assign weights1[60][85] = 16'b1111111111111011;
    assign weights1[60][86] = 16'b1111111111110101;
    assign weights1[60][87] = 16'b1111111111100101;
    assign weights1[60][88] = 16'b1111111111010111;
    assign weights1[60][89] = 16'b1111111111001110;
    assign weights1[60][90] = 16'b1111111110111100;
    assign weights1[60][91] = 16'b1111111110111110;
    assign weights1[60][92] = 16'b1111111110111111;
    assign weights1[60][93] = 16'b1111111110101101;
    assign weights1[60][94] = 16'b1111111110011010;
    assign weights1[60][95] = 16'b1111111110110000;
    assign weights1[60][96] = 16'b1111111110111101;
    assign weights1[60][97] = 16'b1111111110110100;
    assign weights1[60][98] = 16'b1111111110110001;
    assign weights1[60][99] = 16'b1111111110111100;
    assign weights1[60][100] = 16'b1111111111000100;
    assign weights1[60][101] = 16'b1111111111000110;
    assign weights1[60][102] = 16'b1111111111001100;
    assign weights1[60][103] = 16'b1111111111010000;
    assign weights1[60][104] = 16'b1111111111010111;
    assign weights1[60][105] = 16'b1111111111010100;
    assign weights1[60][106] = 16'b1111111111101101;
    assign weights1[60][107] = 16'b1111111111101001;
    assign weights1[60][108] = 16'b1111111111101101;
    assign weights1[60][109] = 16'b1111111111111000;
    assign weights1[60][110] = 16'b1111111111111010;
    assign weights1[60][111] = 16'b1111111111111010;
    assign weights1[60][112] = 16'b1111111111111110;
    assign weights1[60][113] = 16'b1111111111110010;
    assign weights1[60][114] = 16'b1111111111101010;
    assign weights1[60][115] = 16'b1111111111100000;
    assign weights1[60][116] = 16'b1111111111010000;
    assign weights1[60][117] = 16'b1111111110111010;
    assign weights1[60][118] = 16'b1111111110101110;
    assign weights1[60][119] = 16'b1111111110100000;
    assign weights1[60][120] = 16'b1111111110100011;
    assign weights1[60][121] = 16'b1111111110010110;
    assign weights1[60][122] = 16'b1111111110000100;
    assign weights1[60][123] = 16'b1111111110001010;
    assign weights1[60][124] = 16'b1111111110010100;
    assign weights1[60][125] = 16'b1111111110010010;
    assign weights1[60][126] = 16'b1111111110011011;
    assign weights1[60][127] = 16'b1111111110100110;
    assign weights1[60][128] = 16'b1111111110110011;
    assign weights1[60][129] = 16'b1111111110101110;
    assign weights1[60][130] = 16'b1111111110101010;
    assign weights1[60][131] = 16'b1111111110110111;
    assign weights1[60][132] = 16'b1111111110111110;
    assign weights1[60][133] = 16'b1111111111001010;
    assign weights1[60][134] = 16'b1111111111001010;
    assign weights1[60][135] = 16'b1111111111011000;
    assign weights1[60][136] = 16'b1111111111011111;
    assign weights1[60][137] = 16'b1111111111100001;
    assign weights1[60][138] = 16'b1111111111110000;
    assign weights1[60][139] = 16'b1111111111110001;
    assign weights1[60][140] = 16'b1111111111111011;
    assign weights1[60][141] = 16'b1111111111110111;
    assign weights1[60][142] = 16'b1111111111100111;
    assign weights1[60][143] = 16'b1111111111011100;
    assign weights1[60][144] = 16'b1111111111010100;
    assign weights1[60][145] = 16'b1111111110111001;
    assign weights1[60][146] = 16'b1111111110100110;
    assign weights1[60][147] = 16'b1111111110101101;
    assign weights1[60][148] = 16'b1111111110101011;
    assign weights1[60][149] = 16'b1111111110010010;
    assign weights1[60][150] = 16'b1111111110000000;
    assign weights1[60][151] = 16'b1111111110000011;
    assign weights1[60][152] = 16'b1111111110011101;
    assign weights1[60][153] = 16'b1111111110010010;
    assign weights1[60][154] = 16'b1111111110010111;
    assign weights1[60][155] = 16'b1111111111000010;
    assign weights1[60][156] = 16'b1111111110000110;
    assign weights1[60][157] = 16'b1111111110010100;
    assign weights1[60][158] = 16'b1111111110100000;
    assign weights1[60][159] = 16'b1111111110011001;
    assign weights1[60][160] = 16'b1111111110001011;
    assign weights1[60][161] = 16'b1111111110100010;
    assign weights1[60][162] = 16'b1111111110111000;
    assign weights1[60][163] = 16'b1111111110101100;
    assign weights1[60][164] = 16'b1111111110111110;
    assign weights1[60][165] = 16'b1111111111010110;
    assign weights1[60][166] = 16'b1111111111011010;
    assign weights1[60][167] = 16'b1111111111101011;
    assign weights1[60][168] = 16'b1111111111111011;
    assign weights1[60][169] = 16'b1111111111111010;
    assign weights1[60][170] = 16'b1111111111110011;
    assign weights1[60][171] = 16'b1111111111110110;
    assign weights1[60][172] = 16'b1111111111111010;
    assign weights1[60][173] = 16'b1111111111101011;
    assign weights1[60][174] = 16'b1111111111101111;
    assign weights1[60][175] = 16'b1111111111001001;
    assign weights1[60][176] = 16'b1111111111010000;
    assign weights1[60][177] = 16'b1111111111011101;
    assign weights1[60][178] = 16'b1111111111011101;
    assign weights1[60][179] = 16'b1111111111011110;
    assign weights1[60][180] = 16'b1111111111000101;
    assign weights1[60][181] = 16'b1111111110111101;
    assign weights1[60][182] = 16'b1111111111000100;
    assign weights1[60][183] = 16'b1111111110101101;
    assign weights1[60][184] = 16'b1111111110110111;
    assign weights1[60][185] = 16'b1111111111100011;
    assign weights1[60][186] = 16'b1111111110111100;
    assign weights1[60][187] = 16'b1111111110110100;
    assign weights1[60][188] = 16'b1111111110101010;
    assign weights1[60][189] = 16'b1111111111010110;
    assign weights1[60][190] = 16'b1111111111000111;
    assign weights1[60][191] = 16'b1111111110111001;
    assign weights1[60][192] = 16'b1111111111001011;
    assign weights1[60][193] = 16'b1111111111011000;
    assign weights1[60][194] = 16'b1111111111011110;
    assign weights1[60][195] = 16'b1111111111101011;
    assign weights1[60][196] = 16'b0000000000000001;
    assign weights1[60][197] = 16'b1111111111111110;
    assign weights1[60][198] = 16'b1111111111111101;
    assign weights1[60][199] = 16'b1111111111110100;
    assign weights1[60][200] = 16'b0000000000001100;
    assign weights1[60][201] = 16'b0000000000001110;
    assign weights1[60][202] = 16'b0000000000011111;
    assign weights1[60][203] = 16'b0000000000100101;
    assign weights1[60][204] = 16'b0000000000011001;
    assign weights1[60][205] = 16'b0000000000011101;
    assign weights1[60][206] = 16'b0000000000001000;
    assign weights1[60][207] = 16'b0000000000000001;
    assign weights1[60][208] = 16'b1111111111111001;
    assign weights1[60][209] = 16'b1111111111101111;
    assign weights1[60][210] = 16'b0000000000001111;
    assign weights1[60][211] = 16'b1111111111100000;
    assign weights1[60][212] = 16'b1111111111101100;
    assign weights1[60][213] = 16'b1111111111110110;
    assign weights1[60][214] = 16'b1111111111100111;
    assign weights1[60][215] = 16'b1111111111110110;
    assign weights1[60][216] = 16'b1111111111101011;
    assign weights1[60][217] = 16'b1111111111101100;
    assign weights1[60][218] = 16'b1111111111111001;
    assign weights1[60][219] = 16'b0000000000001010;
    assign weights1[60][220] = 16'b0000000000000010;
    assign weights1[60][221] = 16'b1111111111100100;
    assign weights1[60][222] = 16'b1111111111110111;
    assign weights1[60][223] = 16'b1111111111111011;
    assign weights1[60][224] = 16'b1111111111111100;
    assign weights1[60][225] = 16'b1111111111111110;
    assign weights1[60][226] = 16'b1111111111111101;
    assign weights1[60][227] = 16'b0000000000000000;
    assign weights1[60][228] = 16'b0000000000000101;
    assign weights1[60][229] = 16'b0000000000100011;
    assign weights1[60][230] = 16'b0000000000001001;
    assign weights1[60][231] = 16'b0000000000110110;
    assign weights1[60][232] = 16'b0000000000110000;
    assign weights1[60][233] = 16'b0000000000100100;
    assign weights1[60][234] = 16'b0000000000101100;
    assign weights1[60][235] = 16'b0000000000100111;
    assign weights1[60][236] = 16'b0000000000110001;
    assign weights1[60][237] = 16'b0000000000010111;
    assign weights1[60][238] = 16'b0000000000010000;
    assign weights1[60][239] = 16'b0000000000001110;
    assign weights1[60][240] = 16'b1111111111111110;
    assign weights1[60][241] = 16'b0000000000010101;
    assign weights1[60][242] = 16'b0000000000010101;
    assign weights1[60][243] = 16'b0000000000010101;
    assign weights1[60][244] = 16'b0000000000100010;
    assign weights1[60][245] = 16'b0000000000011001;
    assign weights1[60][246] = 16'b0000000000001110;
    assign weights1[60][247] = 16'b0000000000100000;
    assign weights1[60][248] = 16'b0000000000011100;
    assign weights1[60][249] = 16'b0000000000100000;
    assign weights1[60][250] = 16'b0000000000001111;
    assign weights1[60][251] = 16'b0000000000001110;
    assign weights1[60][252] = 16'b0000000000000011;
    assign weights1[60][253] = 16'b0000000000000100;
    assign weights1[60][254] = 16'b0000000000000111;
    assign weights1[60][255] = 16'b0000000000000101;
    assign weights1[60][256] = 16'b0000000000000001;
    assign weights1[60][257] = 16'b0000000000010011;
    assign weights1[60][258] = 16'b0000000000010111;
    assign weights1[60][259] = 16'b0000000000010101;
    assign weights1[60][260] = 16'b0000000000101101;
    assign weights1[60][261] = 16'b0000000000111100;
    assign weights1[60][262] = 16'b0000000000110101;
    assign weights1[60][263] = 16'b0000000000101110;
    assign weights1[60][264] = 16'b0000000001000010;
    assign weights1[60][265] = 16'b0000000000011111;
    assign weights1[60][266] = 16'b0000000000100101;
    assign weights1[60][267] = 16'b0000000000010001;
    assign weights1[60][268] = 16'b0000000000100101;
    assign weights1[60][269] = 16'b0000000000011001;
    assign weights1[60][270] = 16'b0000000000010001;
    assign weights1[60][271] = 16'b0000000000010100;
    assign weights1[60][272] = 16'b0000000000010111;
    assign weights1[60][273] = 16'b0000000000001110;
    assign weights1[60][274] = 16'b0000000000011010;
    assign weights1[60][275] = 16'b1111111111111110;
    assign weights1[60][276] = 16'b0000000000100100;
    assign weights1[60][277] = 16'b0000000000011101;
    assign weights1[60][278] = 16'b0000000000000100;
    assign weights1[60][279] = 16'b0000000000010100;
    assign weights1[60][280] = 16'b0000000000001000;
    assign weights1[60][281] = 16'b0000000000000100;
    assign weights1[60][282] = 16'b0000000000000100;
    assign weights1[60][283] = 16'b1111111111111110;
    assign weights1[60][284] = 16'b0000000000000110;
    assign weights1[60][285] = 16'b1111111111111110;
    assign weights1[60][286] = 16'b0000000000010010;
    assign weights1[60][287] = 16'b0000000000001001;
    assign weights1[60][288] = 16'b0000000000001111;
    assign weights1[60][289] = 16'b0000000000011111;
    assign weights1[60][290] = 16'b0000000000011101;
    assign weights1[60][291] = 16'b0000000000101010;
    assign weights1[60][292] = 16'b0000000000101001;
    assign weights1[60][293] = 16'b0000000001011001;
    assign weights1[60][294] = 16'b0000000000111100;
    assign weights1[60][295] = 16'b0000000001000101;
    assign weights1[60][296] = 16'b0000000000111010;
    assign weights1[60][297] = 16'b0000000000100010;
    assign weights1[60][298] = 16'b0000000000110001;
    assign weights1[60][299] = 16'b0000000000101100;
    assign weights1[60][300] = 16'b0000000000001001;
    assign weights1[60][301] = 16'b0000000000010110;
    assign weights1[60][302] = 16'b0000000000001000;
    assign weights1[60][303] = 16'b0000000000010101;
    assign weights1[60][304] = 16'b0000000000001110;
    assign weights1[60][305] = 16'b0000000000001110;
    assign weights1[60][306] = 16'b0000000000001110;
    assign weights1[60][307] = 16'b0000000000001100;
    assign weights1[60][308] = 16'b0000000000000111;
    assign weights1[60][309] = 16'b0000000000000011;
    assign weights1[60][310] = 16'b0000000000001010;
    assign weights1[60][311] = 16'b1111111111110111;
    assign weights1[60][312] = 16'b1111111111110110;
    assign weights1[60][313] = 16'b1111111111100110;
    assign weights1[60][314] = 16'b0000000000000111;
    assign weights1[60][315] = 16'b0000000000000101;
    assign weights1[60][316] = 16'b1111111111101110;
    assign weights1[60][317] = 16'b0000000000001000;
    assign weights1[60][318] = 16'b1111111111110100;
    assign weights1[60][319] = 16'b0000000000100000;
    assign weights1[60][320] = 16'b0000000000011100;
    assign weights1[60][321] = 16'b0000000000100110;
    assign weights1[60][322] = 16'b0000000000111000;
    assign weights1[60][323] = 16'b0000000000111011;
    assign weights1[60][324] = 16'b0000000000111010;
    assign weights1[60][325] = 16'b0000000000111010;
    assign weights1[60][326] = 16'b0000000000011100;
    assign weights1[60][327] = 16'b0000000000111000;
    assign weights1[60][328] = 16'b0000000000100000;
    assign weights1[60][329] = 16'b0000000000001010;
    assign weights1[60][330] = 16'b0000000000011010;
    assign weights1[60][331] = 16'b0000000000000100;
    assign weights1[60][332] = 16'b1111111111111111;
    assign weights1[60][333] = 16'b0000000000001010;
    assign weights1[60][334] = 16'b1111111111111101;
    assign weights1[60][335] = 16'b0000000000001000;
    assign weights1[60][336] = 16'b0000000000000011;
    assign weights1[60][337] = 16'b1111111111110111;
    assign weights1[60][338] = 16'b0000000000000010;
    assign weights1[60][339] = 16'b1111111111110111;
    assign weights1[60][340] = 16'b1111111111110110;
    assign weights1[60][341] = 16'b1111111111101110;
    assign weights1[60][342] = 16'b0000000000001101;
    assign weights1[60][343] = 16'b1111111111110001;
    assign weights1[60][344] = 16'b1111111111111001;
    assign weights1[60][345] = 16'b1111111111110000;
    assign weights1[60][346] = 16'b1111111111101110;
    assign weights1[60][347] = 16'b1111111111101101;
    assign weights1[60][348] = 16'b1111111111011100;
    assign weights1[60][349] = 16'b1111111111110110;
    assign weights1[60][350] = 16'b0000000000001100;
    assign weights1[60][351] = 16'b0000000000010010;
    assign weights1[60][352] = 16'b0000000000011011;
    assign weights1[60][353] = 16'b1111111111111101;
    assign weights1[60][354] = 16'b1111111111111101;
    assign weights1[60][355] = 16'b0000000000010110;
    assign weights1[60][356] = 16'b0000000000000001;
    assign weights1[60][357] = 16'b1111111111101101;
    assign weights1[60][358] = 16'b0000000000000000;
    assign weights1[60][359] = 16'b1111111111111001;
    assign weights1[60][360] = 16'b1111111111111001;
    assign weights1[60][361] = 16'b0000000000010010;
    assign weights1[60][362] = 16'b1111111111110000;
    assign weights1[60][363] = 16'b1111111111111101;
    assign weights1[60][364] = 16'b0000000000000111;
    assign weights1[60][365] = 16'b1111111111110001;
    assign weights1[60][366] = 16'b0000000000001110;
    assign weights1[60][367] = 16'b1111111111110100;
    assign weights1[60][368] = 16'b1111111111110011;
    assign weights1[60][369] = 16'b1111111111111010;
    assign weights1[60][370] = 16'b1111111111111111;
    assign weights1[60][371] = 16'b1111111111111001;
    assign weights1[60][372] = 16'b1111111111111101;
    assign weights1[60][373] = 16'b1111111111111111;
    assign weights1[60][374] = 16'b1111111111101110;
    assign weights1[60][375] = 16'b1111111111101110;
    assign weights1[60][376] = 16'b1111111111101010;
    assign weights1[60][377] = 16'b1111111111100100;
    assign weights1[60][378] = 16'b1111111111010100;
    assign weights1[60][379] = 16'b1111111111100110;
    assign weights1[60][380] = 16'b1111111111101011;
    assign weights1[60][381] = 16'b1111111111110100;
    assign weights1[60][382] = 16'b1111111111111001;
    assign weights1[60][383] = 16'b1111111111101000;
    assign weights1[60][384] = 16'b1111111111101010;
    assign weights1[60][385] = 16'b0000000000001101;
    assign weights1[60][386] = 16'b0000000000001001;
    assign weights1[60][387] = 16'b1111111111111101;
    assign weights1[60][388] = 16'b1111111111101000;
    assign weights1[60][389] = 16'b0000000000000010;
    assign weights1[60][390] = 16'b1111111111111101;
    assign weights1[60][391] = 16'b1111111111111101;
    assign weights1[60][392] = 16'b0000000000000000;
    assign weights1[60][393] = 16'b1111111111110111;
    assign weights1[60][394] = 16'b0000000000000000;
    assign weights1[60][395] = 16'b0000000000011010;
    assign weights1[60][396] = 16'b0000000000000000;
    assign weights1[60][397] = 16'b1111111111111010;
    assign weights1[60][398] = 16'b1111111111111111;
    assign weights1[60][399] = 16'b1111111111111111;
    assign weights1[60][400] = 16'b1111111111111110;
    assign weights1[60][401] = 16'b1111111111110101;
    assign weights1[60][402] = 16'b0000000000000100;
    assign weights1[60][403] = 16'b0000000000000010;
    assign weights1[60][404] = 16'b1111111111101011;
    assign weights1[60][405] = 16'b1111111111101101;
    assign weights1[60][406] = 16'b1111111111100111;
    assign weights1[60][407] = 16'b1111111111010010;
    assign weights1[60][408] = 16'b1111111111100101;
    assign weights1[60][409] = 16'b0000000000001101;
    assign weights1[60][410] = 16'b1111111111101111;
    assign weights1[60][411] = 16'b1111111111111010;
    assign weights1[60][412] = 16'b0000000000000000;
    assign weights1[60][413] = 16'b1111111111110110;
    assign weights1[60][414] = 16'b1111111111111111;
    assign weights1[60][415] = 16'b0000000000001001;
    assign weights1[60][416] = 16'b0000000000010011;
    assign weights1[60][417] = 16'b1111111111101111;
    assign weights1[60][418] = 16'b1111111111111010;
    assign weights1[60][419] = 16'b1111111111111011;
    assign weights1[60][420] = 16'b0000000000000010;
    assign weights1[60][421] = 16'b0000000000000011;
    assign weights1[60][422] = 16'b1111111111111111;
    assign weights1[60][423] = 16'b0000000000100000;
    assign weights1[60][424] = 16'b0000000000100000;
    assign weights1[60][425] = 16'b1111111111111001;
    assign weights1[60][426] = 16'b0000000000011110;
    assign weights1[60][427] = 16'b0000000000010101;
    assign weights1[60][428] = 16'b1111111111110111;
    assign weights1[60][429] = 16'b0000000000000100;
    assign weights1[60][430] = 16'b0000000000000100;
    assign weights1[60][431] = 16'b1111111111110101;
    assign weights1[60][432] = 16'b1111111111110001;
    assign weights1[60][433] = 16'b1111111111101000;
    assign weights1[60][434] = 16'b1111111111100000;
    assign weights1[60][435] = 16'b1111111111111000;
    assign weights1[60][436] = 16'b1111111111011101;
    assign weights1[60][437] = 16'b1111111111100110;
    assign weights1[60][438] = 16'b1111111111111011;
    assign weights1[60][439] = 16'b0000000000000001;
    assign weights1[60][440] = 16'b0000000000000101;
    assign weights1[60][441] = 16'b0000000000100011;
    assign weights1[60][442] = 16'b1111111111101001;
    assign weights1[60][443] = 16'b0000000000001001;
    assign weights1[60][444] = 16'b0000000000100110;
    assign weights1[60][445] = 16'b0000000000000000;
    assign weights1[60][446] = 16'b1111111111101100;
    assign weights1[60][447] = 16'b0000000000000110;
    assign weights1[60][448] = 16'b0000000000000101;
    assign weights1[60][449] = 16'b0000000000001100;
    assign weights1[60][450] = 16'b0000000000010100;
    assign weights1[60][451] = 16'b0000000000010001;
    assign weights1[60][452] = 16'b0000000000000110;
    assign weights1[60][453] = 16'b1111111111100011;
    assign weights1[60][454] = 16'b0000000000000011;
    assign weights1[60][455] = 16'b1111111111110100;
    assign weights1[60][456] = 16'b1111111111111010;
    assign weights1[60][457] = 16'b1111111111111000;
    assign weights1[60][458] = 16'b1111111111110001;
    assign weights1[60][459] = 16'b1111111111011000;
    assign weights1[60][460] = 16'b1111111111110101;
    assign weights1[60][461] = 16'b1111111111101001;
    assign weights1[60][462] = 16'b1111111111101111;
    assign weights1[60][463] = 16'b1111111111111001;
    assign weights1[60][464] = 16'b1111111111110110;
    assign weights1[60][465] = 16'b0000000000000111;
    assign weights1[60][466] = 16'b1111111111110111;
    assign weights1[60][467] = 16'b1111111111110111;
    assign weights1[60][468] = 16'b0000000000001011;
    assign weights1[60][469] = 16'b0000000000000010;
    assign weights1[60][470] = 16'b0000000000001101;
    assign weights1[60][471] = 16'b1111111111111011;
    assign weights1[60][472] = 16'b1111111111111000;
    assign weights1[60][473] = 16'b1111111111111000;
    assign weights1[60][474] = 16'b0000000000000010;
    assign weights1[60][475] = 16'b0000000000010001;
    assign weights1[60][476] = 16'b1111111111110110;
    assign weights1[60][477] = 16'b0000000000000011;
    assign weights1[60][478] = 16'b0000000000010111;
    assign weights1[60][479] = 16'b0000000000010111;
    assign weights1[60][480] = 16'b0000000000010010;
    assign weights1[60][481] = 16'b0000000000010111;
    assign weights1[60][482] = 16'b0000000000000100;
    assign weights1[60][483] = 16'b1111111111111100;
    assign weights1[60][484] = 16'b1111111111111100;
    assign weights1[60][485] = 16'b1111111111110001;
    assign weights1[60][486] = 16'b0000000000000011;
    assign weights1[60][487] = 16'b0000000000000011;
    assign weights1[60][488] = 16'b1111111111111100;
    assign weights1[60][489] = 16'b0000000000000001;
    assign weights1[60][490] = 16'b0000000000000000;
    assign weights1[60][491] = 16'b1111111111110101;
    assign weights1[60][492] = 16'b1111111111110101;
    assign weights1[60][493] = 16'b1111111111111111;
    assign weights1[60][494] = 16'b0000000000000010;
    assign weights1[60][495] = 16'b1111111111111010;
    assign weights1[60][496] = 16'b1111111111111111;
    assign weights1[60][497] = 16'b0000000000000001;
    assign weights1[60][498] = 16'b0000000000000101;
    assign weights1[60][499] = 16'b0000000000010010;
    assign weights1[60][500] = 16'b0000000000000100;
    assign weights1[60][501] = 16'b0000000000000000;
    assign weights1[60][502] = 16'b0000000000000011;
    assign weights1[60][503] = 16'b0000000000000011;
    assign weights1[60][504] = 16'b1111111111110110;
    assign weights1[60][505] = 16'b0000000000000101;
    assign weights1[60][506] = 16'b0000000000010000;
    assign weights1[60][507] = 16'b1111111111111100;
    assign weights1[60][508] = 16'b0000000000000011;
    assign weights1[60][509] = 16'b0000000000000000;
    assign weights1[60][510] = 16'b0000000000001010;
    assign weights1[60][511] = 16'b1111111111110111;
    assign weights1[60][512] = 16'b1111111111110111;
    assign weights1[60][513] = 16'b1111111111111001;
    assign weights1[60][514] = 16'b1111111111111100;
    assign weights1[60][515] = 16'b0000000000010011;
    assign weights1[60][516] = 16'b0000000000001110;
    assign weights1[60][517] = 16'b1111111111110010;
    assign weights1[60][518] = 16'b0000000000010100;
    assign weights1[60][519] = 16'b1111111111110000;
    assign weights1[60][520] = 16'b1111111111101101;
    assign weights1[60][521] = 16'b1111111111111011;
    assign weights1[60][522] = 16'b0000000000000000;
    assign weights1[60][523] = 16'b1111111111110111;
    assign weights1[60][524] = 16'b1111111111111101;
    assign weights1[60][525] = 16'b0000000000000100;
    assign weights1[60][526] = 16'b0000000000001000;
    assign weights1[60][527] = 16'b0000000000000101;
    assign weights1[60][528] = 16'b1111111111110101;
    assign weights1[60][529] = 16'b1111111111110100;
    assign weights1[60][530] = 16'b1111111111111100;
    assign weights1[60][531] = 16'b0000000000001010;
    assign weights1[60][532] = 16'b1111111111101110;
    assign weights1[60][533] = 16'b1111111111111000;
    assign weights1[60][534] = 16'b1111111111111100;
    assign weights1[60][535] = 16'b1111111111101100;
    assign weights1[60][536] = 16'b1111111111100100;
    assign weights1[60][537] = 16'b1111111111101110;
    assign weights1[60][538] = 16'b1111111111110000;
    assign weights1[60][539] = 16'b0000000000000111;
    assign weights1[60][540] = 16'b0000000000010011;
    assign weights1[60][541] = 16'b0000000000001001;
    assign weights1[60][542] = 16'b1111111111111101;
    assign weights1[60][543] = 16'b0000000000000000;
    assign weights1[60][544] = 16'b0000000000010001;
    assign weights1[60][545] = 16'b1111111111111000;
    assign weights1[60][546] = 16'b0000000000010001;
    assign weights1[60][547] = 16'b1111111111111010;
    assign weights1[60][548] = 16'b1111111111111011;
    assign weights1[60][549] = 16'b0000000000000100;
    assign weights1[60][550] = 16'b1111111111110110;
    assign weights1[60][551] = 16'b1111111111111111;
    assign weights1[60][552] = 16'b1111111111111111;
    assign weights1[60][553] = 16'b1111111111110111;
    assign weights1[60][554] = 16'b1111111111111100;
    assign weights1[60][555] = 16'b0000000000001001;
    assign weights1[60][556] = 16'b1111111111111101;
    assign weights1[60][557] = 16'b0000000000000110;
    assign weights1[60][558] = 16'b1111111111111000;
    assign weights1[60][559] = 16'b1111111111111111;
    assign weights1[60][560] = 16'b1111111111101111;
    assign weights1[60][561] = 16'b1111111111110001;
    assign weights1[60][562] = 16'b1111111111110100;
    assign weights1[60][563] = 16'b1111111111110101;
    assign weights1[60][564] = 16'b1111111111100100;
    assign weights1[60][565] = 16'b0000000000000100;
    assign weights1[60][566] = 16'b0000000000000111;
    assign weights1[60][567] = 16'b1111111111101001;
    assign weights1[60][568] = 16'b1111111111111101;
    assign weights1[60][569] = 16'b0000000000010001;
    assign weights1[60][570] = 16'b0000000000010001;
    assign weights1[60][571] = 16'b0000000000010001;
    assign weights1[60][572] = 16'b0000000000001010;
    assign weights1[60][573] = 16'b1111111111111000;
    assign weights1[60][574] = 16'b0000000000000010;
    assign weights1[60][575] = 16'b0000000000001010;
    assign weights1[60][576] = 16'b1111111111110001;
    assign weights1[60][577] = 16'b1111111111111100;
    assign weights1[60][578] = 16'b1111111111111100;
    assign weights1[60][579] = 16'b1111111111101110;
    assign weights1[60][580] = 16'b0000000000000101;
    assign weights1[60][581] = 16'b1111111111101111;
    assign weights1[60][582] = 16'b0000000000001001;
    assign weights1[60][583] = 16'b1111111111110011;
    assign weights1[60][584] = 16'b1111111111111101;
    assign weights1[60][585] = 16'b0000000000000010;
    assign weights1[60][586] = 16'b1111111111110010;
    assign weights1[60][587] = 16'b1111111111101101;
    assign weights1[60][588] = 16'b1111111111110011;
    assign weights1[60][589] = 16'b1111111111101011;
    assign weights1[60][590] = 16'b1111111111110100;
    assign weights1[60][591] = 16'b1111111111110111;
    assign weights1[60][592] = 16'b1111111111110100;
    assign weights1[60][593] = 16'b1111111111101111;
    assign weights1[60][594] = 16'b1111111111110011;
    assign weights1[60][595] = 16'b1111111111011001;
    assign weights1[60][596] = 16'b1111111111101100;
    assign weights1[60][597] = 16'b1111111111111011;
    assign weights1[60][598] = 16'b1111111111011110;
    assign weights1[60][599] = 16'b1111111111111001;
    assign weights1[60][600] = 16'b1111111111111011;
    assign weights1[60][601] = 16'b0000000000000110;
    assign weights1[60][602] = 16'b1111111111111110;
    assign weights1[60][603] = 16'b1111111111110111;
    assign weights1[60][604] = 16'b1111111111110111;
    assign weights1[60][605] = 16'b0000000000001011;
    assign weights1[60][606] = 16'b1111111111101101;
    assign weights1[60][607] = 16'b0000000000000000;
    assign weights1[60][608] = 16'b1111111111110111;
    assign weights1[60][609] = 16'b0000000000000111;
    assign weights1[60][610] = 16'b0000000000001000;
    assign weights1[60][611] = 16'b1111111111101110;
    assign weights1[60][612] = 16'b1111111111111000;
    assign weights1[60][613] = 16'b1111111111110010;
    assign weights1[60][614] = 16'b1111111111110110;
    assign weights1[60][615] = 16'b1111111111110101;
    assign weights1[60][616] = 16'b1111111111101110;
    assign weights1[60][617] = 16'b1111111111101110;
    assign weights1[60][618] = 16'b1111111111110110;
    assign weights1[60][619] = 16'b0000000000001111;
    assign weights1[60][620] = 16'b1111111111111000;
    assign weights1[60][621] = 16'b1111111111100011;
    assign weights1[60][622] = 16'b1111111111111100;
    assign weights1[60][623] = 16'b1111111111100110;
    assign weights1[60][624] = 16'b1111111111111111;
    assign weights1[60][625] = 16'b1111111111111010;
    assign weights1[60][626] = 16'b1111111111110110;
    assign weights1[60][627] = 16'b1111111111100010;
    assign weights1[60][628] = 16'b1111111111110101;
    assign weights1[60][629] = 16'b1111111111100110;
    assign weights1[60][630] = 16'b0000000000000010;
    assign weights1[60][631] = 16'b1111111111111100;
    assign weights1[60][632] = 16'b1111111111111010;
    assign weights1[60][633] = 16'b1111111111110100;
    assign weights1[60][634] = 16'b1111111111111011;
    assign weights1[60][635] = 16'b1111111111111101;
    assign weights1[60][636] = 16'b1111111111111110;
    assign weights1[60][637] = 16'b1111111111111110;
    assign weights1[60][638] = 16'b0000000000000000;
    assign weights1[60][639] = 16'b1111111111110010;
    assign weights1[60][640] = 16'b0000000000000011;
    assign weights1[60][641] = 16'b1111111111110000;
    assign weights1[60][642] = 16'b1111111111110011;
    assign weights1[60][643] = 16'b1111111111110101;
    assign weights1[60][644] = 16'b1111111111110110;
    assign weights1[60][645] = 16'b1111111111110101;
    assign weights1[60][646] = 16'b1111111111110111;
    assign weights1[60][647] = 16'b1111111111111000;
    assign weights1[60][648] = 16'b1111111111110111;
    assign weights1[60][649] = 16'b0000000000000000;
    assign weights1[60][650] = 16'b1111111111011101;
    assign weights1[60][651] = 16'b1111111111111001;
    assign weights1[60][652] = 16'b1111111111111111;
    assign weights1[60][653] = 16'b1111111111011001;
    assign weights1[60][654] = 16'b1111111111110001;
    assign weights1[60][655] = 16'b0000000000000001;
    assign weights1[60][656] = 16'b1111111111101101;
    assign weights1[60][657] = 16'b1111111111110010;
    assign weights1[60][658] = 16'b1111111111111111;
    assign weights1[60][659] = 16'b1111111111101110;
    assign weights1[60][660] = 16'b0000000000001000;
    assign weights1[60][661] = 16'b1111111111111100;
    assign weights1[60][662] = 16'b1111111111111010;
    assign weights1[60][663] = 16'b1111111111111100;
    assign weights1[60][664] = 16'b1111111111110101;
    assign weights1[60][665] = 16'b0000000000000110;
    assign weights1[60][666] = 16'b1111111111110110;
    assign weights1[60][667] = 16'b1111111111111000;
    assign weights1[60][668] = 16'b1111111111101101;
    assign weights1[60][669] = 16'b1111111111101100;
    assign weights1[60][670] = 16'b1111111111111000;
    assign weights1[60][671] = 16'b1111111111111000;
    assign weights1[60][672] = 16'b1111111111111010;
    assign weights1[60][673] = 16'b1111111111111010;
    assign weights1[60][674] = 16'b1111111111101110;
    assign weights1[60][675] = 16'b1111111111110101;
    assign weights1[60][676] = 16'b1111111111101000;
    assign weights1[60][677] = 16'b1111111111111100;
    assign weights1[60][678] = 16'b1111111111011000;
    assign weights1[60][679] = 16'b1111111111101101;
    assign weights1[60][680] = 16'b1111111111101111;
    assign weights1[60][681] = 16'b1111111111100110;
    assign weights1[60][682] = 16'b1111111111110111;
    assign weights1[60][683] = 16'b1111111111101100;
    assign weights1[60][684] = 16'b0000000000000011;
    assign weights1[60][685] = 16'b1111111111111110;
    assign weights1[60][686] = 16'b1111111111110111;
    assign weights1[60][687] = 16'b1111111111110001;
    assign weights1[60][688] = 16'b0000000000000000;
    assign weights1[60][689] = 16'b1111111111110000;
    assign weights1[60][690] = 16'b1111111111110011;
    assign weights1[60][691] = 16'b1111111111110101;
    assign weights1[60][692] = 16'b1111111111100010;
    assign weights1[60][693] = 16'b1111111111100111;
    assign weights1[60][694] = 16'b1111111111111001;
    assign weights1[60][695] = 16'b1111111111110111;
    assign weights1[60][696] = 16'b1111111111101011;
    assign weights1[60][697] = 16'b1111111111100011;
    assign weights1[60][698] = 16'b1111111111110001;
    assign weights1[60][699] = 16'b1111111111110111;
    assign weights1[60][700] = 16'b1111111111111101;
    assign weights1[60][701] = 16'b1111111111110101;
    assign weights1[60][702] = 16'b1111111111110100;
    assign weights1[60][703] = 16'b1111111111101011;
    assign weights1[60][704] = 16'b1111111111101011;
    assign weights1[60][705] = 16'b1111111111100001;
    assign weights1[60][706] = 16'b1111111111101111;
    assign weights1[60][707] = 16'b0000000000001000;
    assign weights1[60][708] = 16'b1111111111100111;
    assign weights1[60][709] = 16'b1111111111101110;
    assign weights1[60][710] = 16'b1111111111100101;
    assign weights1[60][711] = 16'b0000000000000010;
    assign weights1[60][712] = 16'b0000000000000110;
    assign weights1[60][713] = 16'b1111111111101110;
    assign weights1[60][714] = 16'b1111111111110100;
    assign weights1[60][715] = 16'b1111111111110010;
    assign weights1[60][716] = 16'b0000000000000110;
    assign weights1[60][717] = 16'b1111111111011001;
    assign weights1[60][718] = 16'b1111111111111100;
    assign weights1[60][719] = 16'b0000000000000011;
    assign weights1[60][720] = 16'b1111111111101010;
    assign weights1[60][721] = 16'b1111111111101011;
    assign weights1[60][722] = 16'b1111111111110110;
    assign weights1[60][723] = 16'b1111111111111100;
    assign weights1[60][724] = 16'b1111111111110110;
    assign weights1[60][725] = 16'b1111111111100111;
    assign weights1[60][726] = 16'b1111111111110101;
    assign weights1[60][727] = 16'b1111111111111110;
    assign weights1[60][728] = 16'b1111111111111110;
    assign weights1[60][729] = 16'b1111111111110101;
    assign weights1[60][730] = 16'b1111111111110011;
    assign weights1[60][731] = 16'b1111111111101101;
    assign weights1[60][732] = 16'b1111111111101010;
    assign weights1[60][733] = 16'b1111111111011100;
    assign weights1[60][734] = 16'b1111111111101111;
    assign weights1[60][735] = 16'b0000000000000001;
    assign weights1[60][736] = 16'b0000000000001000;
    assign weights1[60][737] = 16'b0000000000001010;
    assign weights1[60][738] = 16'b1111111111101111;
    assign weights1[60][739] = 16'b1111111111110110;
    assign weights1[60][740] = 16'b1111111111111110;
    assign weights1[60][741] = 16'b0000000000001011;
    assign weights1[60][742] = 16'b1111111111101101;
    assign weights1[60][743] = 16'b1111111111110100;
    assign weights1[60][744] = 16'b1111111111111111;
    assign weights1[60][745] = 16'b1111111111111011;
    assign weights1[60][746] = 16'b1111111111110101;
    assign weights1[60][747] = 16'b0000000000000000;
    assign weights1[60][748] = 16'b1111111111101110;
    assign weights1[60][749] = 16'b1111111111110101;
    assign weights1[60][750] = 16'b1111111111110100;
    assign weights1[60][751] = 16'b1111111111101010;
    assign weights1[60][752] = 16'b0000000000000000;
    assign weights1[60][753] = 16'b0000000000000000;
    assign weights1[60][754] = 16'b0000000000000101;
    assign weights1[60][755] = 16'b0000000000000001;
    assign weights1[60][756] = 16'b1111111111111101;
    assign weights1[60][757] = 16'b1111111111111000;
    assign weights1[60][758] = 16'b1111111111110000;
    assign weights1[60][759] = 16'b1111111111110100;
    assign weights1[60][760] = 16'b1111111111110110;
    assign weights1[60][761] = 16'b1111111111111101;
    assign weights1[60][762] = 16'b1111111111111011;
    assign weights1[60][763] = 16'b1111111111110101;
    assign weights1[60][764] = 16'b1111111111110000;
    assign weights1[60][765] = 16'b1111111111110001;
    assign weights1[60][766] = 16'b1111111111110101;
    assign weights1[60][767] = 16'b1111111111101010;
    assign weights1[60][768] = 16'b1111111111011100;
    assign weights1[60][769] = 16'b1111111111110001;
    assign weights1[60][770] = 16'b1111111111111001;
    assign weights1[60][771] = 16'b1111111111110001;
    assign weights1[60][772] = 16'b1111111111101011;
    assign weights1[60][773] = 16'b1111111111100011;
    assign weights1[60][774] = 16'b0000000000001101;
    assign weights1[60][775] = 16'b1111111111110010;
    assign weights1[60][776] = 16'b1111111111101000;
    assign weights1[60][777] = 16'b1111111111110000;
    assign weights1[60][778] = 16'b0000000000000001;
    assign weights1[60][779] = 16'b1111111111110111;
    assign weights1[60][780] = 16'b1111111111111101;
    assign weights1[60][781] = 16'b1111111111111101;
    assign weights1[60][782] = 16'b0000000000001010;
    assign weights1[60][783] = 16'b0000000000000101;
    assign weights1[61][0] = 16'b0000000000000000;
    assign weights1[61][1] = 16'b0000000000000000;
    assign weights1[61][2] = 16'b0000000000000000;
    assign weights1[61][3] = 16'b0000000000000001;
    assign weights1[61][4] = 16'b0000000000000010;
    assign weights1[61][5] = 16'b0000000000000010;
    assign weights1[61][6] = 16'b0000000000000000;
    assign weights1[61][7] = 16'b0000000000000001;
    assign weights1[61][8] = 16'b1111111111111110;
    assign weights1[61][9] = 16'b1111111111110010;
    assign weights1[61][10] = 16'b1111111111101101;
    assign weights1[61][11] = 16'b1111111111100101;
    assign weights1[61][12] = 16'b1111111111100100;
    assign weights1[61][13] = 16'b1111111111100001;
    assign weights1[61][14] = 16'b1111111111011101;
    assign weights1[61][15] = 16'b1111111111011110;
    assign weights1[61][16] = 16'b1111111111100010;
    assign weights1[61][17] = 16'b1111111111101001;
    assign weights1[61][18] = 16'b1111111111111000;
    assign weights1[61][19] = 16'b1111111111110010;
    assign weights1[61][20] = 16'b0000000000000100;
    assign weights1[61][21] = 16'b0000000000000110;
    assign weights1[61][22] = 16'b0000000000000000;
    assign weights1[61][23] = 16'b1111111111111010;
    assign weights1[61][24] = 16'b1111111111111110;
    assign weights1[61][25] = 16'b0000000000000100;
    assign weights1[61][26] = 16'b0000000000000111;
    assign weights1[61][27] = 16'b0000000000000101;
    assign weights1[61][28] = 16'b0000000000000000;
    assign weights1[61][29] = 16'b0000000000000000;
    assign weights1[61][30] = 16'b0000000000000001;
    assign weights1[61][31] = 16'b0000000000000010;
    assign weights1[61][32] = 16'b0000000000000100;
    assign weights1[61][33] = 16'b0000000000000011;
    assign weights1[61][34] = 16'b1111111111111100;
    assign weights1[61][35] = 16'b1111111111111010;
    assign weights1[61][36] = 16'b1111111111110101;
    assign weights1[61][37] = 16'b1111111111101010;
    assign weights1[61][38] = 16'b1111111111100011;
    assign weights1[61][39] = 16'b1111111111100110;
    assign weights1[61][40] = 16'b1111111111100101;
    assign weights1[61][41] = 16'b1111111111100011;
    assign weights1[61][42] = 16'b1111111111101010;
    assign weights1[61][43] = 16'b1111111111011011;
    assign weights1[61][44] = 16'b1111111111100011;
    assign weights1[61][45] = 16'b1111111111100010;
    assign weights1[61][46] = 16'b1111111111110010;
    assign weights1[61][47] = 16'b1111111111110101;
    assign weights1[61][48] = 16'b1111111111110101;
    assign weights1[61][49] = 16'b1111111111111110;
    assign weights1[61][50] = 16'b0000000000000101;
    assign weights1[61][51] = 16'b1111111111111111;
    assign weights1[61][52] = 16'b0000000000000000;
    assign weights1[61][53] = 16'b0000000000000111;
    assign weights1[61][54] = 16'b0000000000001000;
    assign weights1[61][55] = 16'b0000000000000110;
    assign weights1[61][56] = 16'b0000000000000000;
    assign weights1[61][57] = 16'b0000000000000100;
    assign weights1[61][58] = 16'b0000000000000100;
    assign weights1[61][59] = 16'b0000000000000011;
    assign weights1[61][60] = 16'b0000000000000010;
    assign weights1[61][61] = 16'b1111111111111111;
    assign weights1[61][62] = 16'b1111111111110111;
    assign weights1[61][63] = 16'b1111111111111010;
    assign weights1[61][64] = 16'b1111111111110000;
    assign weights1[61][65] = 16'b1111111111100100;
    assign weights1[61][66] = 16'b1111111111011010;
    assign weights1[61][67] = 16'b1111111111011010;
    assign weights1[61][68] = 16'b1111111111100011;
    assign weights1[61][69] = 16'b1111111111101000;
    assign weights1[61][70] = 16'b1111111111101000;
    assign weights1[61][71] = 16'b1111111111101111;
    assign weights1[61][72] = 16'b1111111111101111;
    assign weights1[61][73] = 16'b1111111111100101;
    assign weights1[61][74] = 16'b1111111111111101;
    assign weights1[61][75] = 16'b1111111111111101;
    assign weights1[61][76] = 16'b1111111111110101;
    assign weights1[61][77] = 16'b0000000000001001;
    assign weights1[61][78] = 16'b1111111111111101;
    assign weights1[61][79] = 16'b0000000000001100;
    assign weights1[61][80] = 16'b0000000000001011;
    assign weights1[61][81] = 16'b0000000000001100;
    assign weights1[61][82] = 16'b0000000000001101;
    assign weights1[61][83] = 16'b0000000000000110;
    assign weights1[61][84] = 16'b0000000000000000;
    assign weights1[61][85] = 16'b0000000000000010;
    assign weights1[61][86] = 16'b0000000000000011;
    assign weights1[61][87] = 16'b0000000000000000;
    assign weights1[61][88] = 16'b1111111111111111;
    assign weights1[61][89] = 16'b0000000000000000;
    assign weights1[61][90] = 16'b1111111111111101;
    assign weights1[61][91] = 16'b1111111111111100;
    assign weights1[61][92] = 16'b1111111111110000;
    assign weights1[61][93] = 16'b1111111111100100;
    assign weights1[61][94] = 16'b1111111111011001;
    assign weights1[61][95] = 16'b1111111111010111;
    assign weights1[61][96] = 16'b1111111111100111;
    assign weights1[61][97] = 16'b1111111111011110;
    assign weights1[61][98] = 16'b1111111111100001;
    assign weights1[61][99] = 16'b1111111111101011;
    assign weights1[61][100] = 16'b1111111111101101;
    assign weights1[61][101] = 16'b1111111111101001;
    assign weights1[61][102] = 16'b1111111111111101;
    assign weights1[61][103] = 16'b0000000000010001;
    assign weights1[61][104] = 16'b1111111111111101;
    assign weights1[61][105] = 16'b1111111111111101;
    assign weights1[61][106] = 16'b0000000000000110;
    assign weights1[61][107] = 16'b0000000000001101;
    assign weights1[61][108] = 16'b0000000000011000;
    assign weights1[61][109] = 16'b0000000000010100;
    assign weights1[61][110] = 16'b0000000000011011;
    assign weights1[61][111] = 16'b0000000000001100;
    assign weights1[61][112] = 16'b0000000000000001;
    assign weights1[61][113] = 16'b0000000000000001;
    assign weights1[61][114] = 16'b0000000000000010;
    assign weights1[61][115] = 16'b1111111111111011;
    assign weights1[61][116] = 16'b1111111111111000;
    assign weights1[61][117] = 16'b1111111111111010;
    assign weights1[61][118] = 16'b0000000000000000;
    assign weights1[61][119] = 16'b1111111111110010;
    assign weights1[61][120] = 16'b1111111111100000;
    assign weights1[61][121] = 16'b1111111111101001;
    assign weights1[61][122] = 16'b1111111111001000;
    assign weights1[61][123] = 16'b1111111111001001;
    assign weights1[61][124] = 16'b1111111110111110;
    assign weights1[61][125] = 16'b1111111111010100;
    assign weights1[61][126] = 16'b1111111111010110;
    assign weights1[61][127] = 16'b1111111111110010;
    assign weights1[61][128] = 16'b1111111111011101;
    assign weights1[61][129] = 16'b1111111111111100;
    assign weights1[61][130] = 16'b0000000000000000;
    assign weights1[61][131] = 16'b1111111111111101;
    assign weights1[61][132] = 16'b0000000000000111;
    assign weights1[61][133] = 16'b0000000000100011;
    assign weights1[61][134] = 16'b0000000000110111;
    assign weights1[61][135] = 16'b0000000000101101;
    assign weights1[61][136] = 16'b0000000000011011;
    assign weights1[61][137] = 16'b0000000000001011;
    assign weights1[61][138] = 16'b0000000000010010;
    assign weights1[61][139] = 16'b0000000000001010;
    assign weights1[61][140] = 16'b0000000000000001;
    assign weights1[61][141] = 16'b0000000000000001;
    assign weights1[61][142] = 16'b1111111111111100;
    assign weights1[61][143] = 16'b1111111111110101;
    assign weights1[61][144] = 16'b1111111111110011;
    assign weights1[61][145] = 16'b1111111111111100;
    assign weights1[61][146] = 16'b1111111111111011;
    assign weights1[61][147] = 16'b1111111111001011;
    assign weights1[61][148] = 16'b1111111111001010;
    assign weights1[61][149] = 16'b1111111110111111;
    assign weights1[61][150] = 16'b1111111110111110;
    assign weights1[61][151] = 16'b1111111111011101;
    assign weights1[61][152] = 16'b1111111111111111;
    assign weights1[61][153] = 16'b0000000000001011;
    assign weights1[61][154] = 16'b1111111111110111;
    assign weights1[61][155] = 16'b1111111111110000;
    assign weights1[61][156] = 16'b1111111111101111;
    assign weights1[61][157] = 16'b0000000000000111;
    assign weights1[61][158] = 16'b0000000000100000;
    assign weights1[61][159] = 16'b0000000000000011;
    assign weights1[61][160] = 16'b0000000000100000;
    assign weights1[61][161] = 16'b0000000000100100;
    assign weights1[61][162] = 16'b0000000000010101;
    assign weights1[61][163] = 16'b0000000000011110;
    assign weights1[61][164] = 16'b0000000000101011;
    assign weights1[61][165] = 16'b0000000000100000;
    assign weights1[61][166] = 16'b0000000000011110;
    assign weights1[61][167] = 16'b0000000000011001;
    assign weights1[61][168] = 16'b0000000000000000;
    assign weights1[61][169] = 16'b1111111111111111;
    assign weights1[61][170] = 16'b1111111111111010;
    assign weights1[61][171] = 16'b1111111111111001;
    assign weights1[61][172] = 16'b1111111111110111;
    assign weights1[61][173] = 16'b1111111111111101;
    assign weights1[61][174] = 16'b1111111111111100;
    assign weights1[61][175] = 16'b1111111111011100;
    assign weights1[61][176] = 16'b1111111110111001;
    assign weights1[61][177] = 16'b1111111110111001;
    assign weights1[61][178] = 16'b1111111111010101;
    assign weights1[61][179] = 16'b1111111110110101;
    assign weights1[61][180] = 16'b1111111111110111;
    assign weights1[61][181] = 16'b0000000000101100;
    assign weights1[61][182] = 16'b0000000000010111;
    assign weights1[61][183] = 16'b0000000000010010;
    assign weights1[61][184] = 16'b1111111111110111;
    assign weights1[61][185] = 16'b0000000000011100;
    assign weights1[61][186] = 16'b0000000000001010;
    assign weights1[61][187] = 16'b0000000000100010;
    assign weights1[61][188] = 16'b0000000000100011;
    assign weights1[61][189] = 16'b0000000000011101;
    assign weights1[61][190] = 16'b0000000000011011;
    assign weights1[61][191] = 16'b1111111111111011;
    assign weights1[61][192] = 16'b0000000000101000;
    assign weights1[61][193] = 16'b0000000000100011;
    assign weights1[61][194] = 16'b0000000000110111;
    assign weights1[61][195] = 16'b0000000000101010;
    assign weights1[61][196] = 16'b1111111111111111;
    assign weights1[61][197] = 16'b1111111111111110;
    assign weights1[61][198] = 16'b1111111111111001;
    assign weights1[61][199] = 16'b1111111111111011;
    assign weights1[61][200] = 16'b1111111111110111;
    assign weights1[61][201] = 16'b1111111111111101;
    assign weights1[61][202] = 16'b1111111111101000;
    assign weights1[61][203] = 16'b1111111111001101;
    assign weights1[61][204] = 16'b1111111111001111;
    assign weights1[61][205] = 16'b1111111110111110;
    assign weights1[61][206] = 16'b1111111111101000;
    assign weights1[61][207] = 16'b0000000000101100;
    assign weights1[61][208] = 16'b0000000000100011;
    assign weights1[61][209] = 16'b0000000000110100;
    assign weights1[61][210] = 16'b0000000000001011;
    assign weights1[61][211] = 16'b0000000000100000;
    assign weights1[61][212] = 16'b0000000000011010;
    assign weights1[61][213] = 16'b0000000000011011;
    assign weights1[61][214] = 16'b0000000000011001;
    assign weights1[61][215] = 16'b0000000000010001;
    assign weights1[61][216] = 16'b0000000000010010;
    assign weights1[61][217] = 16'b0000000000001100;
    assign weights1[61][218] = 16'b0000000000011111;
    assign weights1[61][219] = 16'b0000000000010110;
    assign weights1[61][220] = 16'b0000000000100111;
    assign weights1[61][221] = 16'b0000000000100001;
    assign weights1[61][222] = 16'b0000000000100100;
    assign weights1[61][223] = 16'b0000000000110010;
    assign weights1[61][224] = 16'b1111111111111110;
    assign weights1[61][225] = 16'b1111111111111100;
    assign weights1[61][226] = 16'b0000000000000000;
    assign weights1[61][227] = 16'b1111111111110100;
    assign weights1[61][228] = 16'b1111111111101100;
    assign weights1[61][229] = 16'b1111111111101011;
    assign weights1[61][230] = 16'b1111111111010011;
    assign weights1[61][231] = 16'b1111111110101111;
    assign weights1[61][232] = 16'b1111111110011011;
    assign weights1[61][233] = 16'b1111111111010110;
    assign weights1[61][234] = 16'b1111111111101101;
    assign weights1[61][235] = 16'b0000000000101010;
    assign weights1[61][236] = 16'b0000000000110111;
    assign weights1[61][237] = 16'b0000000000011111;
    assign weights1[61][238] = 16'b0000000000110011;
    assign weights1[61][239] = 16'b0000000000001111;
    assign weights1[61][240] = 16'b0000000000101111;
    assign weights1[61][241] = 16'b0000000000100000;
    assign weights1[61][242] = 16'b0000000000001011;
    assign weights1[61][243] = 16'b0000000000011000;
    assign weights1[61][244] = 16'b0000000000011011;
    assign weights1[61][245] = 16'b0000000000001111;
    assign weights1[61][246] = 16'b0000000000001101;
    assign weights1[61][247] = 16'b0000000001000110;
    assign weights1[61][248] = 16'b0000000000101010;
    assign weights1[61][249] = 16'b0000000000100110;
    assign weights1[61][250] = 16'b0000000000010100;
    assign weights1[61][251] = 16'b0000000000100111;
    assign weights1[61][252] = 16'b1111111111111100;
    assign weights1[61][253] = 16'b1111111111111010;
    assign weights1[61][254] = 16'b1111111111111010;
    assign weights1[61][255] = 16'b1111111111110011;
    assign weights1[61][256] = 16'b1111111111101010;
    assign weights1[61][257] = 16'b1111111111100011;
    assign weights1[61][258] = 16'b1111111111000001;
    assign weights1[61][259] = 16'b1111111110110001;
    assign weights1[61][260] = 16'b1111111111000100;
    assign weights1[61][261] = 16'b1111111111101101;
    assign weights1[61][262] = 16'b0000000000000010;
    assign weights1[61][263] = 16'b0000000000011110;
    assign weights1[61][264] = 16'b0000000000101001;
    assign weights1[61][265] = 16'b0000000001001111;
    assign weights1[61][266] = 16'b0000000000110110;
    assign weights1[61][267] = 16'b0000000000001011;
    assign weights1[61][268] = 16'b1111111111110100;
    assign weights1[61][269] = 16'b0000000000101001;
    assign weights1[61][270] = 16'b0000000000110011;
    assign weights1[61][271] = 16'b0000000000010000;
    assign weights1[61][272] = 16'b0000000000010100;
    assign weights1[61][273] = 16'b0000000000011100;
    assign weights1[61][274] = 16'b1111111111111100;
    assign weights1[61][275] = 16'b0000000000001011;
    assign weights1[61][276] = 16'b0000000000010111;
    assign weights1[61][277] = 16'b0000000000011100;
    assign weights1[61][278] = 16'b0000000000000111;
    assign weights1[61][279] = 16'b0000000000101110;
    assign weights1[61][280] = 16'b1111111111111010;
    assign weights1[61][281] = 16'b1111111111111011;
    assign weights1[61][282] = 16'b1111111111111100;
    assign weights1[61][283] = 16'b1111111111110000;
    assign weights1[61][284] = 16'b1111111111101100;
    assign weights1[61][285] = 16'b1111111111010101;
    assign weights1[61][286] = 16'b1111111110111010;
    assign weights1[61][287] = 16'b1111111111001001;
    assign weights1[61][288] = 16'b1111111111100110;
    assign weights1[61][289] = 16'b0000000000000101;
    assign weights1[61][290] = 16'b0000000000001010;
    assign weights1[61][291] = 16'b0000000000111011;
    assign weights1[61][292] = 16'b0000000000110101;
    assign weights1[61][293] = 16'b0000000000111011;
    assign weights1[61][294] = 16'b0000000000001010;
    assign weights1[61][295] = 16'b1111111111101010;
    assign weights1[61][296] = 16'b1111111111011110;
    assign weights1[61][297] = 16'b1111111111101110;
    assign weights1[61][298] = 16'b1111111111110001;
    assign weights1[61][299] = 16'b1111111111010001;
    assign weights1[61][300] = 16'b1111111111110101;
    assign weights1[61][301] = 16'b1111111111011111;
    assign weights1[61][302] = 16'b1111111111100111;
    assign weights1[61][303] = 16'b1111111111100111;
    assign weights1[61][304] = 16'b1111111111101011;
    assign weights1[61][305] = 16'b0000000000000011;
    assign weights1[61][306] = 16'b0000000000001101;
    assign weights1[61][307] = 16'b0000000000000110;
    assign weights1[61][308] = 16'b1111111111111010;
    assign weights1[61][309] = 16'b1111111111111100;
    assign weights1[61][310] = 16'b1111111111111001;
    assign weights1[61][311] = 16'b1111111111101110;
    assign weights1[61][312] = 16'b1111111111100101;
    assign weights1[61][313] = 16'b1111111111010110;
    assign weights1[61][314] = 16'b1111111110111111;
    assign weights1[61][315] = 16'b1111111111001011;
    assign weights1[61][316] = 16'b1111111111111000;
    assign weights1[61][317] = 16'b1111111111111110;
    assign weights1[61][318] = 16'b0000000000010010;
    assign weights1[61][319] = 16'b0000000000000110;
    assign weights1[61][320] = 16'b0000000001001000;
    assign weights1[61][321] = 16'b0000000000111110;
    assign weights1[61][322] = 16'b1111111111101110;
    assign weights1[61][323] = 16'b1111111110011111;
    assign weights1[61][324] = 16'b1111111110100000;
    assign weights1[61][325] = 16'b1111111111000000;
    assign weights1[61][326] = 16'b1111111111110101;
    assign weights1[61][327] = 16'b1111111111110100;
    assign weights1[61][328] = 16'b1111111111010110;
    assign weights1[61][329] = 16'b1111111111100010;
    assign weights1[61][330] = 16'b1111111111101001;
    assign weights1[61][331] = 16'b1111111111100100;
    assign weights1[61][332] = 16'b1111111111101010;
    assign weights1[61][333] = 16'b0000000000000110;
    assign weights1[61][334] = 16'b0000000000000001;
    assign weights1[61][335] = 16'b1111111111111101;
    assign weights1[61][336] = 16'b1111111111111011;
    assign weights1[61][337] = 16'b1111111111111111;
    assign weights1[61][338] = 16'b1111111111111101;
    assign weights1[61][339] = 16'b1111111111100110;
    assign weights1[61][340] = 16'b1111111111010001;
    assign weights1[61][341] = 16'b1111111111000111;
    assign weights1[61][342] = 16'b1111111111010110;
    assign weights1[61][343] = 16'b1111111111010011;
    assign weights1[61][344] = 16'b0000000000010000;
    assign weights1[61][345] = 16'b1111111111111001;
    assign weights1[61][346] = 16'b0000000000100101;
    assign weights1[61][347] = 16'b0000000000100111;
    assign weights1[61][348] = 16'b0000000000100011;
    assign weights1[61][349] = 16'b0000000001000011;
    assign weights1[61][350] = 16'b1111111111101001;
    assign weights1[61][351] = 16'b1111111110010011;
    assign weights1[61][352] = 16'b1111111110101010;
    assign weights1[61][353] = 16'b1111111111100111;
    assign weights1[61][354] = 16'b1111111111110100;
    assign weights1[61][355] = 16'b1111111111101010;
    assign weights1[61][356] = 16'b1111111111101100;
    assign weights1[61][357] = 16'b1111111111011101;
    assign weights1[61][358] = 16'b1111111111011111;
    assign weights1[61][359] = 16'b1111111111100010;
    assign weights1[61][360] = 16'b1111111111111101;
    assign weights1[61][361] = 16'b1111111111110110;
    assign weights1[61][362] = 16'b1111111111110100;
    assign weights1[61][363] = 16'b0000000000000100;
    assign weights1[61][364] = 16'b1111111111111010;
    assign weights1[61][365] = 16'b1111111111110111;
    assign weights1[61][366] = 16'b1111111111110111;
    assign weights1[61][367] = 16'b1111111111100000;
    assign weights1[61][368] = 16'b1111111111001101;
    assign weights1[61][369] = 16'b1111111111101001;
    assign weights1[61][370] = 16'b0000000000000001;
    assign weights1[61][371] = 16'b1111111111101110;
    assign weights1[61][372] = 16'b0000000000001011;
    assign weights1[61][373] = 16'b1111111111111111;
    assign weights1[61][374] = 16'b0000000000011111;
    assign weights1[61][375] = 16'b0000000000010001;
    assign weights1[61][376] = 16'b0000000000111010;
    assign weights1[61][377] = 16'b0000000000011111;
    assign weights1[61][378] = 16'b1111111110111110;
    assign weights1[61][379] = 16'b1111111110000101;
    assign weights1[61][380] = 16'b1111111111000110;
    assign weights1[61][381] = 16'b1111111111011001;
    assign weights1[61][382] = 16'b1111111111011100;
    assign weights1[61][383] = 16'b1111111111101011;
    assign weights1[61][384] = 16'b1111111111101111;
    assign weights1[61][385] = 16'b1111111111100010;
    assign weights1[61][386] = 16'b1111111111101011;
    assign weights1[61][387] = 16'b1111111111110000;
    assign weights1[61][388] = 16'b0000000000000100;
    assign weights1[61][389] = 16'b1111111111110100;
    assign weights1[61][390] = 16'b0000000000010011;
    assign weights1[61][391] = 16'b0000000000011000;
    assign weights1[61][392] = 16'b1111111111110111;
    assign weights1[61][393] = 16'b1111111111110010;
    assign weights1[61][394] = 16'b1111111111110011;
    assign weights1[61][395] = 16'b1111111111101111;
    assign weights1[61][396] = 16'b1111111111001100;
    assign weights1[61][397] = 16'b1111111111101111;
    assign weights1[61][398] = 16'b1111111111011110;
    assign weights1[61][399] = 16'b1111111111111111;
    assign weights1[61][400] = 16'b0000000000001000;
    assign weights1[61][401] = 16'b0000000000100110;
    assign weights1[61][402] = 16'b0000000000101011;
    assign weights1[61][403] = 16'b0000000000000010;
    assign weights1[61][404] = 16'b0000000000001110;
    assign weights1[61][405] = 16'b1111111111101011;
    assign weights1[61][406] = 16'b1111111110100001;
    assign weights1[61][407] = 16'b1111111110011110;
    assign weights1[61][408] = 16'b1111111111000011;
    assign weights1[61][409] = 16'b1111111111101001;
    assign weights1[61][410] = 16'b1111111111110011;
    assign weights1[61][411] = 16'b1111111111100111;
    assign weights1[61][412] = 16'b1111111111010101;
    assign weights1[61][413] = 16'b1111111111110010;
    assign weights1[61][414] = 16'b0000000000000010;
    assign weights1[61][415] = 16'b1111111111100011;
    assign weights1[61][416] = 16'b1111111111111101;
    assign weights1[61][417] = 16'b0000000000010001;
    assign weights1[61][418] = 16'b0000000000011100;
    assign weights1[61][419] = 16'b0000000000010011;
    assign weights1[61][420] = 16'b1111111111110001;
    assign weights1[61][421] = 16'b1111111111101111;
    assign weights1[61][422] = 16'b1111111111101111;
    assign weights1[61][423] = 16'b1111111111101000;
    assign weights1[61][424] = 16'b1111111111010111;
    assign weights1[61][425] = 16'b0000000000000011;
    assign weights1[61][426] = 16'b1111111111101001;
    assign weights1[61][427] = 16'b0000000000001010;
    assign weights1[61][428] = 16'b1111111111110100;
    assign weights1[61][429] = 16'b0000000000010100;
    assign weights1[61][430] = 16'b0000000000001101;
    assign weights1[61][431] = 16'b0000000000000000;
    assign weights1[61][432] = 16'b0000000000000010;
    assign weights1[61][433] = 16'b1111111111001111;
    assign weights1[61][434] = 16'b1111111110001001;
    assign weights1[61][435] = 16'b1111111110110111;
    assign weights1[61][436] = 16'b1111111111010100;
    assign weights1[61][437] = 16'b1111111111011101;
    assign weights1[61][438] = 16'b1111111111101010;
    assign weights1[61][439] = 16'b1111111111010111;
    assign weights1[61][440] = 16'b0000000000000000;
    assign weights1[61][441] = 16'b1111111111110111;
    assign weights1[61][442] = 16'b1111111111100011;
    assign weights1[61][443] = 16'b0000000000000000;
    assign weights1[61][444] = 16'b1111111111101001;
    assign weights1[61][445] = 16'b0000000000010000;
    assign weights1[61][446] = 16'b1111111111111010;
    assign weights1[61][447] = 16'b0000000000001011;
    assign weights1[61][448] = 16'b1111111111110100;
    assign weights1[61][449] = 16'b1111111111111010;
    assign weights1[61][450] = 16'b1111111111101011;
    assign weights1[61][451] = 16'b1111111111100001;
    assign weights1[61][452] = 16'b1111111111011111;
    assign weights1[61][453] = 16'b1111111111111101;
    assign weights1[61][454] = 16'b1111111111101111;
    assign weights1[61][455] = 16'b1111111111100101;
    assign weights1[61][456] = 16'b1111111111111101;
    assign weights1[61][457] = 16'b0000000000000010;
    assign weights1[61][458] = 16'b0000000000001000;
    assign weights1[61][459] = 16'b0000000000001110;
    assign weights1[61][460] = 16'b1111111111100000;
    assign weights1[61][461] = 16'b1111111110110010;
    assign weights1[61][462] = 16'b1111111110110000;
    assign weights1[61][463] = 16'b1111111111000011;
    assign weights1[61][464] = 16'b1111111111001111;
    assign weights1[61][465] = 16'b1111111111100101;
    assign weights1[61][466] = 16'b1111111111111011;
    assign weights1[61][467] = 16'b1111111111111011;
    assign weights1[61][468] = 16'b1111111111101110;
    assign weights1[61][469] = 16'b0000000000001101;
    assign weights1[61][470] = 16'b0000000000001000;
    assign weights1[61][471] = 16'b1111111111111110;
    assign weights1[61][472] = 16'b0000000000000110;
    assign weights1[61][473] = 16'b0000000000000001;
    assign weights1[61][474] = 16'b0000000000000111;
    assign weights1[61][475] = 16'b0000000000000000;
    assign weights1[61][476] = 16'b1111111111111010;
    assign weights1[61][477] = 16'b1111111111110111;
    assign weights1[61][478] = 16'b1111111111101111;
    assign weights1[61][479] = 16'b1111111111100011;
    assign weights1[61][480] = 16'b1111111111011011;
    assign weights1[61][481] = 16'b1111111111111110;
    assign weights1[61][482] = 16'b1111111111111100;
    assign weights1[61][483] = 16'b1111111111110001;
    assign weights1[61][484] = 16'b1111111111110010;
    assign weights1[61][485] = 16'b1111111111001111;
    assign weights1[61][486] = 16'b1111111111110011;
    assign weights1[61][487] = 16'b0000000000000010;
    assign weights1[61][488] = 16'b1111111111010100;
    assign weights1[61][489] = 16'b1111111111001101;
    assign weights1[61][490] = 16'b1111111110111000;
    assign weights1[61][491] = 16'b1111111111011111;
    assign weights1[61][492] = 16'b1111111111101111;
    assign weights1[61][493] = 16'b1111111111111001;
    assign weights1[61][494] = 16'b0000000000010110;
    assign weights1[61][495] = 16'b1111111111111111;
    assign weights1[61][496] = 16'b0000000000001000;
    assign weights1[61][497] = 16'b1111111111111010;
    assign weights1[61][498] = 16'b0000000000000011;
    assign weights1[61][499] = 16'b0000000000000010;
    assign weights1[61][500] = 16'b1111111111111001;
    assign weights1[61][501] = 16'b0000000000000011;
    assign weights1[61][502] = 16'b0000000000001010;
    assign weights1[61][503] = 16'b0000000000001010;
    assign weights1[61][504] = 16'b1111111111111111;
    assign weights1[61][505] = 16'b0000000000000000;
    assign weights1[61][506] = 16'b1111111111111100;
    assign weights1[61][507] = 16'b1111111111110010;
    assign weights1[61][508] = 16'b1111111111101100;
    assign weights1[61][509] = 16'b1111111111111000;
    assign weights1[61][510] = 16'b0000000000010111;
    assign weights1[61][511] = 16'b1111111111111101;
    assign weights1[61][512] = 16'b1111111111111000;
    assign weights1[61][513] = 16'b1111111111111100;
    assign weights1[61][514] = 16'b1111111111110000;
    assign weights1[61][515] = 16'b1111111111110101;
    assign weights1[61][516] = 16'b1111111111001011;
    assign weights1[61][517] = 16'b1111111111101110;
    assign weights1[61][518] = 16'b1111111111001010;
    assign weights1[61][519] = 16'b1111111111110001;
    assign weights1[61][520] = 16'b0000000000001011;
    assign weights1[61][521] = 16'b1111111111111111;
    assign weights1[61][522] = 16'b1111111111101010;
    assign weights1[61][523] = 16'b1111111111111010;
    assign weights1[61][524] = 16'b0000000000000001;
    assign weights1[61][525] = 16'b1111111111100011;
    assign weights1[61][526] = 16'b0000000000000110;
    assign weights1[61][527] = 16'b1111111111110111;
    assign weights1[61][528] = 16'b1111111111110011;
    assign weights1[61][529] = 16'b0000000000001111;
    assign weights1[61][530] = 16'b1111111111111101;
    assign weights1[61][531] = 16'b0000000000000101;
    assign weights1[61][532] = 16'b0000000000000011;
    assign weights1[61][533] = 16'b0000000000000111;
    assign weights1[61][534] = 16'b0000000000000110;
    assign weights1[61][535] = 16'b1111111111100110;
    assign weights1[61][536] = 16'b1111111111111010;
    assign weights1[61][537] = 16'b1111111111111111;
    assign weights1[61][538] = 16'b0000000000010111;
    assign weights1[61][539] = 16'b0000000000100111;
    assign weights1[61][540] = 16'b1111111111101111;
    assign weights1[61][541] = 16'b0000000000000101;
    assign weights1[61][542] = 16'b1111111111111111;
    assign weights1[61][543] = 16'b0000000000001100;
    assign weights1[61][544] = 16'b1111111111111000;
    assign weights1[61][545] = 16'b1111111111111100;
    assign weights1[61][546] = 16'b0000000000010100;
    assign weights1[61][547] = 16'b1111111111110111;
    assign weights1[61][548] = 16'b1111111111110101;
    assign weights1[61][549] = 16'b1111111111110011;
    assign weights1[61][550] = 16'b0000000000001110;
    assign weights1[61][551] = 16'b1111111111110111;
    assign weights1[61][552] = 16'b0000000000010010;
    assign weights1[61][553] = 16'b1111111111110100;
    assign weights1[61][554] = 16'b0000000000000001;
    assign weights1[61][555] = 16'b0000000000000010;
    assign weights1[61][556] = 16'b0000000000000010;
    assign weights1[61][557] = 16'b1111111111111111;
    assign weights1[61][558] = 16'b1111111111110110;
    assign weights1[61][559] = 16'b1111111111110111;
    assign weights1[61][560] = 16'b0000000000000000;
    assign weights1[61][561] = 16'b0000000000001110;
    assign weights1[61][562] = 16'b0000000000000010;
    assign weights1[61][563] = 16'b1111111111011011;
    assign weights1[61][564] = 16'b0000000000000110;
    assign weights1[61][565] = 16'b0000000000000001;
    assign weights1[61][566] = 16'b0000000000100000;
    assign weights1[61][567] = 16'b1111111111110101;
    assign weights1[61][568] = 16'b0000000000010101;
    assign weights1[61][569] = 16'b0000000000001010;
    assign weights1[61][570] = 16'b0000000000010111;
    assign weights1[61][571] = 16'b0000000000000110;
    assign weights1[61][572] = 16'b0000000000000010;
    assign weights1[61][573] = 16'b1111111111111110;
    assign weights1[61][574] = 16'b1111111111011101;
    assign weights1[61][575] = 16'b0000000000000101;
    assign weights1[61][576] = 16'b0000000000000001;
    assign weights1[61][577] = 16'b1111111111110010;
    assign weights1[61][578] = 16'b0000000000001101;
    assign weights1[61][579] = 16'b0000000000001001;
    assign weights1[61][580] = 16'b1111111111111011;
    assign weights1[61][581] = 16'b0000000000000100;
    assign weights1[61][582] = 16'b1111111111110100;
    assign weights1[61][583] = 16'b1111111111101011;
    assign weights1[61][584] = 16'b1111111111110110;
    assign weights1[61][585] = 16'b1111111111110011;
    assign weights1[61][586] = 16'b1111111111110001;
    assign weights1[61][587] = 16'b1111111111101111;
    assign weights1[61][588] = 16'b1111111111111101;
    assign weights1[61][589] = 16'b0000000000000010;
    assign weights1[61][590] = 16'b1111111111111101;
    assign weights1[61][591] = 16'b1111111111101011;
    assign weights1[61][592] = 16'b1111111111110110;
    assign weights1[61][593] = 16'b1111111111101000;
    assign weights1[61][594] = 16'b1111111111100111;
    assign weights1[61][595] = 16'b1111111111111101;
    assign weights1[61][596] = 16'b0000000000010100;
    assign weights1[61][597] = 16'b0000000000000100;
    assign weights1[61][598] = 16'b1111111111111100;
    assign weights1[61][599] = 16'b0000000000011000;
    assign weights1[61][600] = 16'b0000000000000111;
    assign weights1[61][601] = 16'b0000000000000110;
    assign weights1[61][602] = 16'b1111111111111010;
    assign weights1[61][603] = 16'b1111111111111000;
    assign weights1[61][604] = 16'b1111111111111100;
    assign weights1[61][605] = 16'b1111111111110000;
    assign weights1[61][606] = 16'b0000000000010001;
    assign weights1[61][607] = 16'b0000000000000001;
    assign weights1[61][608] = 16'b1111111111110011;
    assign weights1[61][609] = 16'b1111111111111100;
    assign weights1[61][610] = 16'b1111111111111101;
    assign weights1[61][611] = 16'b1111111111100100;
    assign weights1[61][612] = 16'b1111111111110000;
    assign weights1[61][613] = 16'b1111111111101111;
    assign weights1[61][614] = 16'b1111111111110110;
    assign weights1[61][615] = 16'b1111111111101101;
    assign weights1[61][616] = 16'b1111111111111101;
    assign weights1[61][617] = 16'b1111111111111101;
    assign weights1[61][618] = 16'b1111111111110100;
    assign weights1[61][619] = 16'b1111111111100110;
    assign weights1[61][620] = 16'b1111111111101000;
    assign weights1[61][621] = 16'b1111111111011100;
    assign weights1[61][622] = 16'b1111111111110111;
    assign weights1[61][623] = 16'b1111111111101111;
    assign weights1[61][624] = 16'b0000000000001000;
    assign weights1[61][625] = 16'b0000000000000001;
    assign weights1[61][626] = 16'b0000000000001000;
    assign weights1[61][627] = 16'b0000000000001011;
    assign weights1[61][628] = 16'b0000000000001110;
    assign weights1[61][629] = 16'b1111111111101100;
    assign weights1[61][630] = 16'b0000000000000111;
    assign weights1[61][631] = 16'b0000000000000111;
    assign weights1[61][632] = 16'b0000000000001010;
    assign weights1[61][633] = 16'b0000000000001101;
    assign weights1[61][634] = 16'b0000000000001010;
    assign weights1[61][635] = 16'b1111111111111001;
    assign weights1[61][636] = 16'b1111111111111100;
    assign weights1[61][637] = 16'b1111111111110010;
    assign weights1[61][638] = 16'b1111111111110011;
    assign weights1[61][639] = 16'b1111111111011111;
    assign weights1[61][640] = 16'b1111111111101100;
    assign weights1[61][641] = 16'b1111111111101100;
    assign weights1[61][642] = 16'b1111111111110000;
    assign weights1[61][643] = 16'b1111111111110010;
    assign weights1[61][644] = 16'b0000000000000000;
    assign weights1[61][645] = 16'b1111111111111101;
    assign weights1[61][646] = 16'b1111111111110110;
    assign weights1[61][647] = 16'b1111111111100110;
    assign weights1[61][648] = 16'b1111111111110000;
    assign weights1[61][649] = 16'b1111111111110101;
    assign weights1[61][650] = 16'b0000000000001101;
    assign weights1[61][651] = 16'b1111111111110100;
    assign weights1[61][652] = 16'b1111111111011100;
    assign weights1[61][653] = 16'b1111111111100100;
    assign weights1[61][654] = 16'b0000000000100001;
    assign weights1[61][655] = 16'b0000000000001101;
    assign weights1[61][656] = 16'b1111111111111101;
    assign weights1[61][657] = 16'b0000000000001110;
    assign weights1[61][658] = 16'b0000000000011001;
    assign weights1[61][659] = 16'b1111111111110010;
    assign weights1[61][660] = 16'b0000000000010010;
    assign weights1[61][661] = 16'b1111111111110001;
    assign weights1[61][662] = 16'b1111111111011111;
    assign weights1[61][663] = 16'b1111111111110101;
    assign weights1[61][664] = 16'b1111111111111111;
    assign weights1[61][665] = 16'b1111111111111001;
    assign weights1[61][666] = 16'b1111111111101010;
    assign weights1[61][667] = 16'b1111111111110001;
    assign weights1[61][668] = 16'b1111111111101001;
    assign weights1[61][669] = 16'b1111111111101111;
    assign weights1[61][670] = 16'b1111111111101101;
    assign weights1[61][671] = 16'b1111111111110001;
    assign weights1[61][672] = 16'b1111111111111110;
    assign weights1[61][673] = 16'b1111111111111011;
    assign weights1[61][674] = 16'b0000000000000001;
    assign weights1[61][675] = 16'b1111111111110100;
    assign weights1[61][676] = 16'b1111111111101100;
    assign weights1[61][677] = 16'b1111111111011110;
    assign weights1[61][678] = 16'b1111111111110101;
    assign weights1[61][679] = 16'b1111111111101101;
    assign weights1[61][680] = 16'b1111111111111001;
    assign weights1[61][681] = 16'b0000000000000100;
    assign weights1[61][682] = 16'b1111111111110011;
    assign weights1[61][683] = 16'b1111111111011111;
    assign weights1[61][684] = 16'b0000000000001101;
    assign weights1[61][685] = 16'b1111111111111010;
    assign weights1[61][686] = 16'b1111111111110110;
    assign weights1[61][687] = 16'b0000000000010110;
    assign weights1[61][688] = 16'b1111111111101101;
    assign weights1[61][689] = 16'b0000000000001111;
    assign weights1[61][690] = 16'b0000000000000010;
    assign weights1[61][691] = 16'b1111111111111100;
    assign weights1[61][692] = 16'b1111111111011100;
    assign weights1[61][693] = 16'b1111111111101110;
    assign weights1[61][694] = 16'b1111111111100101;
    assign weights1[61][695] = 16'b1111111111100100;
    assign weights1[61][696] = 16'b1111111111100011;
    assign weights1[61][697] = 16'b1111111111101011;
    assign weights1[61][698] = 16'b1111111111110001;
    assign weights1[61][699] = 16'b1111111111110101;
    assign weights1[61][700] = 16'b1111111111111111;
    assign weights1[61][701] = 16'b1111111111111101;
    assign weights1[61][702] = 16'b1111111111111100;
    assign weights1[61][703] = 16'b1111111111111001;
    assign weights1[61][704] = 16'b1111111111110101;
    assign weights1[61][705] = 16'b1111111111100000;
    assign weights1[61][706] = 16'b0000000000000100;
    assign weights1[61][707] = 16'b0000000000001011;
    assign weights1[61][708] = 16'b1111111111111110;
    assign weights1[61][709] = 16'b0000000000000010;
    assign weights1[61][710] = 16'b1111111111110010;
    assign weights1[61][711] = 16'b0000000000010010;
    assign weights1[61][712] = 16'b0000000000001010;
    assign weights1[61][713] = 16'b0000000000001001;
    assign weights1[61][714] = 16'b1111111111011100;
    assign weights1[61][715] = 16'b1111111111111001;
    assign weights1[61][716] = 16'b1111111111100011;
    assign weights1[61][717] = 16'b1111111111110111;
    assign weights1[61][718] = 16'b1111111111101001;
    assign weights1[61][719] = 16'b1111111111110010;
    assign weights1[61][720] = 16'b1111111111011111;
    assign weights1[61][721] = 16'b1111111111100000;
    assign weights1[61][722] = 16'b1111111111011000;
    assign weights1[61][723] = 16'b1111111111101001;
    assign weights1[61][724] = 16'b1111111111101000;
    assign weights1[61][725] = 16'b1111111111110000;
    assign weights1[61][726] = 16'b1111111111110001;
    assign weights1[61][727] = 16'b1111111111111011;
    assign weights1[61][728] = 16'b1111111111111111;
    assign weights1[61][729] = 16'b1111111111111100;
    assign weights1[61][730] = 16'b1111111111111000;
    assign weights1[61][731] = 16'b1111111111111010;
    assign weights1[61][732] = 16'b0000000000000001;
    assign weights1[61][733] = 16'b1111111111110111;
    assign weights1[61][734] = 16'b0000000000000001;
    assign weights1[61][735] = 16'b0000000000011010;
    assign weights1[61][736] = 16'b0000000000100100;
    assign weights1[61][737] = 16'b0000000000001100;
    assign weights1[61][738] = 16'b1111111111110010;
    assign weights1[61][739] = 16'b0000000000000110;
    assign weights1[61][740] = 16'b0000000000001010;
    assign weights1[61][741] = 16'b0000000000000000;
    assign weights1[61][742] = 16'b0000000000000101;
    assign weights1[61][743] = 16'b1111111111111010;
    assign weights1[61][744] = 16'b1111111111101110;
    assign weights1[61][745] = 16'b1111111111100000;
    assign weights1[61][746] = 16'b1111111111110000;
    assign weights1[61][747] = 16'b1111111111100101;
    assign weights1[61][748] = 16'b1111111111100111;
    assign weights1[61][749] = 16'b1111111111101000;
    assign weights1[61][750] = 16'b1111111111101001;
    assign weights1[61][751] = 16'b1111111111100100;
    assign weights1[61][752] = 16'b1111111111101101;
    assign weights1[61][753] = 16'b1111111111110011;
    assign weights1[61][754] = 16'b1111111111111000;
    assign weights1[61][755] = 16'b1111111111111100;
    assign weights1[61][756] = 16'b1111111111111111;
    assign weights1[61][757] = 16'b1111111111111110;
    assign weights1[61][758] = 16'b1111111111111010;
    assign weights1[61][759] = 16'b1111111111111101;
    assign weights1[61][760] = 16'b1111111111111100;
    assign weights1[61][761] = 16'b1111111111110100;
    assign weights1[61][762] = 16'b1111111111110011;
    assign weights1[61][763] = 16'b1111111111110011;
    assign weights1[61][764] = 16'b1111111111111100;
    assign weights1[61][765] = 16'b1111111111100111;
    assign weights1[61][766] = 16'b1111111111101110;
    assign weights1[61][767] = 16'b1111111111101111;
    assign weights1[61][768] = 16'b1111111111111000;
    assign weights1[61][769] = 16'b1111111111101110;
    assign weights1[61][770] = 16'b1111111111110011;
    assign weights1[61][771] = 16'b1111111111000011;
    assign weights1[61][772] = 16'b1111111111000111;
    assign weights1[61][773] = 16'b1111111111000111;
    assign weights1[61][774] = 16'b1111111111001100;
    assign weights1[61][775] = 16'b1111111111011101;
    assign weights1[61][776] = 16'b1111111111101001;
    assign weights1[61][777] = 16'b1111111111011010;
    assign weights1[61][778] = 16'b1111111111101010;
    assign weights1[61][779] = 16'b1111111111101111;
    assign weights1[61][780] = 16'b1111111111110010;
    assign weights1[61][781] = 16'b1111111111111101;
    assign weights1[61][782] = 16'b1111111111111110;
    assign weights1[61][783] = 16'b1111111111111110;
    assign weights1[62][0] = 16'b0000000000000001;
    assign weights1[62][1] = 16'b1111111111111111;
    assign weights1[62][2] = 16'b1111111111111111;
    assign weights1[62][3] = 16'b1111111111111101;
    assign weights1[62][4] = 16'b1111111111111011;
    assign weights1[62][5] = 16'b1111111111111011;
    assign weights1[62][6] = 16'b0000000000000111;
    assign weights1[62][7] = 16'b0000000000000100;
    assign weights1[62][8] = 16'b0000000000000101;
    assign weights1[62][9] = 16'b0000000000001000;
    assign weights1[62][10] = 16'b0000000000010001;
    assign weights1[62][11] = 16'b0000000000001100;
    assign weights1[62][12] = 16'b0000000000000011;
    assign weights1[62][13] = 16'b1111111111111110;
    assign weights1[62][14] = 16'b0000000000000000;
    assign weights1[62][15] = 16'b1111111111111101;
    assign weights1[62][16] = 16'b0000000000000000;
    assign weights1[62][17] = 16'b0000000000001101;
    assign weights1[62][18] = 16'b1111111111111101;
    assign weights1[62][19] = 16'b0000000000001011;
    assign weights1[62][20] = 16'b0000000000010101;
    assign weights1[62][21] = 16'b0000000000010000;
    assign weights1[62][22] = 16'b1111111111111111;
    assign weights1[62][23] = 16'b0000000000000011;
    assign weights1[62][24] = 16'b1111111111111111;
    assign weights1[62][25] = 16'b1111111111110011;
    assign weights1[62][26] = 16'b1111111111111001;
    assign weights1[62][27] = 16'b0000000000000001;
    assign weights1[62][28] = 16'b0000000000000001;
    assign weights1[62][29] = 16'b0000000000000000;
    assign weights1[62][30] = 16'b1111111111111001;
    assign weights1[62][31] = 16'b1111111111111100;
    assign weights1[62][32] = 16'b1111111111111110;
    assign weights1[62][33] = 16'b1111111111111111;
    assign weights1[62][34] = 16'b1111111111110001;
    assign weights1[62][35] = 16'b0000000000000001;
    assign weights1[62][36] = 16'b1111111111101110;
    assign weights1[62][37] = 16'b0000000000000010;
    assign weights1[62][38] = 16'b1111111111111010;
    assign weights1[62][39] = 16'b1111111111111010;
    assign weights1[62][40] = 16'b1111111111111101;
    assign weights1[62][41] = 16'b0000000000000000;
    assign weights1[62][42] = 16'b1111111111110010;
    assign weights1[62][43] = 16'b0000000000000111;
    assign weights1[62][44] = 16'b1111111111110101;
    assign weights1[62][45] = 16'b1111111111111011;
    assign weights1[62][46] = 16'b1111111111111101;
    assign weights1[62][47] = 16'b1111111111110111;
    assign weights1[62][48] = 16'b0000000000000011;
    assign weights1[62][49] = 16'b1111111111111011;
    assign weights1[62][50] = 16'b1111111111110110;
    assign weights1[62][51] = 16'b1111111111111110;
    assign weights1[62][52] = 16'b1111111111111110;
    assign weights1[62][53] = 16'b0000000000000001;
    assign weights1[62][54] = 16'b1111111111111111;
    assign weights1[62][55] = 16'b1111111111111110;
    assign weights1[62][56] = 16'b0000000000000010;
    assign weights1[62][57] = 16'b1111111111111101;
    assign weights1[62][58] = 16'b1111111111111001;
    assign weights1[62][59] = 16'b1111111111110100;
    assign weights1[62][60] = 16'b1111111111111011;
    assign weights1[62][61] = 16'b1111111111110010;
    assign weights1[62][62] = 16'b1111111111110000;
    assign weights1[62][63] = 16'b1111111111111011;
    assign weights1[62][64] = 16'b1111111111101110;
    assign weights1[62][65] = 16'b0000000000000101;
    assign weights1[62][66] = 16'b1111111111111000;
    assign weights1[62][67] = 16'b0000000000000000;
    assign weights1[62][68] = 16'b1111111111111100;
    assign weights1[62][69] = 16'b1111111111111000;
    assign weights1[62][70] = 16'b0000000000000001;
    assign weights1[62][71] = 16'b0000000000010001;
    assign weights1[62][72] = 16'b1111111111111111;
    assign weights1[62][73] = 16'b0000000000000100;
    assign weights1[62][74] = 16'b1111111111110111;
    assign weights1[62][75] = 16'b0000000000001010;
    assign weights1[62][76] = 16'b1111111111111101;
    assign weights1[62][77] = 16'b0000000000000100;
    assign weights1[62][78] = 16'b1111111111111010;
    assign weights1[62][79] = 16'b0000000000000111;
    assign weights1[62][80] = 16'b0000000000001100;
    assign weights1[62][81] = 16'b0000000000001000;
    assign weights1[62][82] = 16'b0000000000000101;
    assign weights1[62][83] = 16'b0000000000000011;
    assign weights1[62][84] = 16'b0000000000000011;
    assign weights1[62][85] = 16'b0000000000000011;
    assign weights1[62][86] = 16'b1111111111110110;
    assign weights1[62][87] = 16'b1111111111111001;
    assign weights1[62][88] = 16'b1111111111111111;
    assign weights1[62][89] = 16'b1111111111110111;
    assign weights1[62][90] = 16'b1111111111111100;
    assign weights1[62][91] = 16'b0000000000000001;
    assign weights1[62][92] = 16'b0000000000001100;
    assign weights1[62][93] = 16'b1111111111111111;
    assign weights1[62][94] = 16'b0000000000001001;
    assign weights1[62][95] = 16'b0000000000000011;
    assign weights1[62][96] = 16'b1111111111111011;
    assign weights1[62][97] = 16'b1111111111111110;
    assign weights1[62][98] = 16'b1111111111110110;
    assign weights1[62][99] = 16'b1111111111110101;
    assign weights1[62][100] = 16'b1111111111111110;
    assign weights1[62][101] = 16'b0000000000000101;
    assign weights1[62][102] = 16'b1111111111110010;
    assign weights1[62][103] = 16'b1111111111111100;
    assign weights1[62][104] = 16'b0000000000000010;
    assign weights1[62][105] = 16'b0000000000000011;
    assign weights1[62][106] = 16'b0000000000000001;
    assign weights1[62][107] = 16'b0000000000001101;
    assign weights1[62][108] = 16'b0000000000010001;
    assign weights1[62][109] = 16'b0000000000000101;
    assign weights1[62][110] = 16'b0000000000001110;
    assign weights1[62][111] = 16'b0000000000001100;
    assign weights1[62][112] = 16'b1111111111111110;
    assign weights1[62][113] = 16'b1111111111111100;
    assign weights1[62][114] = 16'b1111111111111101;
    assign weights1[62][115] = 16'b0000000000000001;
    assign weights1[62][116] = 16'b1111111111111110;
    assign weights1[62][117] = 16'b1111111111111100;
    assign weights1[62][118] = 16'b0000000000000000;
    assign weights1[62][119] = 16'b0000000000001011;
    assign weights1[62][120] = 16'b1111111111111001;
    assign weights1[62][121] = 16'b1111111111101111;
    assign weights1[62][122] = 16'b0000000000000010;
    assign weights1[62][123] = 16'b0000000000000110;
    assign weights1[62][124] = 16'b0000000000000001;
    assign weights1[62][125] = 16'b1111111111111100;
    assign weights1[62][126] = 16'b0000000000001100;
    assign weights1[62][127] = 16'b0000000000001110;
    assign weights1[62][128] = 16'b1111111111110011;
    assign weights1[62][129] = 16'b0000000000001110;
    assign weights1[62][130] = 16'b0000000000000000;
    assign weights1[62][131] = 16'b0000000000001111;
    assign weights1[62][132] = 16'b1111111111110100;
    assign weights1[62][133] = 16'b1111111111111000;
    assign weights1[62][134] = 16'b1111111111100000;
    assign weights1[62][135] = 16'b0000000000000000;
    assign weights1[62][136] = 16'b1111111111101101;
    assign weights1[62][137] = 16'b1111111111110111;
    assign weights1[62][138] = 16'b1111111111111101;
    assign weights1[62][139] = 16'b0000000000000000;
    assign weights1[62][140] = 16'b1111111111111111;
    assign weights1[62][141] = 16'b1111111111110110;
    assign weights1[62][142] = 16'b1111111111111110;
    assign weights1[62][143] = 16'b1111111111111001;
    assign weights1[62][144] = 16'b1111111111110111;
    assign weights1[62][145] = 16'b0000000000001101;
    assign weights1[62][146] = 16'b1111111111110000;
    assign weights1[62][147] = 16'b0000000000001010;
    assign weights1[62][148] = 16'b0000000000001101;
    assign weights1[62][149] = 16'b1111111111111011;
    assign weights1[62][150] = 16'b1111111111110100;
    assign weights1[62][151] = 16'b0000000000000111;
    assign weights1[62][152] = 16'b1111111111110110;
    assign weights1[62][153] = 16'b0000000000000100;
    assign weights1[62][154] = 16'b1111111111110011;
    assign weights1[62][155] = 16'b0000000000000010;
    assign weights1[62][156] = 16'b1111111111111110;
    assign weights1[62][157] = 16'b1111111111111000;
    assign weights1[62][158] = 16'b1111111111110100;
    assign weights1[62][159] = 16'b0000000000000000;
    assign weights1[62][160] = 16'b1111111111110110;
    assign weights1[62][161] = 16'b1111111111111010;
    assign weights1[62][162] = 16'b1111111111110100;
    assign weights1[62][163] = 16'b1111111111111100;
    assign weights1[62][164] = 16'b1111111111110101;
    assign weights1[62][165] = 16'b0000000000001100;
    assign weights1[62][166] = 16'b1111111111110100;
    assign weights1[62][167] = 16'b1111111111110001;
    assign weights1[62][168] = 16'b0000000000000011;
    assign weights1[62][169] = 16'b0000000000000011;
    assign weights1[62][170] = 16'b1111111111111100;
    assign weights1[62][171] = 16'b0000000000001101;
    assign weights1[62][172] = 16'b1111111111111100;
    assign weights1[62][173] = 16'b0000000000001110;
    assign weights1[62][174] = 16'b0000000000000010;
    assign weights1[62][175] = 16'b1111111111111101;
    assign weights1[62][176] = 16'b1111111111111110;
    assign weights1[62][177] = 16'b0000000000000001;
    assign weights1[62][178] = 16'b1111111111111001;
    assign weights1[62][179] = 16'b0000000000000011;
    assign weights1[62][180] = 16'b1111111111111001;
    assign weights1[62][181] = 16'b1111111111111011;
    assign weights1[62][182] = 16'b1111111111110010;
    assign weights1[62][183] = 16'b1111111111110111;
    assign weights1[62][184] = 16'b0000000000000101;
    assign weights1[62][185] = 16'b1111111111111010;
    assign weights1[62][186] = 16'b0000000000000100;
    assign weights1[62][187] = 16'b1111111111110110;
    assign weights1[62][188] = 16'b1111111111110000;
    assign weights1[62][189] = 16'b1111111111111101;
    assign weights1[62][190] = 16'b1111111111110110;
    assign weights1[62][191] = 16'b1111111111110101;
    assign weights1[62][192] = 16'b1111111111011100;
    assign weights1[62][193] = 16'b1111111111110000;
    assign weights1[62][194] = 16'b1111111111111100;
    assign weights1[62][195] = 16'b1111111111110011;
    assign weights1[62][196] = 16'b1111111111111111;
    assign weights1[62][197] = 16'b0000000000000001;
    assign weights1[62][198] = 16'b0000000000010000;
    assign weights1[62][199] = 16'b0000000000000001;
    assign weights1[62][200] = 16'b1111111111111010;
    assign weights1[62][201] = 16'b1111111111101110;
    assign weights1[62][202] = 16'b1111111111100111;
    assign weights1[62][203] = 16'b0000000000000110;
    assign weights1[62][204] = 16'b1111111111111111;
    assign weights1[62][205] = 16'b1111111111111001;
    assign weights1[62][206] = 16'b1111111111111001;
    assign weights1[62][207] = 16'b0000000000000101;
    assign weights1[62][208] = 16'b0000000000000001;
    assign weights1[62][209] = 16'b0000000000000011;
    assign weights1[62][210] = 16'b1111111111111111;
    assign weights1[62][211] = 16'b1111111111110010;
    assign weights1[62][212] = 16'b0000000000001011;
    assign weights1[62][213] = 16'b1111111111101111;
    assign weights1[62][214] = 16'b1111111111110100;
    assign weights1[62][215] = 16'b1111111111111010;
    assign weights1[62][216] = 16'b1111111111110110;
    assign weights1[62][217] = 16'b1111111111111101;
    assign weights1[62][218] = 16'b1111111111101010;
    assign weights1[62][219] = 16'b1111111111011111;
    assign weights1[62][220] = 16'b0000000000011110;
    assign weights1[62][221] = 16'b1111111111111110;
    assign weights1[62][222] = 16'b1111111111101010;
    assign weights1[62][223] = 16'b1111111111101110;
    assign weights1[62][224] = 16'b1111111111111000;
    assign weights1[62][225] = 16'b1111111111111110;
    assign weights1[62][226] = 16'b0000000000000010;
    assign weights1[62][227] = 16'b1111111111111100;
    assign weights1[62][228] = 16'b1111111111111000;
    assign weights1[62][229] = 16'b1111111111111011;
    assign weights1[62][230] = 16'b0000000000000111;
    assign weights1[62][231] = 16'b1111111111111000;
    assign weights1[62][232] = 16'b0000000000001001;
    assign weights1[62][233] = 16'b0000000000000110;
    assign weights1[62][234] = 16'b1111111111111110;
    assign weights1[62][235] = 16'b1111111111110111;
    assign weights1[62][236] = 16'b1111111111111101;
    assign weights1[62][237] = 16'b1111111111101010;
    assign weights1[62][238] = 16'b0000000000000001;
    assign weights1[62][239] = 16'b1111111111110010;
    assign weights1[62][240] = 16'b1111111111110011;
    assign weights1[62][241] = 16'b1111111111111001;
    assign weights1[62][242] = 16'b1111111111101011;
    assign weights1[62][243] = 16'b1111111111110000;
    assign weights1[62][244] = 16'b1111111111101110;
    assign weights1[62][245] = 16'b1111111111111010;
    assign weights1[62][246] = 16'b1111111111110001;
    assign weights1[62][247] = 16'b1111111111111000;
    assign weights1[62][248] = 16'b1111111111100000;
    assign weights1[62][249] = 16'b1111111111111010;
    assign weights1[62][250] = 16'b1111111111110001;
    assign weights1[62][251] = 16'b1111111111101000;
    assign weights1[62][252] = 16'b1111111111111011;
    assign weights1[62][253] = 16'b1111111111111110;
    assign weights1[62][254] = 16'b0000000000001110;
    assign weights1[62][255] = 16'b0000000000000010;
    assign weights1[62][256] = 16'b0000000000000011;
    assign weights1[62][257] = 16'b1111111111111010;
    assign weights1[62][258] = 16'b1111111111110101;
    assign weights1[62][259] = 16'b1111111111111101;
    assign weights1[62][260] = 16'b1111111111111000;
    assign weights1[62][261] = 16'b1111111111111100;
    assign weights1[62][262] = 16'b0000000000000010;
    assign weights1[62][263] = 16'b0000000000001010;
    assign weights1[62][264] = 16'b1111111111111100;
    assign weights1[62][265] = 16'b1111111111111001;
    assign weights1[62][266] = 16'b0000000000001010;
    assign weights1[62][267] = 16'b1111111111111110;
    assign weights1[62][268] = 16'b1111111111111111;
    assign weights1[62][269] = 16'b1111111111111010;
    assign weights1[62][270] = 16'b0000000000000001;
    assign weights1[62][271] = 16'b1111111111110111;
    assign weights1[62][272] = 16'b0000000000001110;
    assign weights1[62][273] = 16'b1111111111101111;
    assign weights1[62][274] = 16'b1111111111111100;
    assign weights1[62][275] = 16'b1111111111100101;
    assign weights1[62][276] = 16'b1111111111101011;
    assign weights1[62][277] = 16'b1111111111011011;
    assign weights1[62][278] = 16'b1111111111011101;
    assign weights1[62][279] = 16'b1111111111100001;
    assign weights1[62][280] = 16'b1111111111111110;
    assign weights1[62][281] = 16'b1111111111111000;
    assign weights1[62][282] = 16'b1111111111110100;
    assign weights1[62][283] = 16'b0000000000001011;
    assign weights1[62][284] = 16'b0000000000000111;
    assign weights1[62][285] = 16'b0000000000000010;
    assign weights1[62][286] = 16'b0000000000001000;
    assign weights1[62][287] = 16'b1111111111110000;
    assign weights1[62][288] = 16'b0000000000010110;
    assign weights1[62][289] = 16'b0000000000000010;
    assign weights1[62][290] = 16'b0000000000001000;
    assign weights1[62][291] = 16'b0000000000000010;
    assign weights1[62][292] = 16'b0000000000000010;
    assign weights1[62][293] = 16'b1111111111111100;
    assign weights1[62][294] = 16'b0000000000000011;
    assign weights1[62][295] = 16'b0000000000001001;
    assign weights1[62][296] = 16'b1111111111111101;
    assign weights1[62][297] = 16'b0000000000000111;
    assign weights1[62][298] = 16'b0000000000000100;
    assign weights1[62][299] = 16'b1111111111111111;
    assign weights1[62][300] = 16'b1111111111110101;
    assign weights1[62][301] = 16'b0000000000000111;
    assign weights1[62][302] = 16'b1111111111111000;
    assign weights1[62][303] = 16'b0000000000010000;
    assign weights1[62][304] = 16'b1111111111111111;
    assign weights1[62][305] = 16'b1111111111101000;
    assign weights1[62][306] = 16'b1111111111110101;
    assign weights1[62][307] = 16'b1111111111110000;
    assign weights1[62][308] = 16'b1111111111111100;
    assign weights1[62][309] = 16'b1111111111111001;
    assign weights1[62][310] = 16'b0000000000000110;
    assign weights1[62][311] = 16'b1111111111111000;
    assign weights1[62][312] = 16'b1111111111101010;
    assign weights1[62][313] = 16'b1111111111111000;
    assign weights1[62][314] = 16'b1111111111111110;
    assign weights1[62][315] = 16'b1111111111110111;
    assign weights1[62][316] = 16'b1111111111111001;
    assign weights1[62][317] = 16'b1111111111110010;
    assign weights1[62][318] = 16'b1111111111110101;
    assign weights1[62][319] = 16'b1111111111111101;
    assign weights1[62][320] = 16'b1111111111110110;
    assign weights1[62][321] = 16'b1111111111110110;
    assign weights1[62][322] = 16'b1111111111111011;
    assign weights1[62][323] = 16'b1111111111111001;
    assign weights1[62][324] = 16'b1111111111111100;
    assign weights1[62][325] = 16'b1111111111110011;
    assign weights1[62][326] = 16'b1111111111111101;
    assign weights1[62][327] = 16'b0000000000000000;
    assign weights1[62][328] = 16'b1111111111111011;
    assign weights1[62][329] = 16'b1111111111111001;
    assign weights1[62][330] = 16'b1111111111110001;
    assign weights1[62][331] = 16'b1111111111111111;
    assign weights1[62][332] = 16'b1111111111100010;
    assign weights1[62][333] = 16'b1111111111110010;
    assign weights1[62][334] = 16'b1111111111011010;
    assign weights1[62][335] = 16'b0000000000000000;
    assign weights1[62][336] = 16'b1111111111110101;
    assign weights1[62][337] = 16'b0000000000000100;
    assign weights1[62][338] = 16'b1111111111110111;
    assign weights1[62][339] = 16'b0000000000001000;
    assign weights1[62][340] = 16'b1111111111101100;
    assign weights1[62][341] = 16'b1111111111110101;
    assign weights1[62][342] = 16'b0000000000000010;
    assign weights1[62][343] = 16'b0000000000010010;
    assign weights1[62][344] = 16'b0000000000000011;
    assign weights1[62][345] = 16'b1111111111110111;
    assign weights1[62][346] = 16'b1111111111111100;
    assign weights1[62][347] = 16'b0000000000000110;
    assign weights1[62][348] = 16'b1111111111111010;
    assign weights1[62][349] = 16'b1111111111111110;
    assign weights1[62][350] = 16'b0000000000000010;
    assign weights1[62][351] = 16'b0000000000000010;
    assign weights1[62][352] = 16'b0000000000001000;
    assign weights1[62][353] = 16'b1111111111111011;
    assign weights1[62][354] = 16'b0000000000000010;
    assign weights1[62][355] = 16'b1111111111110101;
    assign weights1[62][356] = 16'b0000000000001100;
    assign weights1[62][357] = 16'b1111111111111000;
    assign weights1[62][358] = 16'b0000000000000100;
    assign weights1[62][359] = 16'b1111111111110011;
    assign weights1[62][360] = 16'b0000000000001100;
    assign weights1[62][361] = 16'b1111111111111001;
    assign weights1[62][362] = 16'b0000000000001001;
    assign weights1[62][363] = 16'b0000000000001111;
    assign weights1[62][364] = 16'b0000000000000111;
    assign weights1[62][365] = 16'b0000000000001001;
    assign weights1[62][366] = 16'b0000000000000110;
    assign weights1[62][367] = 16'b1111111111111110;
    assign weights1[62][368] = 16'b1111111111111010;
    assign weights1[62][369] = 16'b0000000000001000;
    assign weights1[62][370] = 16'b0000000000010000;
    assign weights1[62][371] = 16'b1111111111111100;
    assign weights1[62][372] = 16'b1111111111111101;
    assign weights1[62][373] = 16'b1111111111101110;
    assign weights1[62][374] = 16'b1111111111110111;
    assign weights1[62][375] = 16'b0000000000000001;
    assign weights1[62][376] = 16'b0000000000000010;
    assign weights1[62][377] = 16'b0000000000000010;
    assign weights1[62][378] = 16'b1111111111111001;
    assign weights1[62][379] = 16'b1111111111110001;
    assign weights1[62][380] = 16'b1111111111111000;
    assign weights1[62][381] = 16'b1111111111111100;
    assign weights1[62][382] = 16'b1111111111110111;
    assign weights1[62][383] = 16'b1111111111111011;
    assign weights1[62][384] = 16'b1111111111111000;
    assign weights1[62][385] = 16'b0000000000000101;
    assign weights1[62][386] = 16'b0000000000000110;
    assign weights1[62][387] = 16'b0000000000010011;
    assign weights1[62][388] = 16'b0000000000001101;
    assign weights1[62][389] = 16'b0000000000011010;
    assign weights1[62][390] = 16'b0000000000001011;
    assign weights1[62][391] = 16'b0000000000001001;
    assign weights1[62][392] = 16'b0000000000001100;
    assign weights1[62][393] = 16'b1111111111111010;
    assign weights1[62][394] = 16'b1111111111110000;
    assign weights1[62][395] = 16'b0000000000000010;
    assign weights1[62][396] = 16'b1111111111110110;
    assign weights1[62][397] = 16'b1111111111111110;
    assign weights1[62][398] = 16'b1111111111110100;
    assign weights1[62][399] = 16'b1111111111111000;
    assign weights1[62][400] = 16'b1111111111110100;
    assign weights1[62][401] = 16'b1111111111110111;
    assign weights1[62][402] = 16'b1111111111111100;
    assign weights1[62][403] = 16'b1111111111111101;
    assign weights1[62][404] = 16'b1111111111101110;
    assign weights1[62][405] = 16'b1111111111110111;
    assign weights1[62][406] = 16'b0000000000000100;
    assign weights1[62][407] = 16'b1111111111110101;
    assign weights1[62][408] = 16'b0000000000000000;
    assign weights1[62][409] = 16'b1111111111110111;
    assign weights1[62][410] = 16'b0000000000000101;
    assign weights1[62][411] = 16'b1111111111111111;
    assign weights1[62][412] = 16'b0000000000000010;
    assign weights1[62][413] = 16'b1111111111111101;
    assign weights1[62][414] = 16'b0000000000010010;
    assign weights1[62][415] = 16'b0000000000000110;
    assign weights1[62][416] = 16'b0000000000001111;
    assign weights1[62][417] = 16'b0000000000001010;
    assign weights1[62][418] = 16'b0000000000101011;
    assign weights1[62][419] = 16'b0000000000001111;
    assign weights1[62][420] = 16'b0000000000011001;
    assign weights1[62][421] = 16'b0000000000001011;
    assign weights1[62][422] = 16'b1111111111111100;
    assign weights1[62][423] = 16'b1111111111110111;
    assign weights1[62][424] = 16'b1111111111100101;
    assign weights1[62][425] = 16'b1111111111101011;
    assign weights1[62][426] = 16'b0000000000000001;
    assign weights1[62][427] = 16'b1111111111110001;
    assign weights1[62][428] = 16'b1111111111111010;
    assign weights1[62][429] = 16'b1111111111110100;
    assign weights1[62][430] = 16'b0000000000000111;
    assign weights1[62][431] = 16'b1111111111110010;
    assign weights1[62][432] = 16'b1111111111110010;
    assign weights1[62][433] = 16'b1111111111111111;
    assign weights1[62][434] = 16'b1111111111101111;
    assign weights1[62][435] = 16'b1111111111110110;
    assign weights1[62][436] = 16'b1111111111110000;
    assign weights1[62][437] = 16'b1111111111110010;
    assign weights1[62][438] = 16'b1111111111110101;
    assign weights1[62][439] = 16'b0000000000010000;
    assign weights1[62][440] = 16'b0000000000010100;
    assign weights1[62][441] = 16'b0000000000001110;
    assign weights1[62][442] = 16'b0000000000011010;
    assign weights1[62][443] = 16'b0000000000000101;
    assign weights1[62][444] = 16'b0000000000011100;
    assign weights1[62][445] = 16'b0000000000101000;
    assign weights1[62][446] = 16'b0000000000011010;
    assign weights1[62][447] = 16'b0000000000001110;
    assign weights1[62][448] = 16'b0000000000010110;
    assign weights1[62][449] = 16'b0000000000010011;
    assign weights1[62][450] = 16'b0000000000000101;
    assign weights1[62][451] = 16'b0000000000000111;
    assign weights1[62][452] = 16'b0000000000001011;
    assign weights1[62][453] = 16'b1111111111110110;
    assign weights1[62][454] = 16'b1111111111110110;
    assign weights1[62][455] = 16'b0000000000000110;
    assign weights1[62][456] = 16'b1111111111111100;
    assign weights1[62][457] = 16'b0000000000000000;
    assign weights1[62][458] = 16'b1111111111111110;
    assign weights1[62][459] = 16'b1111111111110011;
    assign weights1[62][460] = 16'b1111111111110001;
    assign weights1[62][461] = 16'b0000000000000001;
    assign weights1[62][462] = 16'b1111111111111110;
    assign weights1[62][463] = 16'b0000000000000000;
    assign weights1[62][464] = 16'b0000000000000000;
    assign weights1[62][465] = 16'b0000000000000010;
    assign weights1[62][466] = 16'b0000000000001110;
    assign weights1[62][467] = 16'b0000000000010010;
    assign weights1[62][468] = 16'b0000000000001100;
    assign weights1[62][469] = 16'b0000000000100101;
    assign weights1[62][470] = 16'b0000000000010001;
    assign weights1[62][471] = 16'b0000000000001100;
    assign weights1[62][472] = 16'b0000000000011010;
    assign weights1[62][473] = 16'b0000000000011100;
    assign weights1[62][474] = 16'b0000000000011000;
    assign weights1[62][475] = 16'b0000000000000110;
    assign weights1[62][476] = 16'b0000000000011101;
    assign weights1[62][477] = 16'b0000000000010110;
    assign weights1[62][478] = 16'b0000000000010110;
    assign weights1[62][479] = 16'b0000000000001001;
    assign weights1[62][480] = 16'b0000000000100011;
    assign weights1[62][481] = 16'b0000000000001100;
    assign weights1[62][482] = 16'b1111111111111111;
    assign weights1[62][483] = 16'b1111111111110101;
    assign weights1[62][484] = 16'b1111111111111100;
    assign weights1[62][485] = 16'b1111111111110110;
    assign weights1[62][486] = 16'b0000000000000110;
    assign weights1[62][487] = 16'b0000000000001010;
    assign weights1[62][488] = 16'b0000000000000110;
    assign weights1[62][489] = 16'b0000000000001001;
    assign weights1[62][490] = 16'b0000000000000010;
    assign weights1[62][491] = 16'b0000000000001101;
    assign weights1[62][492] = 16'b0000000000010101;
    assign weights1[62][493] = 16'b0000000000100011;
    assign weights1[62][494] = 16'b0000000000011000;
    assign weights1[62][495] = 16'b0000000000000111;
    assign weights1[62][496] = 16'b0000000000011010;
    assign weights1[62][497] = 16'b0000000000001001;
    assign weights1[62][498] = 16'b0000000000001001;
    assign weights1[62][499] = 16'b1111111111111111;
    assign weights1[62][500] = 16'b0000000000000001;
    assign weights1[62][501] = 16'b0000000000011011;
    assign weights1[62][502] = 16'b0000000000001101;
    assign weights1[62][503] = 16'b0000000000001001;
    assign weights1[62][504] = 16'b0000000000010101;
    assign weights1[62][505] = 16'b0000000000011001;
    assign weights1[62][506] = 16'b0000000000100001;
    assign weights1[62][507] = 16'b0000000000101010;
    assign weights1[62][508] = 16'b0000000000010101;
    assign weights1[62][509] = 16'b0000000000011000;
    assign weights1[62][510] = 16'b0000000000011011;
    assign weights1[62][511] = 16'b0000000000001111;
    assign weights1[62][512] = 16'b0000000000010100;
    assign weights1[62][513] = 16'b0000000000010111;
    assign weights1[62][514] = 16'b0000000000010110;
    assign weights1[62][515] = 16'b0000000000010010;
    assign weights1[62][516] = 16'b0000000000011001;
    assign weights1[62][517] = 16'b0000000000011000;
    assign weights1[62][518] = 16'b0000000000101010;
    assign weights1[62][519] = 16'b0000000000011110;
    assign weights1[62][520] = 16'b0000000000101001;
    assign weights1[62][521] = 16'b0000000000010110;
    assign weights1[62][522] = 16'b0000000000001111;
    assign weights1[62][523] = 16'b0000000000011101;
    assign weights1[62][524] = 16'b0000000000001001;
    assign weights1[62][525] = 16'b0000000000000100;
    assign weights1[62][526] = 16'b0000000000010010;
    assign weights1[62][527] = 16'b1111111111111111;
    assign weights1[62][528] = 16'b0000000000011001;
    assign weights1[62][529] = 16'b0000000000010010;
    assign weights1[62][530] = 16'b0000000000001000;
    assign weights1[62][531] = 16'b1111111111110001;
    assign weights1[62][532] = 16'b0000000000010101;
    assign weights1[62][533] = 16'b0000000000001001;
    assign weights1[62][534] = 16'b0000000000011100;
    assign weights1[62][535] = 16'b0000000000010101;
    assign weights1[62][536] = 16'b0000000000111011;
    assign weights1[62][537] = 16'b0000000000010110;
    assign weights1[62][538] = 16'b0000000000101000;
    assign weights1[62][539] = 16'b0000000000100111;
    assign weights1[62][540] = 16'b0000000000011111;
    assign weights1[62][541] = 16'b0000000000011101;
    assign weights1[62][542] = 16'b0000000000100000;
    assign weights1[62][543] = 16'b0000000000011001;
    assign weights1[62][544] = 16'b0000000000011100;
    assign weights1[62][545] = 16'b0000000000100001;
    assign weights1[62][546] = 16'b0000000000010111;
    assign weights1[62][547] = 16'b0000000000010000;
    assign weights1[62][548] = 16'b0000000000010110;
    assign weights1[62][549] = 16'b0000000000011100;
    assign weights1[62][550] = 16'b0000000000101001;
    assign weights1[62][551] = 16'b0000000000010011;
    assign weights1[62][552] = 16'b0000000000011010;
    assign weights1[62][553] = 16'b0000000000001100;
    assign weights1[62][554] = 16'b0000000000100000;
    assign weights1[62][555] = 16'b1111111111110101;
    assign weights1[62][556] = 16'b0000000000000000;
    assign weights1[62][557] = 16'b1111111111101010;
    assign weights1[62][558] = 16'b1111111111101101;
    assign weights1[62][559] = 16'b1111111111010111;
    assign weights1[62][560] = 16'b0000000000011111;
    assign weights1[62][561] = 16'b0000000000001110;
    assign weights1[62][562] = 16'b0000000000001110;
    assign weights1[62][563] = 16'b0000000000010000;
    assign weights1[62][564] = 16'b0000000000011111;
    assign weights1[62][565] = 16'b0000000000010001;
    assign weights1[62][566] = 16'b0000000000010001;
    assign weights1[62][567] = 16'b0000000000011110;
    assign weights1[62][568] = 16'b0000000000011111;
    assign weights1[62][569] = 16'b0000000000001110;
    assign weights1[62][570] = 16'b0000000000011101;
    assign weights1[62][571] = 16'b0000000000010111;
    assign weights1[62][572] = 16'b0000000000010011;
    assign weights1[62][573] = 16'b0000000000011100;
    assign weights1[62][574] = 16'b0000000000011010;
    assign weights1[62][575] = 16'b1111111111111100;
    assign weights1[62][576] = 16'b0000000000101000;
    assign weights1[62][577] = 16'b0000000000000010;
    assign weights1[62][578] = 16'b0000000000011111;
    assign weights1[62][579] = 16'b0000000000001001;
    assign weights1[62][580] = 16'b0000000000001100;
    assign weights1[62][581] = 16'b0000000000011001;
    assign weights1[62][582] = 16'b0000000000001100;
    assign weights1[62][583] = 16'b1111111111110100;
    assign weights1[62][584] = 16'b1111111111100010;
    assign weights1[62][585] = 16'b1111111111000000;
    assign weights1[62][586] = 16'b1111111111000011;
    assign weights1[62][587] = 16'b1111111111001011;
    assign weights1[62][588] = 16'b0000000000000010;
    assign weights1[62][589] = 16'b0000000000001101;
    assign weights1[62][590] = 16'b1111111111111001;
    assign weights1[62][591] = 16'b1111111111111000;
    assign weights1[62][592] = 16'b0000000000001100;
    assign weights1[62][593] = 16'b0000000000010111;
    assign weights1[62][594] = 16'b1111111111111000;
    assign weights1[62][595] = 16'b0000000000001001;
    assign weights1[62][596] = 16'b0000000000000011;
    assign weights1[62][597] = 16'b0000000000010100;
    assign weights1[62][598] = 16'b0000000000000101;
    assign weights1[62][599] = 16'b0000000000001011;
    assign weights1[62][600] = 16'b0000000000001001;
    assign weights1[62][601] = 16'b1111111111110101;
    assign weights1[62][602] = 16'b0000000000001011;
    assign weights1[62][603] = 16'b0000000000000111;
    assign weights1[62][604] = 16'b0000000000010100;
    assign weights1[62][605] = 16'b1111111111111001;
    assign weights1[62][606] = 16'b1111111111101110;
    assign weights1[62][607] = 16'b0000000000011000;
    assign weights1[62][608] = 16'b1111111111110001;
    assign weights1[62][609] = 16'b1111111111110000;
    assign weights1[62][610] = 16'b1111111111100000;
    assign weights1[62][611] = 16'b1111111111000011;
    assign weights1[62][612] = 16'b1111111110110100;
    assign weights1[62][613] = 16'b1111111111000110;
    assign weights1[62][614] = 16'b1111111110111010;
    assign weights1[62][615] = 16'b1111111111010011;
    assign weights1[62][616] = 16'b1111111111101110;
    assign weights1[62][617] = 16'b1111111111101111;
    assign weights1[62][618] = 16'b1111111111100011;
    assign weights1[62][619] = 16'b1111111111011111;
    assign weights1[62][620] = 16'b0000000000000010;
    assign weights1[62][621] = 16'b1111111111111011;
    assign weights1[62][622] = 16'b0000000000000000;
    assign weights1[62][623] = 16'b0000000000000000;
    assign weights1[62][624] = 16'b1111111111111110;
    assign weights1[62][625] = 16'b1111111111110010;
    assign weights1[62][626] = 16'b0000000000001011;
    assign weights1[62][627] = 16'b1111111111111101;
    assign weights1[62][628] = 16'b0000000000001001;
    assign weights1[62][629] = 16'b1111111111111011;
    assign weights1[62][630] = 16'b0000000000001110;
    assign weights1[62][631] = 16'b1111111111110100;
    assign weights1[62][632] = 16'b1111111111100111;
    assign weights1[62][633] = 16'b1111111111001111;
    assign weights1[62][634] = 16'b1111111110111110;
    assign weights1[62][635] = 16'b1111111111000001;
    assign weights1[62][636] = 16'b1111111110110000;
    assign weights1[62][637] = 16'b1111111110011101;
    assign weights1[62][638] = 16'b1111111110011111;
    assign weights1[62][639] = 16'b1111111110100000;
    assign weights1[62][640] = 16'b1111111110011100;
    assign weights1[62][641] = 16'b1111111111000000;
    assign weights1[62][642] = 16'b1111111111001010;
    assign weights1[62][643] = 16'b1111111111011010;
    assign weights1[62][644] = 16'b1111111111101010;
    assign weights1[62][645] = 16'b1111111111100100;
    assign weights1[62][646] = 16'b1111111111010001;
    assign weights1[62][647] = 16'b1111111111010011;
    assign weights1[62][648] = 16'b1111111110111101;
    assign weights1[62][649] = 16'b1111111111001011;
    assign weights1[62][650] = 16'b1111111111011010;
    assign weights1[62][651] = 16'b1111111111010100;
    assign weights1[62][652] = 16'b1111111111000100;
    assign weights1[62][653] = 16'b1111111111001100;
    assign weights1[62][654] = 16'b1111111111101101;
    assign weights1[62][655] = 16'b1111111111001011;
    assign weights1[62][656] = 16'b1111111110110010;
    assign weights1[62][657] = 16'b1111111110100110;
    assign weights1[62][658] = 16'b1111111110011000;
    assign weights1[62][659] = 16'b1111111101111001;
    assign weights1[62][660] = 16'b1111111100100100;
    assign weights1[62][661] = 16'b1111111101000011;
    assign weights1[62][662] = 16'b1111111101101011;
    assign weights1[62][663] = 16'b1111111101110000;
    assign weights1[62][664] = 16'b1111111101111000;
    assign weights1[62][665] = 16'b1111111110011100;
    assign weights1[62][666] = 16'b1111111110100110;
    assign weights1[62][667] = 16'b1111111110111000;
    assign weights1[62][668] = 16'b1111111110101011;
    assign weights1[62][669] = 16'b1111111111001000;
    assign weights1[62][670] = 16'b1111111111010100;
    assign weights1[62][671] = 16'b1111111111100011;
    assign weights1[62][672] = 16'b1111111111110100;
    assign weights1[62][673] = 16'b1111111111101000;
    assign weights1[62][674] = 16'b1111111111011011;
    assign weights1[62][675] = 16'b1111111111001001;
    assign weights1[62][676] = 16'b1111111111001000;
    assign weights1[62][677] = 16'b1111111110110100;
    assign weights1[62][678] = 16'b1111111110110100;
    assign weights1[62][679] = 16'b1111111110100001;
    assign weights1[62][680] = 16'b1111111110010010;
    assign weights1[62][681] = 16'b1111111101110100;
    assign weights1[62][682] = 16'b1111111101011011;
    assign weights1[62][683] = 16'b1111111101011100;
    assign weights1[62][684] = 16'b1111111101110001;
    assign weights1[62][685] = 16'b1111111101110011;
    assign weights1[62][686] = 16'b1111111101100101;
    assign weights1[62][687] = 16'b1111111101110001;
    assign weights1[62][688] = 16'b1111111101111110;
    assign weights1[62][689] = 16'b1111111110011010;
    assign weights1[62][690] = 16'b1111111110100111;
    assign weights1[62][691] = 16'b1111111110101000;
    assign weights1[62][692] = 16'b1111111110001011;
    assign weights1[62][693] = 16'b1111111110101110;
    assign weights1[62][694] = 16'b1111111110110100;
    assign weights1[62][695] = 16'b1111111111000101;
    assign weights1[62][696] = 16'b1111111111001000;
    assign weights1[62][697] = 16'b1111111111011010;
    assign weights1[62][698] = 16'b1111111111100100;
    assign weights1[62][699] = 16'b1111111111101100;
    assign weights1[62][700] = 16'b1111111111110110;
    assign weights1[62][701] = 16'b1111111111110011;
    assign weights1[62][702] = 16'b1111111111101011;
    assign weights1[62][703] = 16'b1111111111011101;
    assign weights1[62][704] = 16'b1111111111010011;
    assign weights1[62][705] = 16'b1111111110111111;
    assign weights1[62][706] = 16'b1111111110111101;
    assign weights1[62][707] = 16'b1111111110110111;
    assign weights1[62][708] = 16'b1111111110110000;
    assign weights1[62][709] = 16'b1111111110011011;
    assign weights1[62][710] = 16'b1111111110110100;
    assign weights1[62][711] = 16'b1111111110111000;
    assign weights1[62][712] = 16'b1111111110101111;
    assign weights1[62][713] = 16'b1111111110110011;
    assign weights1[62][714] = 16'b1111111110111000;
    assign weights1[62][715] = 16'b1111111110101011;
    assign weights1[62][716] = 16'b1111111111000011;
    assign weights1[62][717] = 16'b1111111110111101;
    assign weights1[62][718] = 16'b1111111111000100;
    assign weights1[62][719] = 16'b1111111111001011;
    assign weights1[62][720] = 16'b1111111110111111;
    assign weights1[62][721] = 16'b1111111111010010;
    assign weights1[62][722] = 16'b1111111111011010;
    assign weights1[62][723] = 16'b1111111111010011;
    assign weights1[62][724] = 16'b1111111111011010;
    assign weights1[62][725] = 16'b1111111111101100;
    assign weights1[62][726] = 16'b1111111111101011;
    assign weights1[62][727] = 16'b1111111111111000;
    assign weights1[62][728] = 16'b1111111111111101;
    assign weights1[62][729] = 16'b0000000000000000;
    assign weights1[62][730] = 16'b1111111111111000;
    assign weights1[62][731] = 16'b1111111111110110;
    assign weights1[62][732] = 16'b1111111111100101;
    assign weights1[62][733] = 16'b1111111111011100;
    assign weights1[62][734] = 16'b1111111111011110;
    assign weights1[62][735] = 16'b1111111111001000;
    assign weights1[62][736] = 16'b1111111111001011;
    assign weights1[62][737] = 16'b1111111111010001;
    assign weights1[62][738] = 16'b1111111111011000;
    assign weights1[62][739] = 16'b1111111111000101;
    assign weights1[62][740] = 16'b1111111111001100;
    assign weights1[62][741] = 16'b1111111111010101;
    assign weights1[62][742] = 16'b1111111111010111;
    assign weights1[62][743] = 16'b1111111111010110;
    assign weights1[62][744] = 16'b1111111111011001;
    assign weights1[62][745] = 16'b1111111111010111;
    assign weights1[62][746] = 16'b1111111111001110;
    assign weights1[62][747] = 16'b1111111111011110;
    assign weights1[62][748] = 16'b1111111111011010;
    assign weights1[62][749] = 16'b1111111111100000;
    assign weights1[62][750] = 16'b1111111111101101;
    assign weights1[62][751] = 16'b1111111111101001;
    assign weights1[62][752] = 16'b1111111111101101;
    assign weights1[62][753] = 16'b1111111111110001;
    assign weights1[62][754] = 16'b1111111111111001;
    assign weights1[62][755] = 16'b1111111111111100;
    assign weights1[62][756] = 16'b1111111111111111;
    assign weights1[62][757] = 16'b1111111111111101;
    assign weights1[62][758] = 16'b1111111111111010;
    assign weights1[62][759] = 16'b1111111111111100;
    assign weights1[62][760] = 16'b1111111111110111;
    assign weights1[62][761] = 16'b1111111111110101;
    assign weights1[62][762] = 16'b1111111111101111;
    assign weights1[62][763] = 16'b1111111111101010;
    assign weights1[62][764] = 16'b1111111111101011;
    assign weights1[62][765] = 16'b1111111111100110;
    assign weights1[62][766] = 16'b1111111111100111;
    assign weights1[62][767] = 16'b1111111111101000;
    assign weights1[62][768] = 16'b1111111111101010;
    assign weights1[62][769] = 16'b1111111111101011;
    assign weights1[62][770] = 16'b1111111111100011;
    assign weights1[62][771] = 16'b1111111111101000;
    assign weights1[62][772] = 16'b1111111111100100;
    assign weights1[62][773] = 16'b1111111111100100;
    assign weights1[62][774] = 16'b1111111111011110;
    assign weights1[62][775] = 16'b1111111111100000;
    assign weights1[62][776] = 16'b1111111111110000;
    assign weights1[62][777] = 16'b1111111111100111;
    assign weights1[62][778] = 16'b1111111111110110;
    assign weights1[62][779] = 16'b1111111111110010;
    assign weights1[62][780] = 16'b1111111111110010;
    assign weights1[62][781] = 16'b1111111111110100;
    assign weights1[62][782] = 16'b1111111111111011;
    assign weights1[62][783] = 16'b1111111111111101;
    assign weights1[63][0] = 16'b0000000000000001;
    assign weights1[63][1] = 16'b0000000000000000;
    assign weights1[63][2] = 16'b0000000000000001;
    assign weights1[63][3] = 16'b0000000000000100;
    assign weights1[63][4] = 16'b0000000000000111;
    assign weights1[63][5] = 16'b0000000000001001;
    assign weights1[63][6] = 16'b0000000000010000;
    assign weights1[63][7] = 16'b0000000000011010;
    assign weights1[63][8] = 16'b0000000000011110;
    assign weights1[63][9] = 16'b0000000000100001;
    assign weights1[63][10] = 16'b0000000000110010;
    assign weights1[63][11] = 16'b0000000000111010;
    assign weights1[63][12] = 16'b0000000000101110;
    assign weights1[63][13] = 16'b0000000000110001;
    assign weights1[63][14] = 16'b0000000000001110;
    assign weights1[63][15] = 16'b0000000000100111;
    assign weights1[63][16] = 16'b0000000000110100;
    assign weights1[63][17] = 16'b0000000000101000;
    assign weights1[63][18] = 16'b0000000000101011;
    assign weights1[63][19] = 16'b0000000000100110;
    assign weights1[63][20] = 16'b0000000000010111;
    assign weights1[63][21] = 16'b0000000000100010;
    assign weights1[63][22] = 16'b0000000000010100;
    assign weights1[63][23] = 16'b0000000000001100;
    assign weights1[63][24] = 16'b0000000000001011;
    assign weights1[63][25] = 16'b0000000000000000;
    assign weights1[63][26] = 16'b0000000000001000;
    assign weights1[63][27] = 16'b0000000000000010;
    assign weights1[63][28] = 16'b0000000000000001;
    assign weights1[63][29] = 16'b1111111111111111;
    assign weights1[63][30] = 16'b0000000000000101;
    assign weights1[63][31] = 16'b0000000000000110;
    assign weights1[63][32] = 16'b0000000000001010;
    assign weights1[63][33] = 16'b0000000000001011;
    assign weights1[63][34] = 16'b0000000000010001;
    assign weights1[63][35] = 16'b0000000000001110;
    assign weights1[63][36] = 16'b0000000000010011;
    assign weights1[63][37] = 16'b0000000000001001;
    assign weights1[63][38] = 16'b0000000000001100;
    assign weights1[63][39] = 16'b0000000000010011;
    assign weights1[63][40] = 16'b0000000000000111;
    assign weights1[63][41] = 16'b1111111111101001;
    assign weights1[63][42] = 16'b0000000000000101;
    assign weights1[63][43] = 16'b0000000000010111;
    assign weights1[63][44] = 16'b0000000000010111;
    assign weights1[63][45] = 16'b0000000000000001;
    assign weights1[63][46] = 16'b0000000000010010;
    assign weights1[63][47] = 16'b0000000000010000;
    assign weights1[63][48] = 16'b0000000000010010;
    assign weights1[63][49] = 16'b0000000000001011;
    assign weights1[63][50] = 16'b0000000000010111;
    assign weights1[63][51] = 16'b0000000000001001;
    assign weights1[63][52] = 16'b0000000000001111;
    assign weights1[63][53] = 16'b0000000000000110;
    assign weights1[63][54] = 16'b0000000000001011;
    assign weights1[63][55] = 16'b0000000000000100;
    assign weights1[63][56] = 16'b0000000000000001;
    assign weights1[63][57] = 16'b0000000000000011;
    assign weights1[63][58] = 16'b0000000000001010;
    assign weights1[63][59] = 16'b0000000000000010;
    assign weights1[63][60] = 16'b0000000000001010;
    assign weights1[63][61] = 16'b0000000000001010;
    assign weights1[63][62] = 16'b0000000000001001;
    assign weights1[63][63] = 16'b0000000000001011;
    assign weights1[63][64] = 16'b0000000000000000;
    assign weights1[63][65] = 16'b0000000000000001;
    assign weights1[63][66] = 16'b0000000000000101;
    assign weights1[63][67] = 16'b0000000000010000;
    assign weights1[63][68] = 16'b1111111111111011;
    assign weights1[63][69] = 16'b1111111111101111;
    assign weights1[63][70] = 16'b1111111111111001;
    assign weights1[63][71] = 16'b1111111111110110;
    assign weights1[63][72] = 16'b0000000000000000;
    assign weights1[63][73] = 16'b1111111111110110;
    assign weights1[63][74] = 16'b0000000000000101;
    assign weights1[63][75] = 16'b1111111111110100;
    assign weights1[63][76] = 16'b1111111111111101;
    assign weights1[63][77] = 16'b0000000000001001;
    assign weights1[63][78] = 16'b0000000000010101;
    assign weights1[63][79] = 16'b0000000000001010;
    assign weights1[63][80] = 16'b0000000000001011;
    assign weights1[63][81] = 16'b0000000000010011;
    assign weights1[63][82] = 16'b0000000000010001;
    assign weights1[63][83] = 16'b0000000000001000;
    assign weights1[63][84] = 16'b0000000000000010;
    assign weights1[63][85] = 16'b0000000000000001;
    assign weights1[63][86] = 16'b1111111111111110;
    assign weights1[63][87] = 16'b0000000000001101;
    assign weights1[63][88] = 16'b0000000000000110;
    assign weights1[63][89] = 16'b0000000000000110;
    assign weights1[63][90] = 16'b0000000000000000;
    assign weights1[63][91] = 16'b1111111111111100;
    assign weights1[63][92] = 16'b1111111111101101;
    assign weights1[63][93] = 16'b1111111111111000;
    assign weights1[63][94] = 16'b1111111111111001;
    assign weights1[63][95] = 16'b1111111111111011;
    assign weights1[63][96] = 16'b1111111111101101;
    assign weights1[63][97] = 16'b1111111111111101;
    assign weights1[63][98] = 16'b0000000000000011;
    assign weights1[63][99] = 16'b1111111111110001;
    assign weights1[63][100] = 16'b1111111111100100;
    assign weights1[63][101] = 16'b1111111111111010;
    assign weights1[63][102] = 16'b1111111111111111;
    assign weights1[63][103] = 16'b1111111111101101;
    assign weights1[63][104] = 16'b1111111111100110;
    assign weights1[63][105] = 16'b1111111111110011;
    assign weights1[63][106] = 16'b1111111111111000;
    assign weights1[63][107] = 16'b1111111111110110;
    assign weights1[63][108] = 16'b1111111111111101;
    assign weights1[63][109] = 16'b0000000000001111;
    assign weights1[63][110] = 16'b0000000000001010;
    assign weights1[63][111] = 16'b0000000000001001;
    assign weights1[63][112] = 16'b0000000000000000;
    assign weights1[63][113] = 16'b0000000000000011;
    assign weights1[63][114] = 16'b1111111111111110;
    assign weights1[63][115] = 16'b0000000000000011;
    assign weights1[63][116] = 16'b0000000000001100;
    assign weights1[63][117] = 16'b0000000000000011;
    assign weights1[63][118] = 16'b0000000000000011;
    assign weights1[63][119] = 16'b1111111111111010;
    assign weights1[63][120] = 16'b0000000000001100;
    assign weights1[63][121] = 16'b0000000000000101;
    assign weights1[63][122] = 16'b1111111111101101;
    assign weights1[63][123] = 16'b1111111111101101;
    assign weights1[63][124] = 16'b1111111111100010;
    assign weights1[63][125] = 16'b1111111111111101;
    assign weights1[63][126] = 16'b1111111111111000;
    assign weights1[63][127] = 16'b1111111111111101;
    assign weights1[63][128] = 16'b1111111111101000;
    assign weights1[63][129] = 16'b0000000000000000;
    assign weights1[63][130] = 16'b1111111111111110;
    assign weights1[63][131] = 16'b1111111111110011;
    assign weights1[63][132] = 16'b1111111111101100;
    assign weights1[63][133] = 16'b1111111111111001;
    assign weights1[63][134] = 16'b1111111111110100;
    assign weights1[63][135] = 16'b1111111111100000;
    assign weights1[63][136] = 16'b0000000000000001;
    assign weights1[63][137] = 16'b0000000000000000;
    assign weights1[63][138] = 16'b0000000000000010;
    assign weights1[63][139] = 16'b0000000000000010;
    assign weights1[63][140] = 16'b1111111111111111;
    assign weights1[63][141] = 16'b0000000000000011;
    assign weights1[63][142] = 16'b1111111111111110;
    assign weights1[63][143] = 16'b0000000000000110;
    assign weights1[63][144] = 16'b0000000000011000;
    assign weights1[63][145] = 16'b0000000000011001;
    assign weights1[63][146] = 16'b0000000000000000;
    assign weights1[63][147] = 16'b1111111111111011;
    assign weights1[63][148] = 16'b0000000000011010;
    assign weights1[63][149] = 16'b1111111111101101;
    assign weights1[63][150] = 16'b0000000000001010;
    assign weights1[63][151] = 16'b1111111111101111;
    assign weights1[63][152] = 16'b1111111111110000;
    assign weights1[63][153] = 16'b0000000000001001;
    assign weights1[63][154] = 16'b1111111111111110;
    assign weights1[63][155] = 16'b0000000000010010;
    assign weights1[63][156] = 16'b0000000000010010;
    assign weights1[63][157] = 16'b0000000000011000;
    assign weights1[63][158] = 16'b1111111111100111;
    assign weights1[63][159] = 16'b1111111111100011;
    assign weights1[63][160] = 16'b1111111111110010;
    assign weights1[63][161] = 16'b1111111111100011;
    assign weights1[63][162] = 16'b1111111111110101;
    assign weights1[63][163] = 16'b1111111111110111;
    assign weights1[63][164] = 16'b0000000000001100;
    assign weights1[63][165] = 16'b0000000000000000;
    assign weights1[63][166] = 16'b0000000000000000;
    assign weights1[63][167] = 16'b0000000000000011;
    assign weights1[63][168] = 16'b1111111111111110;
    assign weights1[63][169] = 16'b1111111111111111;
    assign weights1[63][170] = 16'b1111111111110111;
    assign weights1[63][171] = 16'b0000000000000001;
    assign weights1[63][172] = 16'b0000000000001001;
    assign weights1[63][173] = 16'b0000000000010110;
    assign weights1[63][174] = 16'b0000000000000011;
    assign weights1[63][175] = 16'b0000000000010000;
    assign weights1[63][176] = 16'b0000000000001100;
    assign weights1[63][177] = 16'b0000000000000001;
    assign weights1[63][178] = 16'b0000000000000101;
    assign weights1[63][179] = 16'b0000000000000110;
    assign weights1[63][180] = 16'b1111111111101111;
    assign weights1[63][181] = 16'b0000000000001100;
    assign weights1[63][182] = 16'b1111111111111001;
    assign weights1[63][183] = 16'b1111111111110010;
    assign weights1[63][184] = 16'b0000000000001010;
    assign weights1[63][185] = 16'b1111111111111110;
    assign weights1[63][186] = 16'b0000000000010101;
    assign weights1[63][187] = 16'b0000000000000001;
    assign weights1[63][188] = 16'b1111111111111001;
    assign weights1[63][189] = 16'b0000000000000100;
    assign weights1[63][190] = 16'b0000000000000110;
    assign weights1[63][191] = 16'b1111111111011011;
    assign weights1[63][192] = 16'b0000000000001100;
    assign weights1[63][193] = 16'b0000000000000100;
    assign weights1[63][194] = 16'b0000000000001010;
    assign weights1[63][195] = 16'b0000000000000000;
    assign weights1[63][196] = 16'b1111111111111100;
    assign weights1[63][197] = 16'b1111111111111001;
    assign weights1[63][198] = 16'b1111111111110100;
    assign weights1[63][199] = 16'b0000000000001110;
    assign weights1[63][200] = 16'b0000000000001010;
    assign weights1[63][201] = 16'b1111111111111101;
    assign weights1[63][202] = 16'b0000000000000011;
    assign weights1[63][203] = 16'b0000000000011111;
    assign weights1[63][204] = 16'b1111111111111110;
    assign weights1[63][205] = 16'b1111111111100101;
    assign weights1[63][206] = 16'b0000000000001111;
    assign weights1[63][207] = 16'b1111111111111000;
    assign weights1[63][208] = 16'b0000000000001111;
    assign weights1[63][209] = 16'b0000000000010111;
    assign weights1[63][210] = 16'b0000000000000110;
    assign weights1[63][211] = 16'b0000000000001011;
    assign weights1[63][212] = 16'b0000000000000011;
    assign weights1[63][213] = 16'b1111111111110111;
    assign weights1[63][214] = 16'b1111111111101110;
    assign weights1[63][215] = 16'b1111111111111011;
    assign weights1[63][216] = 16'b0000000000000100;
    assign weights1[63][217] = 16'b0000000000001011;
    assign weights1[63][218] = 16'b0000000000001011;
    assign weights1[63][219] = 16'b0000000000001011;
    assign weights1[63][220] = 16'b0000000000001111;
    assign weights1[63][221] = 16'b0000000000010001;
    assign weights1[63][222] = 16'b0000000000000011;
    assign weights1[63][223] = 16'b1111111111111100;
    assign weights1[63][224] = 16'b0000000000000100;
    assign weights1[63][225] = 16'b1111111111111000;
    assign weights1[63][226] = 16'b0000000000001010;
    assign weights1[63][227] = 16'b0000000000000010;
    assign weights1[63][228] = 16'b0000000000001111;
    assign weights1[63][229] = 16'b0000000000010101;
    assign weights1[63][230] = 16'b0000000000010111;
    assign weights1[63][231] = 16'b0000000000011111;
    assign weights1[63][232] = 16'b0000000000011101;
    assign weights1[63][233] = 16'b0000000000000010;
    assign weights1[63][234] = 16'b0000000000011000;
    assign weights1[63][235] = 16'b0000000000001110;
    assign weights1[63][236] = 16'b1111111111100111;
    assign weights1[63][237] = 16'b1111111111110100;
    assign weights1[63][238] = 16'b1111111111110111;
    assign weights1[63][239] = 16'b0000000000011110;
    assign weights1[63][240] = 16'b0000000000000000;
    assign weights1[63][241] = 16'b0000000000001001;
    assign weights1[63][242] = 16'b1111111111111100;
    assign weights1[63][243] = 16'b0000000000000001;
    assign weights1[63][244] = 16'b0000000000010111;
    assign weights1[63][245] = 16'b0000000000010100;
    assign weights1[63][246] = 16'b0000000000010010;
    assign weights1[63][247] = 16'b0000000000001101;
    assign weights1[63][248] = 16'b0000000000001110;
    assign weights1[63][249] = 16'b0000000000001110;
    assign weights1[63][250] = 16'b1111111111111111;
    assign weights1[63][251] = 16'b0000000000000010;
    assign weights1[63][252] = 16'b1111111111111110;
    assign weights1[63][253] = 16'b0000000000001000;
    assign weights1[63][254] = 16'b0000000000000010;
    assign weights1[63][255] = 16'b0000000000000000;
    assign weights1[63][256] = 16'b0000000000010111;
    assign weights1[63][257] = 16'b0000000000000110;
    assign weights1[63][258] = 16'b1111111111111111;
    assign weights1[63][259] = 16'b0000000000011101;
    assign weights1[63][260] = 16'b0000000000101001;
    assign weights1[63][261] = 16'b0000000000001100;
    assign weights1[63][262] = 16'b0000000000001011;
    assign weights1[63][263] = 16'b0000000000010111;
    assign weights1[63][264] = 16'b0000000000000000;
    assign weights1[63][265] = 16'b0000000000000110;
    assign weights1[63][266] = 16'b0000000000010111;
    assign weights1[63][267] = 16'b1111111111101011;
    assign weights1[63][268] = 16'b0000000000001111;
    assign weights1[63][269] = 16'b0000000000001000;
    assign weights1[63][270] = 16'b0000000000010001;
    assign weights1[63][271] = 16'b0000000000000100;
    assign weights1[63][272] = 16'b0000000000011000;
    assign weights1[63][273] = 16'b0000000000000100;
    assign weights1[63][274] = 16'b1111111111111010;
    assign weights1[63][275] = 16'b0000000000001100;
    assign weights1[63][276] = 16'b0000000000010011;
    assign weights1[63][277] = 16'b0000000000001100;
    assign weights1[63][278] = 16'b0000000000011000;
    assign weights1[63][279] = 16'b0000000000010001;
    assign weights1[63][280] = 16'b1111111111111111;
    assign weights1[63][281] = 16'b0000000000001001;
    assign weights1[63][282] = 16'b0000000000010101;
    assign weights1[63][283] = 16'b0000000000010011;
    assign weights1[63][284] = 16'b0000000000010110;
    assign weights1[63][285] = 16'b0000000000010001;
    assign weights1[63][286] = 16'b0000000000000101;
    assign weights1[63][287] = 16'b0000000000010001;
    assign weights1[63][288] = 16'b0000000000011110;
    assign weights1[63][289] = 16'b0000000000001111;
    assign weights1[63][290] = 16'b0000000000100100;
    assign weights1[63][291] = 16'b0000000000001011;
    assign weights1[63][292] = 16'b1111111111111001;
    assign weights1[63][293] = 16'b0000000000010111;
    assign weights1[63][294] = 16'b0000000000011001;
    assign weights1[63][295] = 16'b0000000000011101;
    assign weights1[63][296] = 16'b0000000000010111;
    assign weights1[63][297] = 16'b0000000000010001;
    assign weights1[63][298] = 16'b0000000000000000;
    assign weights1[63][299] = 16'b0000000000011011;
    assign weights1[63][300] = 16'b0000000000010111;
    assign weights1[63][301] = 16'b0000000000011011;
    assign weights1[63][302] = 16'b0000000000001110;
    assign weights1[63][303] = 16'b0000000000001101;
    assign weights1[63][304] = 16'b0000000000001010;
    assign weights1[63][305] = 16'b0000000000011111;
    assign weights1[63][306] = 16'b0000000000001101;
    assign weights1[63][307] = 16'b0000000000001010;
    assign weights1[63][308] = 16'b0000000000000000;
    assign weights1[63][309] = 16'b0000000000001100;
    assign weights1[63][310] = 16'b0000000000011100;
    assign weights1[63][311] = 16'b0000000000010011;
    assign weights1[63][312] = 16'b1111111111111101;
    assign weights1[63][313] = 16'b0000000000001010;
    assign weights1[63][314] = 16'b0000000000011100;
    assign weights1[63][315] = 16'b0000000000010110;
    assign weights1[63][316] = 16'b0000000000101010;
    assign weights1[63][317] = 16'b0000000000010011;
    assign weights1[63][318] = 16'b0000000000100100;
    assign weights1[63][319] = 16'b0000000000101110;
    assign weights1[63][320] = 16'b0000000000100111;
    assign weights1[63][321] = 16'b0000000000100001;
    assign weights1[63][322] = 16'b0000000000011110;
    assign weights1[63][323] = 16'b0000000000010101;
    assign weights1[63][324] = 16'b0000000000101001;
    assign weights1[63][325] = 16'b0000000000100110;
    assign weights1[63][326] = 16'b0000000000100010;
    assign weights1[63][327] = 16'b0000000000001110;
    assign weights1[63][328] = 16'b0000000000101011;
    assign weights1[63][329] = 16'b0000000000010101;
    assign weights1[63][330] = 16'b0000000000010101;
    assign weights1[63][331] = 16'b0000000000101011;
    assign weights1[63][332] = 16'b0000000000000110;
    assign weights1[63][333] = 16'b0000000000010110;
    assign weights1[63][334] = 16'b0000000000001110;
    assign weights1[63][335] = 16'b0000000000000110;
    assign weights1[63][336] = 16'b1111111111111111;
    assign weights1[63][337] = 16'b0000000000000110;
    assign weights1[63][338] = 16'b0000000000010111;
    assign weights1[63][339] = 16'b0000000000011010;
    assign weights1[63][340] = 16'b0000000000010111;
    assign weights1[63][341] = 16'b1111111111110100;
    assign weights1[63][342] = 16'b0000000000010011;
    assign weights1[63][343] = 16'b0000000000010101;
    assign weights1[63][344] = 16'b1111111111111001;
    assign weights1[63][345] = 16'b0000000000100101;
    assign weights1[63][346] = 16'b0000000000100010;
    assign weights1[63][347] = 16'b0000000000100011;
    assign weights1[63][348] = 16'b0000000000100110;
    assign weights1[63][349] = 16'b0000000000011101;
    assign weights1[63][350] = 16'b0000000000011010;
    assign weights1[63][351] = 16'b0000000000011100;
    assign weights1[63][352] = 16'b0000000000100101;
    assign weights1[63][353] = 16'b0000000000011101;
    assign weights1[63][354] = 16'b0000000000100001;
    assign weights1[63][355] = 16'b0000000000101000;
    assign weights1[63][356] = 16'b0000000000011001;
    assign weights1[63][357] = 16'b0000000000101100;
    assign weights1[63][358] = 16'b0000000000001001;
    assign weights1[63][359] = 16'b0000000000101010;
    assign weights1[63][360] = 16'b0000000000100100;
    assign weights1[63][361] = 16'b0000000000100100;
    assign weights1[63][362] = 16'b0000000000010010;
    assign weights1[63][363] = 16'b0000000000001110;
    assign weights1[63][364] = 16'b1111111111111110;
    assign weights1[63][365] = 16'b0000000000001000;
    assign weights1[63][366] = 16'b0000000000010010;
    assign weights1[63][367] = 16'b0000000000100110;
    assign weights1[63][368] = 16'b0000000000011110;
    assign weights1[63][369] = 16'b0000000000001101;
    assign weights1[63][370] = 16'b0000000000001010;
    assign weights1[63][371] = 16'b0000000000001011;
    assign weights1[63][372] = 16'b0000000000001100;
    assign weights1[63][373] = 16'b0000000000001000;
    assign weights1[63][374] = 16'b0000000000011100;
    assign weights1[63][375] = 16'b0000000000100110;
    assign weights1[63][376] = 16'b0000000000110010;
    assign weights1[63][377] = 16'b0000000000100010;
    assign weights1[63][378] = 16'b0000000000011011;
    assign weights1[63][379] = 16'b0000000000010001;
    assign weights1[63][380] = 16'b0000000000100110;
    assign weights1[63][381] = 16'b0000000000101000;
    assign weights1[63][382] = 16'b0000000000001001;
    assign weights1[63][383] = 16'b0000000000101000;
    assign weights1[63][384] = 16'b0000000000100000;
    assign weights1[63][385] = 16'b0000000000010010;
    assign weights1[63][386] = 16'b0000000000011110;
    assign weights1[63][387] = 16'b0000000000100000;
    assign weights1[63][388] = 16'b0000000000100110;
    assign weights1[63][389] = 16'b0000000000010001;
    assign weights1[63][390] = 16'b0000000000010001;
    assign weights1[63][391] = 16'b1111111111111111;
    assign weights1[63][392] = 16'b1111111111111011;
    assign weights1[63][393] = 16'b0000000000000000;
    assign weights1[63][394] = 16'b0000000000001010;
    assign weights1[63][395] = 16'b1111111111111010;
    assign weights1[63][396] = 16'b1111111111111000;
    assign weights1[63][397] = 16'b0000000000011001;
    assign weights1[63][398] = 16'b0000000000001000;
    assign weights1[63][399] = 16'b0000000000011011;
    assign weights1[63][400] = 16'b0000000000100011;
    assign weights1[63][401] = 16'b0000000000100000;
    assign weights1[63][402] = 16'b0000000000100110;
    assign weights1[63][403] = 16'b0000000000110011;
    assign weights1[63][404] = 16'b0000000000101100;
    assign weights1[63][405] = 16'b0000000000100001;
    assign weights1[63][406] = 16'b0000000000100101;
    assign weights1[63][407] = 16'b0000000000110010;
    assign weights1[63][408] = 16'b0000000000011010;
    assign weights1[63][409] = 16'b0000000000011111;
    assign weights1[63][410] = 16'b0000000000010010;
    assign weights1[63][411] = 16'b0000000000010000;
    assign weights1[63][412] = 16'b0000000000100001;
    assign weights1[63][413] = 16'b0000000000100110;
    assign weights1[63][414] = 16'b0000000000101110;
    assign weights1[63][415] = 16'b0000000000001111;
    assign weights1[63][416] = 16'b0000000000000111;
    assign weights1[63][417] = 16'b1111111111111011;
    assign weights1[63][418] = 16'b0000000000000101;
    assign weights1[63][419] = 16'b0000000000000110;
    assign weights1[63][420] = 16'b1111111111111110;
    assign weights1[63][421] = 16'b1111111111101111;
    assign weights1[63][422] = 16'b1111111111100110;
    assign weights1[63][423] = 16'b1111111111100010;
    assign weights1[63][424] = 16'b1111111111101110;
    assign weights1[63][425] = 16'b1111111111110001;
    assign weights1[63][426] = 16'b1111111111101001;
    assign weights1[63][427] = 16'b0000000000000010;
    assign weights1[63][428] = 16'b1111111111110110;
    assign weights1[63][429] = 16'b1111111111111101;
    assign weights1[63][430] = 16'b0000000000001000;
    assign weights1[63][431] = 16'b0000000000010111;
    assign weights1[63][432] = 16'b0000000000101100;
    assign weights1[63][433] = 16'b0000000000111000;
    assign weights1[63][434] = 16'b0000000000111110;
    assign weights1[63][435] = 16'b0000000000101110;
    assign weights1[63][436] = 16'b0000000000101110;
    assign weights1[63][437] = 16'b0000000000100110;
    assign weights1[63][438] = 16'b0000000000110011;
    assign weights1[63][439] = 16'b0000000000101000;
    assign weights1[63][440] = 16'b0000000000010100;
    assign weights1[63][441] = 16'b0000000000001100;
    assign weights1[63][442] = 16'b0000000000000010;
    assign weights1[63][443] = 16'b0000000000010010;
    assign weights1[63][444] = 16'b0000000000001001;
    assign weights1[63][445] = 16'b0000000000000001;
    assign weights1[63][446] = 16'b0000000000000100;
    assign weights1[63][447] = 16'b0000000000001100;
    assign weights1[63][448] = 16'b1111111111110001;
    assign weights1[63][449] = 16'b1111111111100100;
    assign weights1[63][450] = 16'b1111111111101011;
    assign weights1[63][451] = 16'b1111111111011000;
    assign weights1[63][452] = 16'b1111111111011111;
    assign weights1[63][453] = 16'b1111111111001010;
    assign weights1[63][454] = 16'b1111111111101110;
    assign weights1[63][455] = 16'b1111111111111001;
    assign weights1[63][456] = 16'b1111111111011100;
    assign weights1[63][457] = 16'b1111111111101000;
    assign weights1[63][458] = 16'b1111111111101100;
    assign weights1[63][459] = 16'b1111111111100010;
    assign weights1[63][460] = 16'b0000000000000111;
    assign weights1[63][461] = 16'b0000000000001000;
    assign weights1[63][462] = 16'b0000000000110010;
    assign weights1[63][463] = 16'b0000000000010001;
    assign weights1[63][464] = 16'b0000000000011111;
    assign weights1[63][465] = 16'b0000000000010000;
    assign weights1[63][466] = 16'b0000000000010110;
    assign weights1[63][467] = 16'b1111111111110000;
    assign weights1[63][468] = 16'b1111111111100110;
    assign weights1[63][469] = 16'b1111111111111101;
    assign weights1[63][470] = 16'b1111111111011000;
    assign weights1[63][471] = 16'b1111111111101011;
    assign weights1[63][472] = 16'b1111111111111100;
    assign weights1[63][473] = 16'b1111111111111000;
    assign weights1[63][474] = 16'b1111111111111011;
    assign weights1[63][475] = 16'b1111111111111101;
    assign weights1[63][476] = 16'b1111111111101100;
    assign weights1[63][477] = 16'b1111111111011111;
    assign weights1[63][478] = 16'b1111111111001110;
    assign weights1[63][479] = 16'b1111111111001101;
    assign weights1[63][480] = 16'b1111111111001101;
    assign weights1[63][481] = 16'b1111111111010101;
    assign weights1[63][482] = 16'b1111111111011111;
    assign weights1[63][483] = 16'b1111111111000110;
    assign weights1[63][484] = 16'b1111111110111011;
    assign weights1[63][485] = 16'b1111111110110010;
    assign weights1[63][486] = 16'b1111111110101110;
    assign weights1[63][487] = 16'b1111111110101000;
    assign weights1[63][488] = 16'b1111111110110000;
    assign weights1[63][489] = 16'b1111111110110111;
    assign weights1[63][490] = 16'b1111111111001111;
    assign weights1[63][491] = 16'b1111111111010011;
    assign weights1[63][492] = 16'b1111111111011010;
    assign weights1[63][493] = 16'b1111111111100011;
    assign weights1[63][494] = 16'b1111111111001110;
    assign weights1[63][495] = 16'b1111111111010101;
    assign weights1[63][496] = 16'b1111111111001101;
    assign weights1[63][497] = 16'b1111111111010110;
    assign weights1[63][498] = 16'b1111111111000110;
    assign weights1[63][499] = 16'b1111111111001100;
    assign weights1[63][500] = 16'b1111111111001011;
    assign weights1[63][501] = 16'b1111111111011110;
    assign weights1[63][502] = 16'b1111111111100111;
    assign weights1[63][503] = 16'b1111111111111011;
    assign weights1[63][504] = 16'b1111111111101111;
    assign weights1[63][505] = 16'b1111111111011111;
    assign weights1[63][506] = 16'b1111111111010110;
    assign weights1[63][507] = 16'b1111111111011110;
    assign weights1[63][508] = 16'b1111111111010101;
    assign weights1[63][509] = 16'b1111111111010000;
    assign weights1[63][510] = 16'b1111111111001001;
    assign weights1[63][511] = 16'b1111111111010001;
    assign weights1[63][512] = 16'b1111111111011100;
    assign weights1[63][513] = 16'b1111111111010101;
    assign weights1[63][514] = 16'b1111111111000010;
    assign weights1[63][515] = 16'b1111111110101111;
    assign weights1[63][516] = 16'b1111111110011001;
    assign weights1[63][517] = 16'b1111111110010111;
    assign weights1[63][518] = 16'b1111111101111000;
    assign weights1[63][519] = 16'b1111111110100011;
    assign weights1[63][520] = 16'b1111111110100100;
    assign weights1[63][521] = 16'b1111111110100111;
    assign weights1[63][522] = 16'b1111111111000011;
    assign weights1[63][523] = 16'b1111111111011000;
    assign weights1[63][524] = 16'b1111111110110101;
    assign weights1[63][525] = 16'b1111111111011010;
    assign weights1[63][526] = 16'b1111111110110010;
    assign weights1[63][527] = 16'b1111111110111011;
    assign weights1[63][528] = 16'b1111111110110010;
    assign weights1[63][529] = 16'b1111111111001111;
    assign weights1[63][530] = 16'b1111111111100101;
    assign weights1[63][531] = 16'b1111111111110000;
    assign weights1[63][532] = 16'b1111111111101111;
    assign weights1[63][533] = 16'b1111111111100110;
    assign weights1[63][534] = 16'b1111111111100011;
    assign weights1[63][535] = 16'b1111111111100110;
    assign weights1[63][536] = 16'b1111111111100101;
    assign weights1[63][537] = 16'b1111111111100101;
    assign weights1[63][538] = 16'b1111111111011101;
    assign weights1[63][539] = 16'b1111111111010100;
    assign weights1[63][540] = 16'b1111111111011001;
    assign weights1[63][541] = 16'b1111111111010111;
    assign weights1[63][542] = 16'b1111111111001000;
    assign weights1[63][543] = 16'b1111111111010001;
    assign weights1[63][544] = 16'b1111111110111011;
    assign weights1[63][545] = 16'b1111111110111111;
    assign weights1[63][546] = 16'b1111111111001101;
    assign weights1[63][547] = 16'b1111111110111000;
    assign weights1[63][548] = 16'b1111111111000011;
    assign weights1[63][549] = 16'b1111111110111011;
    assign weights1[63][550] = 16'b1111111111000100;
    assign weights1[63][551] = 16'b1111111111001000;
    assign weights1[63][552] = 16'b1111111111001010;
    assign weights1[63][553] = 16'b1111111111010000;
    assign weights1[63][554] = 16'b1111111110101110;
    assign weights1[63][555] = 16'b1111111111000011;
    assign weights1[63][556] = 16'b1111111111000001;
    assign weights1[63][557] = 16'b1111111111010011;
    assign weights1[63][558] = 16'b1111111111011100;
    assign weights1[63][559] = 16'b1111111111110010;
    assign weights1[63][560] = 16'b1111111111110111;
    assign weights1[63][561] = 16'b1111111111101011;
    assign weights1[63][562] = 16'b1111111111100110;
    assign weights1[63][563] = 16'b1111111111101110;
    assign weights1[63][564] = 16'b1111111111100101;
    assign weights1[63][565] = 16'b0000000000000000;
    assign weights1[63][566] = 16'b1111111111110011;
    assign weights1[63][567] = 16'b1111111111011110;
    assign weights1[63][568] = 16'b1111111111010110;
    assign weights1[63][569] = 16'b1111111111010100;
    assign weights1[63][570] = 16'b1111111111011110;
    assign weights1[63][571] = 16'b1111111110111011;
    assign weights1[63][572] = 16'b1111111111000110;
    assign weights1[63][573] = 16'b1111111110111000;
    assign weights1[63][574] = 16'b1111111111001101;
    assign weights1[63][575] = 16'b1111111111000101;
    assign weights1[63][576] = 16'b1111111111010010;
    assign weights1[63][577] = 16'b1111111111000111;
    assign weights1[63][578] = 16'b1111111111010001;
    assign weights1[63][579] = 16'b1111111111010001;
    assign weights1[63][580] = 16'b1111111110111001;
    assign weights1[63][581] = 16'b1111111111001010;
    assign weights1[63][582] = 16'b1111111111001000;
    assign weights1[63][583] = 16'b1111111111010000;
    assign weights1[63][584] = 16'b1111111111010111;
    assign weights1[63][585] = 16'b1111111111011011;
    assign weights1[63][586] = 16'b1111111111100111;
    assign weights1[63][587] = 16'b1111111111111000;
    assign weights1[63][588] = 16'b1111111111111000;
    assign weights1[63][589] = 16'b1111111111111101;
    assign weights1[63][590] = 16'b1111111111110011;
    assign weights1[63][591] = 16'b1111111111111010;
    assign weights1[63][592] = 16'b1111111111111011;
    assign weights1[63][593] = 16'b1111111111101011;
    assign weights1[63][594] = 16'b1111111111101101;
    assign weights1[63][595] = 16'b1111111111010110;
    assign weights1[63][596] = 16'b1111111111011001;
    assign weights1[63][597] = 16'b1111111111011110;
    assign weights1[63][598] = 16'b1111111111110000;
    assign weights1[63][599] = 16'b1111111111010000;
    assign weights1[63][600] = 16'b1111111111000001;
    assign weights1[63][601] = 16'b1111111111000001;
    assign weights1[63][602] = 16'b1111111111001111;
    assign weights1[63][603] = 16'b1111111111001110;
    assign weights1[63][604] = 16'b1111111110111100;
    assign weights1[63][605] = 16'b1111111111000010;
    assign weights1[63][606] = 16'b1111111111001111;
    assign weights1[63][607] = 16'b1111111111010110;
    assign weights1[63][608] = 16'b1111111111001110;
    assign weights1[63][609] = 16'b1111111111011100;
    assign weights1[63][610] = 16'b1111111111011001;
    assign weights1[63][611] = 16'b1111111111011100;
    assign weights1[63][612] = 16'b1111111111100010;
    assign weights1[63][613] = 16'b1111111111011110;
    assign weights1[63][614] = 16'b1111111111101011;
    assign weights1[63][615] = 16'b1111111111110110;
    assign weights1[63][616] = 16'b1111111111111011;
    assign weights1[63][617] = 16'b1111111111111110;
    assign weights1[63][618] = 16'b1111111111110101;
    assign weights1[63][619] = 16'b1111111111111011;
    assign weights1[63][620] = 16'b1111111111110101;
    assign weights1[63][621] = 16'b1111111111110000;
    assign weights1[63][622] = 16'b1111111111101000;
    assign weights1[63][623] = 16'b1111111111100001;
    assign weights1[63][624] = 16'b1111111111111010;
    assign weights1[63][625] = 16'b1111111111011101;
    assign weights1[63][626] = 16'b1111111111101001;
    assign weights1[63][627] = 16'b1111111111100010;
    assign weights1[63][628] = 16'b1111111111000110;
    assign weights1[63][629] = 16'b1111111111101010;
    assign weights1[63][630] = 16'b1111111111011111;
    assign weights1[63][631] = 16'b1111111111011101;
    assign weights1[63][632] = 16'b1111111111011100;
    assign weights1[63][633] = 16'b1111111111010010;
    assign weights1[63][634] = 16'b1111111111100011;
    assign weights1[63][635] = 16'b1111111111010111;
    assign weights1[63][636] = 16'b1111111111100001;
    assign weights1[63][637] = 16'b1111111111110100;
    assign weights1[63][638] = 16'b1111111111101010;
    assign weights1[63][639] = 16'b1111111111010101;
    assign weights1[63][640] = 16'b1111111111101010;
    assign weights1[63][641] = 16'b1111111111101000;
    assign weights1[63][642] = 16'b1111111111110010;
    assign weights1[63][643] = 16'b1111111111110111;
    assign weights1[63][644] = 16'b1111111111111111;
    assign weights1[63][645] = 16'b1111111111111110;
    assign weights1[63][646] = 16'b1111111111110110;
    assign weights1[63][647] = 16'b1111111111111001;
    assign weights1[63][648] = 16'b1111111111101110;
    assign weights1[63][649] = 16'b1111111111100011;
    assign weights1[63][650] = 16'b1111111111110111;
    assign weights1[63][651] = 16'b1111111111011011;
    assign weights1[63][652] = 16'b1111111111011101;
    assign weights1[63][653] = 16'b1111111111101100;
    assign weights1[63][654] = 16'b1111111111101000;
    assign weights1[63][655] = 16'b1111111111101100;
    assign weights1[63][656] = 16'b0000000000001010;
    assign weights1[63][657] = 16'b1111111111110001;
    assign weights1[63][658] = 16'b1111111111011000;
    assign weights1[63][659] = 16'b1111111111010001;
    assign weights1[63][660] = 16'b0000000000000011;
    assign weights1[63][661] = 16'b1111111111101001;
    assign weights1[63][662] = 16'b1111111111011111;
    assign weights1[63][663] = 16'b1111111111111010;
    assign weights1[63][664] = 16'b1111111111011111;
    assign weights1[63][665] = 16'b1111111111101011;
    assign weights1[63][666] = 16'b1111111111101110;
    assign weights1[63][667] = 16'b1111111111101001;
    assign weights1[63][668] = 16'b1111111111101111;
    assign weights1[63][669] = 16'b1111111111110100;
    assign weights1[63][670] = 16'b1111111111110111;
    assign weights1[63][671] = 16'b1111111111111001;
    assign weights1[63][672] = 16'b1111111111111110;
    assign weights1[63][673] = 16'b1111111111111001;
    assign weights1[63][674] = 16'b1111111111110010;
    assign weights1[63][675] = 16'b1111111111110111;
    assign weights1[63][676] = 16'b1111111111110111;
    assign weights1[63][677] = 16'b1111111111100111;
    assign weights1[63][678] = 16'b1111111111101100;
    assign weights1[63][679] = 16'b1111111111001110;
    assign weights1[63][680] = 16'b1111111111010011;
    assign weights1[63][681] = 16'b1111111111100110;
    assign weights1[63][682] = 16'b1111111111101000;
    assign weights1[63][683] = 16'b1111111111110010;
    assign weights1[63][684] = 16'b1111111111111000;
    assign weights1[63][685] = 16'b1111111111101001;
    assign weights1[63][686] = 16'b1111111111100111;
    assign weights1[63][687] = 16'b1111111111011101;
    assign weights1[63][688] = 16'b1111111111101110;
    assign weights1[63][689] = 16'b1111111111011000;
    assign weights1[63][690] = 16'b1111111111101101;
    assign weights1[63][691] = 16'b1111111111100001;
    assign weights1[63][692] = 16'b0000000000000111;
    assign weights1[63][693] = 16'b1111111111110110;
    assign weights1[63][694] = 16'b1111111111110001;
    assign weights1[63][695] = 16'b1111111111101100;
    assign weights1[63][696] = 16'b1111111111110001;
    assign weights1[63][697] = 16'b1111111111111001;
    assign weights1[63][698] = 16'b0000000000000010;
    assign weights1[63][699] = 16'b1111111111111110;
    assign weights1[63][700] = 16'b1111111111111110;
    assign weights1[63][701] = 16'b1111111111111000;
    assign weights1[63][702] = 16'b1111111111111001;
    assign weights1[63][703] = 16'b1111111111110110;
    assign weights1[63][704] = 16'b1111111111111001;
    assign weights1[63][705] = 16'b1111111111101101;
    assign weights1[63][706] = 16'b1111111111010011;
    assign weights1[63][707] = 16'b1111111111001000;
    assign weights1[63][708] = 16'b1111111111010100;
    assign weights1[63][709] = 16'b1111111111100101;
    assign weights1[63][710] = 16'b1111111111001110;
    assign weights1[63][711] = 16'b1111111111000110;
    assign weights1[63][712] = 16'b1111111110011001;
    assign weights1[63][713] = 16'b1111111111001111;
    assign weights1[63][714] = 16'b1111111110111110;
    assign weights1[63][715] = 16'b1111111111100000;
    assign weights1[63][716] = 16'b1111111111000010;
    assign weights1[63][717] = 16'b1111111111000110;
    assign weights1[63][718] = 16'b1111111110101110;
    assign weights1[63][719] = 16'b1111111110101101;
    assign weights1[63][720] = 16'b1111111111001101;
    assign weights1[63][721] = 16'b1111111111010011;
    assign weights1[63][722] = 16'b1111111111101011;
    assign weights1[63][723] = 16'b1111111111110100;
    assign weights1[63][724] = 16'b1111111111110110;
    assign weights1[63][725] = 16'b1111111111111110;
    assign weights1[63][726] = 16'b0000000000000000;
    assign weights1[63][727] = 16'b0000000000000000;
    assign weights1[63][728] = 16'b1111111111111111;
    assign weights1[63][729] = 16'b1111111111111011;
    assign weights1[63][730] = 16'b1111111111111110;
    assign weights1[63][731] = 16'b1111111111111010;
    assign weights1[63][732] = 16'b1111111111111011;
    assign weights1[63][733] = 16'b1111111111111010;
    assign weights1[63][734] = 16'b1111111111110000;
    assign weights1[63][735] = 16'b1111111111100001;
    assign weights1[63][736] = 16'b1111111111001101;
    assign weights1[63][737] = 16'b1111111111001001;
    assign weights1[63][738] = 16'b1111111111010110;
    assign weights1[63][739] = 16'b1111111111001111;
    assign weights1[63][740] = 16'b1111111111010011;
    assign weights1[63][741] = 16'b1111111110111001;
    assign weights1[63][742] = 16'b1111111111001011;
    assign weights1[63][743] = 16'b1111111111010001;
    assign weights1[63][744] = 16'b1111111111000001;
    assign weights1[63][745] = 16'b1111111110111101;
    assign weights1[63][746] = 16'b1111111111001011;
    assign weights1[63][747] = 16'b1111111111000011;
    assign weights1[63][748] = 16'b1111111111010100;
    assign weights1[63][749] = 16'b1111111111011011;
    assign weights1[63][750] = 16'b1111111111100101;
    assign weights1[63][751] = 16'b1111111111110100;
    assign weights1[63][752] = 16'b1111111111111001;
    assign weights1[63][753] = 16'b1111111111111111;
    assign weights1[63][754] = 16'b0000000000000000;
    assign weights1[63][755] = 16'b0000000000000010;
    assign weights1[63][756] = 16'b0000000000000000;
    assign weights1[63][757] = 16'b1111111111111110;
    assign weights1[63][758] = 16'b0000000000000000;
    assign weights1[63][759] = 16'b0000000000000000;
    assign weights1[63][760] = 16'b1111111111111100;
    assign weights1[63][761] = 16'b1111111111111101;
    assign weights1[63][762] = 16'b1111111111111100;
    assign weights1[63][763] = 16'b1111111111110101;
    assign weights1[63][764] = 16'b1111111111101111;
    assign weights1[63][765] = 16'b1111111111100111;
    assign weights1[63][766] = 16'b1111111111100000;
    assign weights1[63][767] = 16'b1111111111101100;
    assign weights1[63][768] = 16'b1111111111110100;
    assign weights1[63][769] = 16'b1111111111101010;
    assign weights1[63][770] = 16'b1111111111011100;
    assign weights1[63][771] = 16'b1111111111100110;
    assign weights1[63][772] = 16'b1111111111011111;
    assign weights1[63][773] = 16'b1111111111011011;
    assign weights1[63][774] = 16'b1111111111010111;
    assign weights1[63][775] = 16'b1111111111100011;
    assign weights1[63][776] = 16'b1111111111100001;
    assign weights1[63][777] = 16'b1111111111100010;
    assign weights1[63][778] = 16'b1111111111110001;
    assign weights1[63][779] = 16'b1111111111110011;
    assign weights1[63][780] = 16'b1111111111111000;
    assign weights1[63][781] = 16'b1111111111111101;
    assign weights1[63][782] = 16'b1111111111111111;
    assign weights1[63][783] = 16'b0000000000000010;
    assign biases1[0] = 16'b0000000001110011;
    assign biases1[1] = 16'b0000000000100101;
    assign biases1[2] = 16'b0000000001000000;
    assign biases1[3] = 16'b0000000001010010;
    assign biases1[4] = 16'b1111111111100000;
    assign biases1[5] = 16'b0000000001000110;
    assign biases1[6] = 16'b0000000000000000;
    assign biases1[7] = 16'b0000000001010000;
    assign biases1[8] = 16'b1111111101110101;
    assign biases1[9] = 16'b1111111110010110;
    assign biases1[10] = 16'b1111111111001111;
    assign biases1[11] = 16'b0000000000011100;
    assign biases1[12] = 16'b0000000001000100;
    assign biases1[13] = 16'b0000000000011010;
    assign biases1[14] = 16'b1111111111111001;
    assign biases1[15] = 16'b1111111110010111;
    assign biases1[16] = 16'b1111111110010011;
    assign biases1[17] = 16'b0000000100011101;
    assign biases1[18] = 16'b0000000000011001;
    assign biases1[19] = 16'b1111111111111010;
    assign biases1[20] = 16'b0000000001001100;
    assign biases1[21] = 16'b0000000100001110;
    assign biases1[22] = 16'b0000000001000101;
    assign biases1[23] = 16'b1111111110100000;
    assign biases1[24] = 16'b0000000001001101;
    assign biases1[25] = 16'b0000000000011000;
    assign biases1[26] = 16'b1111111111101101;
    assign biases1[27] = 16'b0000000001001010;
    assign biases1[28] = 16'b0000000010000110;
    assign biases1[29] = 16'b0000000010011001;
    assign biases1[30] = 16'b0000000000010111;
    assign biases1[31] = 16'b0000000000100101;
    assign biases1[32] = 16'b1111111111110100;
    assign biases1[33] = 16'b1111111111101000;
    assign biases1[34] = 16'b0000000010011111;
    assign biases1[35] = 16'b0000000000110111;
    assign biases1[36] = 16'b0000000000001001;
    assign biases1[37] = 16'b0000000000101001;
    assign biases1[38] = 16'b0000000000011000;
    assign biases1[39] = 16'b0000000010011101;
    assign biases1[40] = 16'b1111111001101000;
    assign biases1[41] = 16'b1111111101011000;
    assign biases1[42] = 16'b0000000010010111;
    assign biases1[43] = 16'b0000000000000001;
    assign biases1[44] = 16'b0000000000011001;
    assign biases1[45] = 16'b1111111110001111;
    assign biases1[46] = 16'b0000000001000110;
    assign biases1[47] = 16'b0000000000101110;
    assign biases1[48] = 16'b0000000000110100;
    assign biases1[49] = 16'b0000000100010011;
    assign biases1[50] = 16'b0000000010000101;
    assign biases1[51] = 16'b1111111111111000;
    assign biases1[52] = 16'b0000000010010001;
    assign biases1[53] = 16'b1111111111110110;
    assign biases1[54] = 16'b0000000000000000;
    assign biases1[55] = 16'b0000000000000010;
    assign biases1[56] = 16'b0000000001000000;
    assign biases1[57] = 16'b0000000001001100;
    assign biases1[58] = 16'b1111111110100001;
    assign biases1[59] = 16'b0000000010010101;
    assign biases1[60] = 16'b1111111111100010;
    assign biases1[61] = 16'b0000000010100000;
    assign biases1[62] = 16'b0000000000001000;
    assign biases1[63] = 16'b1111111111101010;
    assign weights2[0][0] = 16'b0000000000000001;
    assign weights2[0][1] = 16'b1111111101101100;
    assign weights2[0][2] = 16'b0000000000000100;
    assign weights2[0][3] = 16'b1111111111001101;
    assign weights2[0][4] = 16'b0000000000001001;
    assign weights2[0][5] = 16'b1111111111110101;
    assign weights2[0][6] = 16'b0000000000000000;
    assign weights2[0][7] = 16'b1111111111110101;
    assign weights2[0][8] = 16'b0000000000100011;
    assign weights2[0][9] = 16'b0000000000010001;
    assign weights2[0][10] = 16'b1111111110001011;
    assign weights2[0][11] = 16'b0000000000001000;
    assign weights2[0][12] = 16'b1111111111010001;
    assign weights2[0][13] = 16'b1111111100110001;
    assign weights2[0][14] = 16'b1111111110101110;
    assign weights2[0][15] = 16'b0000000000011101;
    assign weights2[0][16] = 16'b0000000000010111;
    assign weights2[0][17] = 16'b0000000000110010;
    assign weights2[0][18] = 16'b1111111111111001;
    assign weights2[0][19] = 16'b1111111111110011;
    assign weights2[0][20] = 16'b1111111110100001;
    assign weights2[0][21] = 16'b0000000000011000;
    assign weights2[0][22] = 16'b0000000000000011;
    assign weights2[0][23] = 16'b0000000000001010;
    assign weights2[0][24] = 16'b1111111110111010;
    assign weights2[0][25] = 16'b0000000000000101;
    assign weights2[0][26] = 16'b0000000000001111;
    assign weights2[0][27] = 16'b1111111111010001;
    assign weights2[0][28] = 16'b1111111111100111;
    assign weights2[0][29] = 16'b0000000000000100;
    assign weights2[0][30] = 16'b0000000000000111;
    assign weights2[0][31] = 16'b1111111110011001;
    assign weights2[0][32] = 16'b0000000000011001;
    assign weights2[0][33] = 16'b0000000001000110;
    assign weights2[0][34] = 16'b1111111110100111;
    assign weights2[0][35] = 16'b1111111111100010;
    assign weights2[0][36] = 16'b1111111111010101;
    assign weights2[0][37] = 16'b1111111110011101;
    assign weights2[0][38] = 16'b1111111111100100;
    assign weights2[0][39] = 16'b1111111110011010;
    assign weights2[0][40] = 16'b0000000000001000;
    assign weights2[0][41] = 16'b1111111101100100;
    assign weights2[0][42] = 16'b0000000000011101;
    assign weights2[0][43] = 16'b1111111111001101;
    assign weights2[0][44] = 16'b0000000000100011;
    assign weights2[0][45] = 16'b0000000000101101;
    assign weights2[0][46] = 16'b1111111111111010;
    assign weights2[0][47] = 16'b1111111111110100;
    assign weights2[0][48] = 16'b0000000000101011;
    assign weights2[0][49] = 16'b0000000000100001;
    assign weights2[0][50] = 16'b1111111111011100;
    assign weights2[0][51] = 16'b0000000000001010;
    assign weights2[0][52] = 16'b0000000000101111;
    assign weights2[0][53] = 16'b1111111100100011;
    assign weights2[0][54] = 16'b0000000000000000;
    assign weights2[0][55] = 16'b0000000000010101;
    assign weights2[0][56] = 16'b1111111100010100;
    assign weights2[0][57] = 16'b1111111111101100;
    assign weights2[0][58] = 16'b1111111101010011;
    assign weights2[0][59] = 16'b1111111111111000;
    assign weights2[0][60] = 16'b0000000000001000;
    assign weights2[0][61] = 16'b0000000000011010;
    assign weights2[0][62] = 16'b0000000000001111;
    assign weights2[0][63] = 16'b1111111110001111;
    assign weights2[1][0] = 16'b1111111111110101;
    assign weights2[1][1] = 16'b0000000001100001;
    assign weights2[1][2] = 16'b1111111111001110;
    assign weights2[1][3] = 16'b1111111101111111;
    assign weights2[1][4] = 16'b1111111110010110;
    assign weights2[1][5] = 16'b0000000000001110;
    assign weights2[1][6] = 16'b0000000000000000;
    assign weights2[1][7] = 16'b0000000001110100;
    assign weights2[1][8] = 16'b0000000000011010;
    assign weights2[1][9] = 16'b1111111110110001;
    assign weights2[1][10] = 16'b0000000000100100;
    assign weights2[1][11] = 16'b1111111111111110;
    assign weights2[1][12] = 16'b0000000001101100;
    assign weights2[1][13] = 16'b0000000001111000;
    assign weights2[1][14] = 16'b1111111111110100;
    assign weights2[1][15] = 16'b0000000000001000;
    assign weights2[1][16] = 16'b0000000000001000;
    assign weights2[1][17] = 16'b1111111110110110;
    assign weights2[1][18] = 16'b1111111111110001;
    assign weights2[1][19] = 16'b1111111111010111;
    assign weights2[1][20] = 16'b1111111110010000;
    assign weights2[1][21] = 16'b1111111111010110;
    assign weights2[1][22] = 16'b1111111111100101;
    assign weights2[1][23] = 16'b1111111110110111;
    assign weights2[1][24] = 16'b1111111110000001;
    assign weights2[1][25] = 16'b1111111111110001;
    assign weights2[1][26] = 16'b1111111110011011;
    assign weights2[1][27] = 16'b0000000000100100;
    assign weights2[1][28] = 16'b0000000010010011;
    assign weights2[1][29] = 16'b1111111111100001;
    assign weights2[1][30] = 16'b1111111111110001;
    assign weights2[1][31] = 16'b1111111111111101;
    assign weights2[1][32] = 16'b1111111111100101;
    assign weights2[1][33] = 16'b1111111101111111;
    assign weights2[1][34] = 16'b1111111110000111;
    assign weights2[1][35] = 16'b1111111110110101;
    assign weights2[1][36] = 16'b0000000001001110;
    assign weights2[1][37] = 16'b1111111111110010;
    assign weights2[1][38] = 16'b1111111111011011;
    assign weights2[1][39] = 16'b0000000000010010;
    assign weights2[1][40] = 16'b0000000000000000;
    assign weights2[1][41] = 16'b0000000000110001;
    assign weights2[1][42] = 16'b1111111111001100;
    assign weights2[1][43] = 16'b1111111101010110;
    assign weights2[1][44] = 16'b0000000000001000;
    assign weights2[1][45] = 16'b1111111111011101;
    assign weights2[1][46] = 16'b0000000001101101;
    assign weights2[1][47] = 16'b0000000001001000;
    assign weights2[1][48] = 16'b0000000000101100;
    assign weights2[1][49] = 16'b1111111110111011;
    assign weights2[1][50] = 16'b0000000001010011;
    assign weights2[1][51] = 16'b0000000000000011;
    assign weights2[1][52] = 16'b1111111111000011;
    assign weights2[1][53] = 16'b0000000000010110;
    assign weights2[1][54] = 16'b0000000000000000;
    assign weights2[1][55] = 16'b1111111110111100;
    assign weights2[1][56] = 16'b0000000001101100;
    assign weights2[1][57] = 16'b1111111110101000;
    assign weights2[1][58] = 16'b0000000000011111;
    assign weights2[1][59] = 16'b1111111111011111;
    assign weights2[1][60] = 16'b1111111111110010;
    assign weights2[1][61] = 16'b1111111111011100;
    assign weights2[1][62] = 16'b0000000000101111;
    assign weights2[1][63] = 16'b1111111110111110;
    assign weights2[2][0] = 16'b0000000001111111;
    assign weights2[2][1] = 16'b1111111110100010;
    assign weights2[2][2] = 16'b0000000000011100;
    assign weights2[2][3] = 16'b0000000000000110;
    assign weights2[2][4] = 16'b1111111101110100;
    assign weights2[2][5] = 16'b0000000000001100;
    assign weights2[2][6] = 16'b0000000000000000;
    assign weights2[2][7] = 16'b1111111111110001;
    assign weights2[2][8] = 16'b0000000001001000;
    assign weights2[2][9] = 16'b1111111110101000;
    assign weights2[2][10] = 16'b1111111111011001;
    assign weights2[2][11] = 16'b1111111111100011;
    assign weights2[2][12] = 16'b1111111111110100;
    assign weights2[2][13] = 16'b1111111110011011;
    assign weights2[2][14] = 16'b0000000000000101;
    assign weights2[2][15] = 16'b0000000000101010;
    assign weights2[2][16] = 16'b0000000000111101;
    assign weights2[2][17] = 16'b0000000001011100;
    assign weights2[2][18] = 16'b0000000000011010;
    assign weights2[2][19] = 16'b0000000010000000;
    assign weights2[2][20] = 16'b0000000000010000;
    assign weights2[2][21] = 16'b0000000000111001;
    assign weights2[2][22] = 16'b0000000001111111;
    assign weights2[2][23] = 16'b0000000001010001;
    assign weights2[2][24] = 16'b1111111111111011;
    assign weights2[2][25] = 16'b0000000000010110;
    assign weights2[2][26] = 16'b1111111101101000;
    assign weights2[2][27] = 16'b0000000000111110;
    assign weights2[2][28] = 16'b1111111110100100;
    assign weights2[2][29] = 16'b1111111111111011;
    assign weights2[2][30] = 16'b0000000001110101;
    assign weights2[2][31] = 16'b1111111111111101;
    assign weights2[2][32] = 16'b0000000000010111;
    assign weights2[2][33] = 16'b1111111110010000;
    assign weights2[2][34] = 16'b1111111111111110;
    assign weights2[2][35] = 16'b1111111111011100;
    assign weights2[2][36] = 16'b1111111111111010;
    assign weights2[2][37] = 16'b1111111111111101;
    assign weights2[2][38] = 16'b0000000000100000;
    assign weights2[2][39] = 16'b1111111111001010;
    assign weights2[2][40] = 16'b0000000000000000;
    assign weights2[2][41] = 16'b1111111111101001;
    assign weights2[2][42] = 16'b0000000000100111;
    assign weights2[2][43] = 16'b0000000000000011;
    assign weights2[2][44] = 16'b0000000000100001;
    assign weights2[2][45] = 16'b0000000000000010;
    assign weights2[2][46] = 16'b1111111110110000;
    assign weights2[2][47] = 16'b1111111111011011;
    assign weights2[2][48] = 16'b0000000001000110;
    assign weights2[2][49] = 16'b0000000000110001;
    assign weights2[2][50] = 16'b1111111111111011;
    assign weights2[2][51] = 16'b1111111111111100;
    assign weights2[2][52] = 16'b0000000001000101;
    assign weights2[2][53] = 16'b1111111111011101;
    assign weights2[2][54] = 16'b0000000000000000;
    assign weights2[2][55] = 16'b1111111111001000;
    assign weights2[2][56] = 16'b1111111111010001;
    assign weights2[2][57] = 16'b1111111111111010;
    assign weights2[2][58] = 16'b1111111111101111;
    assign weights2[2][59] = 16'b0000000000000000;
    assign weights2[2][60] = 16'b0000000000001001;
    assign weights2[2][61] = 16'b0000000000011001;
    assign weights2[2][62] = 16'b0000000000110001;
    assign weights2[2][63] = 16'b1111111101010000;
    assign weights2[3][0] = 16'b1111111111111111;
    assign weights2[3][1] = 16'b1111111101111101;
    assign weights2[3][2] = 16'b1111111111111011;
    assign weights2[3][3] = 16'b1111111111100101;
    assign weights2[3][4] = 16'b1111111111100100;
    assign weights2[3][5] = 16'b1111111111001011;
    assign weights2[3][6] = 16'b0000000000000000;
    assign weights2[3][7] = 16'b1111111100011010;
    assign weights2[3][8] = 16'b1111111111010111;
    assign weights2[3][9] = 16'b1111111111111111;
    assign weights2[3][10] = 16'b1111111110011101;
    assign weights2[3][11] = 16'b1111111101011010;
    assign weights2[3][12] = 16'b1111111111111111;
    assign weights2[3][13] = 16'b1111111110000011;
    assign weights2[3][14] = 16'b1111111101110010;
    assign weights2[3][15] = 16'b0000000000001000;
    assign weights2[3][16] = 16'b1111111111111100;
    assign weights2[3][17] = 16'b1111111110001111;
    assign weights2[3][18] = 16'b1111111110001000;
    assign weights2[3][19] = 16'b1111111101111010;
    assign weights2[3][20] = 16'b1111111111111111;
    assign weights2[3][21] = 16'b1111111110101100;
    assign weights2[3][22] = 16'b1111111110111001;
    assign weights2[3][23] = 16'b1111111110010111;
    assign weights2[3][24] = 16'b0000000000011110;
    assign weights2[3][25] = 16'b0000000000001001;
    assign weights2[3][26] = 16'b1111111111110011;
    assign weights2[3][27] = 16'b1111111101010011;
    assign weights2[3][28] = 16'b0000000000001111;
    assign weights2[3][29] = 16'b0000000000010100;
    assign weights2[3][30] = 16'b1111111111110000;
    assign weights2[3][31] = 16'b1111111110010100;
    assign weights2[3][32] = 16'b0000000000011000;
    assign weights2[3][33] = 16'b1111111111111110;
    assign weights2[3][34] = 16'b1111111111110100;
    assign weights2[3][35] = 16'b1111111111111001;
    assign weights2[3][36] = 16'b1111111100111110;
    assign weights2[3][37] = 16'b1111111101111010;
    assign weights2[3][38] = 16'b1111111111110110;
    assign weights2[3][39] = 16'b1111111101111110;
    assign weights2[3][40] = 16'b1111111111111010;
    assign weights2[3][41] = 16'b1111111101111000;
    assign weights2[3][42] = 16'b0000000000101111;
    assign weights2[3][43] = 16'b0000000000100100;
    assign weights2[3][44] = 16'b0000000000001010;
    assign weights2[3][45] = 16'b0000000000010111;
    assign weights2[3][46] = 16'b0000000000101011;
    assign weights2[3][47] = 16'b1111111101111110;
    assign weights2[3][48] = 16'b0000000000011010;
    assign weights2[3][49] = 16'b0000000000100001;
    assign weights2[3][50] = 16'b0000000000001011;
    assign weights2[3][51] = 16'b0000000000010100;
    assign weights2[3][52] = 16'b0000000000100011;
    assign weights2[3][53] = 16'b1111111101100111;
    assign weights2[3][54] = 16'b0000000000000000;
    assign weights2[3][55] = 16'b0000000000010100;
    assign weights2[3][56] = 16'b1111111110111101;
    assign weights2[3][57] = 16'b0000000000110100;
    assign weights2[3][58] = 16'b1111111101101010;
    assign weights2[3][59] = 16'b0000000000011111;
    assign weights2[3][60] = 16'b1111111111111110;
    assign weights2[3][61] = 16'b0000000000011110;
    assign weights2[3][62] = 16'b0000000000001010;
    assign weights2[3][63] = 16'b1111111110001111;
    assign weights2[4][0] = 16'b1111111111101001;
    assign weights2[4][1] = 16'b1111111110011101;
    assign weights2[4][2] = 16'b0000000000111010;
    assign weights2[4][3] = 16'b0000000000100111;
    assign weights2[4][4] = 16'b0000000000010110;
    assign weights2[4][5] = 16'b0000000000011111;
    assign weights2[4][6] = 16'b0000000000000000;
    assign weights2[4][7] = 16'b1111111110000100;
    assign weights2[4][8] = 16'b1111111110100101;
    assign weights2[4][9] = 16'b0000000000000000;
    assign weights2[4][10] = 16'b0000000000000011;
    assign weights2[4][11] = 16'b0000000000001111;
    assign weights2[4][12] = 16'b1111111101011011;
    assign weights2[4][13] = 16'b1111111111000000;
    assign weights2[4][14] = 16'b0000000001101110;
    assign weights2[4][15] = 16'b1111111100111101;
    assign weights2[4][16] = 16'b1111111111110011;
    assign weights2[4][17] = 16'b0000000000011110;
    assign weights2[4][18] = 16'b1111111111111111;
    assign weights2[4][19] = 16'b0000000000010111;
    assign weights2[4][20] = 16'b0000000000110110;
    assign weights2[4][21] = 16'b0000000001000010;
    assign weights2[4][22] = 16'b0000000000000101;
    assign weights2[4][23] = 16'b1111111110111101;
    assign weights2[4][24] = 16'b0000000000110000;
    assign weights2[4][25] = 16'b0000000000001001;
    assign weights2[4][26] = 16'b1111111111111010;
    assign weights2[4][27] = 16'b1111111111100101;
    assign weights2[4][28] = 16'b1111111111111001;
    assign weights2[4][29] = 16'b0000000000000100;
    assign weights2[4][30] = 16'b0000000000100011;
    assign weights2[4][31] = 16'b0000000001011011;
    assign weights2[4][32] = 16'b0000000000001000;
    assign weights2[4][33] = 16'b1111111111011000;
    assign weights2[4][34] = 16'b0000000000101010;
    assign weights2[4][35] = 16'b1111111110001100;
    assign weights2[4][36] = 16'b1111111110101010;
    assign weights2[4][37] = 16'b0000000001100101;
    assign weights2[4][38] = 16'b0000000000100001;
    assign weights2[4][39] = 16'b0000000000101100;
    assign weights2[4][40] = 16'b1111111111001001;
    assign weights2[4][41] = 16'b0000000000011000;
    assign weights2[4][42] = 16'b0000000000110001;
    assign weights2[4][43] = 16'b0000000000101011;
    assign weights2[4][44] = 16'b0000000000000111;
    assign weights2[4][45] = 16'b1111111111100110;
    assign weights2[4][46] = 16'b0000000000010000;
    assign weights2[4][47] = 16'b1111111111010011;
    assign weights2[4][48] = 16'b1111111100000001;
    assign weights2[4][49] = 16'b0000000001000011;
    assign weights2[4][50] = 16'b0000000000000010;
    assign weights2[4][51] = 16'b0000000000000001;
    assign weights2[4][52] = 16'b1111111111101101;
    assign weights2[4][53] = 16'b0000000000111101;
    assign weights2[4][54] = 16'b0000000000000000;
    assign weights2[4][55] = 16'b1111111110001001;
    assign weights2[4][56] = 16'b0000000000010001;
    assign weights2[4][57] = 16'b0000000000101011;
    assign weights2[4][58] = 16'b0000000000101001;
    assign weights2[4][59] = 16'b0000000000000111;
    assign weights2[4][60] = 16'b1111111111111011;
    assign weights2[4][61] = 16'b0000000000011111;
    assign weights2[4][62] = 16'b1111111011111000;
    assign weights2[4][63] = 16'b1111111111111011;
    assign weights2[5][0] = 16'b0000000000001111;
    assign weights2[5][1] = 16'b1111111110101001;
    assign weights2[5][2] = 16'b0000000001000010;
    assign weights2[5][3] = 16'b0000000000110100;
    assign weights2[5][4] = 16'b0000000000110101;
    assign weights2[5][5] = 16'b0000000000010000;
    assign weights2[5][6] = 16'b0000000000000000;
    assign weights2[5][7] = 16'b1111111100001010;
    assign weights2[5][8] = 16'b1111111111001010;
    assign weights2[5][9] = 16'b0000000000001110;
    assign weights2[5][10] = 16'b1111111110110001;
    assign weights2[5][11] = 16'b0000000000010010;
    assign weights2[5][12] = 16'b1111111110000001;
    assign weights2[5][13] = 16'b1111111110101101;
    assign weights2[5][14] = 16'b0000000001110000;
    assign weights2[5][15] = 16'b1111111101101011;
    assign weights2[5][16] = 16'b0000000000100001;
    assign weights2[5][17] = 16'b1111111111110001;
    assign weights2[5][18] = 16'b0000000000001001;
    assign weights2[5][19] = 16'b0000000000100010;
    assign weights2[5][20] = 16'b0000000000101110;
    assign weights2[5][21] = 16'b0000000000111011;
    assign weights2[5][22] = 16'b0000000000100000;
    assign weights2[5][23] = 16'b1111111110100100;
    assign weights2[5][24] = 16'b0000000000000001;
    assign weights2[5][25] = 16'b0000000000010101;
    assign weights2[5][26] = 16'b0000000000010100;
    assign weights2[5][27] = 16'b1111111111011100;
    assign weights2[5][28] = 16'b1111111100010110;
    assign weights2[5][29] = 16'b1111111111011111;
    assign weights2[5][30] = 16'b1111111111110101;
    assign weights2[5][31] = 16'b0000000001011110;
    assign weights2[5][32] = 16'b0000000000110110;
    assign weights2[5][33] = 16'b0000000000001100;
    assign weights2[5][34] = 16'b0000000000010010;
    assign weights2[5][35] = 16'b1111111111101011;
    assign weights2[5][36] = 16'b1111111100110001;
    assign weights2[5][37] = 16'b0000000001110101;
    assign weights2[5][38] = 16'b1111111111101000;
    assign weights2[5][39] = 16'b0000000000010110;
    assign weights2[5][40] = 16'b1111111111101110;
    assign weights2[5][41] = 16'b0000000000000101;
    assign weights2[5][42] = 16'b0000000001101000;
    assign weights2[5][43] = 16'b1111111111110000;
    assign weights2[5][44] = 16'b0000000000101100;
    assign weights2[5][45] = 16'b0000000000000000;
    assign weights2[5][46] = 16'b1111111101101101;
    assign weights2[5][47] = 16'b1111111111011110;
    assign weights2[5][48] = 16'b1111111111001110;
    assign weights2[5][49] = 16'b0000000001011011;
    assign weights2[5][50] = 16'b1111111110101110;
    assign weights2[5][51] = 16'b0000000000000101;
    assign weights2[5][52] = 16'b0000000000110010;
    assign weights2[5][53] = 16'b0000000000110100;
    assign weights2[5][54] = 16'b0000000000000000;
    assign weights2[5][55] = 16'b1111111111111100;
    assign weights2[5][56] = 16'b0000000000011010;
    assign weights2[5][57] = 16'b1111111111111111;
    assign weights2[5][58] = 16'b1111111111111101;
    assign weights2[5][59] = 16'b0000000000010100;
    assign weights2[5][60] = 16'b0000000000101101;
    assign weights2[5][61] = 16'b0000000001000110;
    assign weights2[5][62] = 16'b1111111111100100;
    assign weights2[5][63] = 16'b0000000000001101;
    assign weights2[6][0] = 16'b0000000000000110;
    assign weights2[6][1] = 16'b0000000001000101;
    assign weights2[6][2] = 16'b1111111111000010;
    assign weights2[6][3] = 16'b0000000000000100;
    assign weights2[6][4] = 16'b1111111111110001;
    assign weights2[6][5] = 16'b1111111111010001;
    assign weights2[6][6] = 16'b0000000000000000;
    assign weights2[6][7] = 16'b1111111100101010;
    assign weights2[6][8] = 16'b1111111101111110;
    assign weights2[6][9] = 16'b0000000000100101;
    assign weights2[6][10] = 16'b1111111110011010;
    assign weights2[6][11] = 16'b1111111100010100;
    assign weights2[6][12] = 16'b0000000000111010;
    assign weights2[6][13] = 16'b0000000000111101;
    assign weights2[6][14] = 16'b1111111111111111;
    assign weights2[6][15] = 16'b1111111110111000;
    assign weights2[6][16] = 16'b0000000000001111;
    assign weights2[6][17] = 16'b1111111100111010;
    assign weights2[6][18] = 16'b1111111101000111;
    assign weights2[6][19] = 16'b1111111101000011;
    assign weights2[6][20] = 16'b1111111111011001;
    assign weights2[6][21] = 16'b1111111101101010;
    assign weights2[6][22] = 16'b1111111110011010;
    assign weights2[6][23] = 16'b1111111101010000;
    assign weights2[6][24] = 16'b0000000000000101;
    assign weights2[6][25] = 16'b1111111111110011;
    assign weights2[6][26] = 16'b1111111111011010;
    assign weights2[6][27] = 16'b1111111111000001;
    assign weights2[6][28] = 16'b1111111101101110;
    assign weights2[6][29] = 16'b0000000000000111;
    assign weights2[6][30] = 16'b1111111110011111;
    assign weights2[6][31] = 16'b1111111111111100;
    assign weights2[6][32] = 16'b0000000000101010;
    assign weights2[6][33] = 16'b1111111111110001;
    assign weights2[6][34] = 16'b1111111111111001;
    assign weights2[6][35] = 16'b1111111111111100;
    assign weights2[6][36] = 16'b1111111110000001;
    assign weights2[6][37] = 16'b0000000000000001;
    assign weights2[6][38] = 16'b1111111111011000;
    assign weights2[6][39] = 16'b1111111110011100;
    assign weights2[6][40] = 16'b1111111111101100;
    assign weights2[6][41] = 16'b1111111111110011;
    assign weights2[6][42] = 16'b1111111111010111;
    assign weights2[6][43] = 16'b0000000000010010;
    assign weights2[6][44] = 16'b0000000000011100;
    assign weights2[6][45] = 16'b0000000000011001;
    assign weights2[6][46] = 16'b1111111111101000;
    assign weights2[6][47] = 16'b1111111110100111;
    assign weights2[6][48] = 16'b1111111111110011;
    assign weights2[6][49] = 16'b1111111110100110;
    assign weights2[6][50] = 16'b1111111111110101;
    assign weights2[6][51] = 16'b0000000000001111;
    assign weights2[6][52] = 16'b1111111110100001;
    assign weights2[6][53] = 16'b0000000000001100;
    assign weights2[6][54] = 16'b0000000000000000;
    assign weights2[6][55] = 16'b0000000001000000;
    assign weights2[6][56] = 16'b0000000000101010;
    assign weights2[6][57] = 16'b0000000000001100;
    assign weights2[6][58] = 16'b1111111101110101;
    assign weights2[6][59] = 16'b0000000000010110;
    assign weights2[6][60] = 16'b1111111111110011;
    assign weights2[6][61] = 16'b1111111111111010;
    assign weights2[6][62] = 16'b0000000000001100;
    assign weights2[6][63] = 16'b0000000000101000;
    assign weights2[7][0] = 16'b0000000000010101;
    assign weights2[7][1] = 16'b1111111101011000;
    assign weights2[7][2] = 16'b0000000000011000;
    assign weights2[7][3] = 16'b1111111111111111;
    assign weights2[7][4] = 16'b1111111100000011;
    assign weights2[7][5] = 16'b1111111111101010;
    assign weights2[7][6] = 16'b0000000000000000;
    assign weights2[7][7] = 16'b1111111111011111;
    assign weights2[7][8] = 16'b0000000001000001;
    assign weights2[7][9] = 16'b1111111100110111;
    assign weights2[7][10] = 16'b0000000000001011;
    assign weights2[7][11] = 16'b1111111111100010;
    assign weights2[7][12] = 16'b1111111101000110;
    assign weights2[7][13] = 16'b1111111101101110;
    assign weights2[7][14] = 16'b0000000000010010;
    assign weights2[7][15] = 16'b1111111111100001;
    assign weights2[7][16] = 16'b0000000000011101;
    assign weights2[7][17] = 16'b0000000000110000;
    assign weights2[7][18] = 16'b0000000000001101;
    assign weights2[7][19] = 16'b0000000000000111;
    assign weights2[7][20] = 16'b1111111111110001;
    assign weights2[7][21] = 16'b0000000000101110;
    assign weights2[7][22] = 16'b0000000000100101;
    assign weights2[7][23] = 16'b0000000001000000;
    assign weights2[7][24] = 16'b0000000000001011;
    assign weights2[7][25] = 16'b0000000000001111;
    assign weights2[7][26] = 16'b1111111100111101;
    assign weights2[7][27] = 16'b1111111111001101;
    assign weights2[7][28] = 16'b1111111110110101;
    assign weights2[7][29] = 16'b1111111111111111;
    assign weights2[7][30] = 16'b1111111111111111;
    assign weights2[7][31] = 16'b0000000000001001;
    assign weights2[7][32] = 16'b1111111111111010;
    assign weights2[7][33] = 16'b1111111110010110;
    assign weights2[7][34] = 16'b0000000000000000;
    assign weights2[7][35] = 16'b1111111110101110;
    assign weights2[7][36] = 16'b0000000000010001;
    assign weights2[7][37] = 16'b0000000000010110;
    assign weights2[7][38] = 16'b0000000000100001;
    assign weights2[7][39] = 16'b1111111111100100;
    assign weights2[7][40] = 16'b1111111111110011;
    assign weights2[7][41] = 16'b1111111111101110;
    assign weights2[7][42] = 16'b0000000000100110;
    assign weights2[7][43] = 16'b0000000000001100;
    assign weights2[7][44] = 16'b1111111111110001;
    assign weights2[7][45] = 16'b0000000000000110;
    assign weights2[7][46] = 16'b1111111111110010;
    assign weights2[7][47] = 16'b1111111110000111;
    assign weights2[7][48] = 16'b1111111111001101;
    assign weights2[7][49] = 16'b0000000000100000;
    assign weights2[7][50] = 16'b0000000000011110;
    assign weights2[7][51] = 16'b0000000000000100;
    assign weights2[7][52] = 16'b0000000000010000;
    assign weights2[7][53] = 16'b1111111111111001;
    assign weights2[7][54] = 16'b0000000000000000;
    assign weights2[7][55] = 16'b1111111100011111;
    assign weights2[7][56] = 16'b1111111110100111;
    assign weights2[7][57] = 16'b0000000000001011;
    assign weights2[7][58] = 16'b0000000000001110;
    assign weights2[7][59] = 16'b0000000000010010;
    assign weights2[7][60] = 16'b0000000000100001;
    assign weights2[7][61] = 16'b0000000000011010;
    assign weights2[7][62] = 16'b1111111111001110;
    assign weights2[7][63] = 16'b1111111110011000;
    assign weights2[8][0] = 16'b1111111111000101;
    assign weights2[8][1] = 16'b0000000000011101;
    assign weights2[8][2] = 16'b1111111111011000;
    assign weights2[8][3] = 16'b1111111111000011;
    assign weights2[8][4] = 16'b1111111111010101;
    assign weights2[8][5] = 16'b1111111111001111;
    assign weights2[8][6] = 16'b0000000000000000;
    assign weights2[8][7] = 16'b0000000010110011;
    assign weights2[8][8] = 16'b0000000000111001;
    assign weights2[8][9] = 16'b1111111111110010;
    assign weights2[8][10] = 16'b0000000001011111;
    assign weights2[8][11] = 16'b0000000000000010;
    assign weights2[8][12] = 16'b0000000000101111;
    assign weights2[8][13] = 16'b0000000000011110;
    assign weights2[8][14] = 16'b1111111110011111;
    assign weights2[8][15] = 16'b0000000000001100;
    assign weights2[8][16] = 16'b1111111111111111;
    assign weights2[8][17] = 16'b0000000000011111;
    assign weights2[8][18] = 16'b0000000000000011;
    assign weights2[8][19] = 16'b0000000000010000;
    assign weights2[8][20] = 16'b1111111101111111;
    assign weights2[8][21] = 16'b1111111111011011;
    assign weights2[8][22] = 16'b0000000000001000;
    assign weights2[8][23] = 16'b0000000000010111;
    assign weights2[8][24] = 16'b0000000000010010;
    assign weights2[8][25] = 16'b1111111111011000;
    assign weights2[8][26] = 16'b1111111111101000;
    assign weights2[8][27] = 16'b0000000000011011;
    assign weights2[8][28] = 16'b0000000010011100;
    assign weights2[8][29] = 16'b0000000000011100;
    assign weights2[8][30] = 16'b0000000000001000;
    assign weights2[8][31] = 16'b1111111111000001;
    assign weights2[8][32] = 16'b1111111110101111;
    assign weights2[8][33] = 16'b0000000000010100;
    assign weights2[8][34] = 16'b1111111110110010;
    assign weights2[8][35] = 16'b1111111111110100;
    assign weights2[8][36] = 16'b0000000001000100;
    assign weights2[8][37] = 16'b1111111101100110;
    assign weights2[8][38] = 16'b1111111111111010;
    assign weights2[8][39] = 16'b1111111110101100;
    assign weights2[8][40] = 16'b0000000000000000;
    assign weights2[8][41] = 16'b0000000000101111;
    assign weights2[8][42] = 16'b1111111110101011;
    assign weights2[8][43] = 16'b0000000000010100;
    assign weights2[8][44] = 16'b1111111111001000;
    assign weights2[8][45] = 16'b0000000000000101;
    assign weights2[8][46] = 16'b0000000010001111;
    assign weights2[8][47] = 16'b0000000000001011;
    assign weights2[8][48] = 16'b0000000000010010;
    assign weights2[8][49] = 16'b1111111111000000;
    assign weights2[8][50] = 16'b0000000010011100;
    assign weights2[8][51] = 16'b1111111111110010;
    assign weights2[8][52] = 16'b1111111110101110;
    assign weights2[8][53] = 16'b1111111110110111;
    assign weights2[8][54] = 16'b1111111111111111;
    assign weights2[8][55] = 16'b1111111111001011;
    assign weights2[8][56] = 16'b0000000000000010;
    assign weights2[8][57] = 16'b0000000000001011;
    assign weights2[8][58] = 16'b0000000000011110;
    assign weights2[8][59] = 16'b1111111111001000;
    assign weights2[8][60] = 16'b1111111111100100;
    assign weights2[8][61] = 16'b1111111111011011;
    assign weights2[8][62] = 16'b0000000000010101;
    assign weights2[8][63] = 16'b1111111101000011;
    assign weights2[9][0] = 16'b0000000000001100;
    assign weights2[9][1] = 16'b1111111110010101;
    assign weights2[9][2] = 16'b0000000001001001;
    assign weights2[9][3] = 16'b0000000000111010;
    assign weights2[9][4] = 16'b0000000000110111;
    assign weights2[9][5] = 16'b0000000000010110;
    assign weights2[9][6] = 16'b0000000000000000;
    assign weights2[9][7] = 16'b0000000000111000;
    assign weights2[9][8] = 16'b0000000000100111;
    assign weights2[9][9] = 16'b0000000000010111;
    assign weights2[9][10] = 16'b1111111111100011;
    assign weights2[9][11] = 16'b0000000001001001;
    assign weights2[9][12] = 16'b1111111110001001;
    assign weights2[9][13] = 16'b1111111110101111;
    assign weights2[9][14] = 16'b0000000000101010;
    assign weights2[9][15] = 16'b1111111111100111;
    assign weights2[9][16] = 16'b1111111111111011;
    assign weights2[9][17] = 16'b0000000010001011;
    assign weights2[9][18] = 16'b0000000000110111;
    assign weights2[9][19] = 16'b0000000000111110;
    assign weights2[9][20] = 16'b1111111101011110;
    assign weights2[9][21] = 16'b0000000001111100;
    assign weights2[9][22] = 16'b0000000001001110;
    assign weights2[9][23] = 16'b0000000000101111;
    assign weights2[9][24] = 16'b0000000000101001;
    assign weights2[9][25] = 16'b1111111111111101;
    assign weights2[9][26] = 16'b0000000001001001;
    assign weights2[9][27] = 16'b0000000000000010;
    assign weights2[9][28] = 16'b0000000000010111;
    assign weights2[9][29] = 16'b1111111111111001;
    assign weights2[9][30] = 16'b0000000000101011;
    assign weights2[9][31] = 16'b0000000000100100;
    assign weights2[9][32] = 16'b1111111111111110;
    assign weights2[9][33] = 16'b0000000010100010;
    assign weights2[9][34] = 16'b0000000000011000;
    assign weights2[9][35] = 16'b1111111111000001;
    assign weights2[9][36] = 16'b0000000000001100;
    assign weights2[9][37] = 16'b0000000000110000;
    assign weights2[9][38] = 16'b0000000000110100;
    assign weights2[9][39] = 16'b0000000000110011;
    assign weights2[9][40] = 16'b1111111111011001;
    assign weights2[9][41] = 16'b1111111111001110;
    assign weights2[9][42] = 16'b0000000000100100;
    assign weights2[9][43] = 16'b0000000000111110;
    assign weights2[9][44] = 16'b0000000000000010;
    assign weights2[9][45] = 16'b0000000000001101;
    assign weights2[9][46] = 16'b0000000000001010;
    assign weights2[9][47] = 16'b0000000000000001;
    assign weights2[9][48] = 16'b1111111111101001;
    assign weights2[9][49] = 16'b0000000000011001;
    assign weights2[9][50] = 16'b0000000000001011;
    assign weights2[9][51] = 16'b1111111111010001;
    assign weights2[9][52] = 16'b0000000001001001;
    assign weights2[9][53] = 16'b0000000000110010;
    assign weights2[9][54] = 16'b0000000000000000;
    assign weights2[9][55] = 16'b0000000000101111;
    assign weights2[9][56] = 16'b1111111110111001;
    assign weights2[9][57] = 16'b0000000000100001;
    assign weights2[9][58] = 16'b1111111111001111;
    assign weights2[9][59] = 16'b0000000000000111;
    assign weights2[9][60] = 16'b1111111111100010;
    assign weights2[9][61] = 16'b0000000000011001;
    assign weights2[9][62] = 16'b1111111111110111;
    assign weights2[9][63] = 16'b0000000001000111;
    assign weights2[10][0] = 16'b0000000000011011;
    assign weights2[10][1] = 16'b0000000001101000;
    assign weights2[10][2] = 16'b1111111111010110;
    assign weights2[10][3] = 16'b1111111110010100;
    assign weights2[10][4] = 16'b1111111111110011;
    assign weights2[10][5] = 16'b0000000000001001;
    assign weights2[10][6] = 16'b0000000000000000;
    assign weights2[10][7] = 16'b0000000000010011;
    assign weights2[10][8] = 16'b0000000000011011;
    assign weights2[10][9] = 16'b0000000000001000;
    assign weights2[10][10] = 16'b0000000000010100;
    assign weights2[10][11] = 16'b0000000001111100;
    assign weights2[10][12] = 16'b0000000001000001;
    assign weights2[10][13] = 16'b0000000001101101;
    assign weights2[10][14] = 16'b0000000000111000;
    assign weights2[10][15] = 16'b1111111111111101;
    assign weights2[10][16] = 16'b0000000000110101;
    assign weights2[10][17] = 16'b0000000000111110;
    assign weights2[10][18] = 16'b0000000001110101;
    assign weights2[10][19] = 16'b0000000001010111;
    assign weights2[10][20] = 16'b0000000000100000;
    assign weights2[10][21] = 16'b0000000000111100;
    assign weights2[10][22] = 16'b0000000001111011;
    assign weights2[10][23] = 16'b0000000000101101;
    assign weights2[10][24] = 16'b1111111101011010;
    assign weights2[10][25] = 16'b1111111111110000;
    assign weights2[10][26] = 16'b0000000000000100;
    assign weights2[10][27] = 16'b0000000010111001;
    assign weights2[10][28] = 16'b1111111111100111;
    assign weights2[10][29] = 16'b1111111110110110;
    assign weights2[10][30] = 16'b1111111111110001;
    assign weights2[10][31] = 16'b0000000000110110;
    assign weights2[10][32] = 16'b0000000000000100;
    assign weights2[10][33] = 16'b1111111111100000;
    assign weights2[10][34] = 16'b1111111110100000;
    assign weights2[10][35] = 16'b1111111110101001;
    assign weights2[10][36] = 16'b0000000000100101;
    assign weights2[10][37] = 16'b0000000000110001;
    assign weights2[10][38] = 16'b1111111111100000;
    assign weights2[10][39] = 16'b1111111111111101;
    assign weights2[10][40] = 16'b1111111111111001;
    assign weights2[10][41] = 16'b0000000000011011;
    assign weights2[10][42] = 16'b1111111111100110;
    assign weights2[10][43] = 16'b1111111101101111;
    assign weights2[10][44] = 16'b1111111111111011;
    assign weights2[10][45] = 16'b1111111111010101;
    assign weights2[10][46] = 16'b0000000000011100;
    assign weights2[10][47] = 16'b0000000001110000;
    assign weights2[10][48] = 16'b1111111111110000;
    assign weights2[10][49] = 16'b1111111111110010;
    assign weights2[10][50] = 16'b0000000000100110;
    assign weights2[10][51] = 16'b1111111111100101;
    assign weights2[10][52] = 16'b1111111111111101;
    assign weights2[10][53] = 16'b0000000000010110;
    assign weights2[10][54] = 16'b0000000000000000;
    assign weights2[10][55] = 16'b1111111111110110;
    assign weights2[10][56] = 16'b0000000000110100;
    assign weights2[10][57] = 16'b1111111110001101;
    assign weights2[10][58] = 16'b0000000000000010;
    assign weights2[10][59] = 16'b1111111111101001;
    assign weights2[10][60] = 16'b0000000001000001;
    assign weights2[10][61] = 16'b1111111111110000;
    assign weights2[10][62] = 16'b1111111111110001;
    assign weights2[10][63] = 16'b1111111111010101;
    assign weights2[11][0] = 16'b0000000000000100;
    assign weights2[11][1] = 16'b1111111101111111;
    assign weights2[11][2] = 16'b1111111111100000;
    assign weights2[11][3] = 16'b1111111111001001;
    assign weights2[11][4] = 16'b0000000000010101;
    assign weights2[11][5] = 16'b1111111111101111;
    assign weights2[11][6] = 16'b0000000000000000;
    assign weights2[11][7] = 16'b0000000000010010;
    assign weights2[11][8] = 16'b0000000000111111;
    assign weights2[11][9] = 16'b0000000000000100;
    assign weights2[11][10] = 16'b1111111111001101;
    assign weights2[11][11] = 16'b1111111111111011;
    assign weights2[11][12] = 16'b1111111111000011;
    assign weights2[11][13] = 16'b1111111101011101;
    assign weights2[11][14] = 16'b1111111110010001;
    assign weights2[11][15] = 16'b1111111111101010;
    assign weights2[11][16] = 16'b0000000000100101;
    assign weights2[11][17] = 16'b1111111111010110;
    assign weights2[11][18] = 16'b0000000000001000;
    assign weights2[11][19] = 16'b1111111111011111;
    assign weights2[11][20] = 16'b1111111100100011;
    assign weights2[11][21] = 16'b0000000000001011;
    assign weights2[11][22] = 16'b0000000000011110;
    assign weights2[11][23] = 16'b0000000000101110;
    assign weights2[11][24] = 16'b1111111111100000;
    assign weights2[11][25] = 16'b1111111111001110;
    assign weights2[11][26] = 16'b0000000000001010;
    assign weights2[11][27] = 16'b1111111110000111;
    assign weights2[11][28] = 16'b1111111111000001;
    assign weights2[11][29] = 16'b1111111110110000;
    assign weights2[11][30] = 16'b1111111110101011;
    assign weights2[11][31] = 16'b1111111110010001;
    assign weights2[11][32] = 16'b1111111111010111;
    assign weights2[11][33] = 16'b0000000000110100;
    assign weights2[11][34] = 16'b1111111111000111;
    assign weights2[11][35] = 16'b0000000000001010;
    assign weights2[11][36] = 16'b0000000000101100;
    assign weights2[11][37] = 16'b1111111111000101;
    assign weights2[11][38] = 16'b1111111111101000;
    assign weights2[11][39] = 16'b1111111111010111;
    assign weights2[11][40] = 16'b0000000000001001;
    assign weights2[11][41] = 16'b1111111111110110;
    assign weights2[11][42] = 16'b1111111101101100;
    assign weights2[11][43] = 16'b1111111111100010;
    assign weights2[11][44] = 16'b1111111111110010;
    assign weights2[11][45] = 16'b0000000000001100;
    assign weights2[11][46] = 16'b1111111111111000;
    assign weights2[11][47] = 16'b1111111111010100;
    assign weights2[11][48] = 16'b1111111111111010;
    assign weights2[11][49] = 16'b1111111111000011;
    assign weights2[11][50] = 16'b1111111111100101;
    assign weights2[11][51] = 16'b0000000000000000;
    assign weights2[11][52] = 16'b1111111111110101;
    assign weights2[11][53] = 16'b1111111111100001;
    assign weights2[11][54] = 16'b0000000000000000;
    assign weights2[11][55] = 16'b1111111111001000;
    assign weights2[11][56] = 16'b1111111110111111;
    assign weights2[11][57] = 16'b1111111111010111;
    assign weights2[11][58] = 16'b1111111111111010;
    assign weights2[11][59] = 16'b1111111111000010;
    assign weights2[11][60] = 16'b1111111111011101;
    assign weights2[11][61] = 16'b1111111110111110;
    assign weights2[11][62] = 16'b0000000000001111;
    assign weights2[11][63] = 16'b0000000000100011;
    assign weights2[12][0] = 16'b1111111101111001;
    assign weights2[12][1] = 16'b0000000000000101;
    assign weights2[12][2] = 16'b0000000001010011;
    assign weights2[12][3] = 16'b0000000000111001;
    assign weights2[12][4] = 16'b1111111111111111;
    assign weights2[12][5] = 16'b1111111101100000;
    assign weights2[12][6] = 16'b0000000000000000;
    assign weights2[12][7] = 16'b0000000000100001;
    assign weights2[12][8] = 16'b0000000000011000;
    assign weights2[12][9] = 16'b1111111111100100;
    assign weights2[12][10] = 16'b1111111111100001;
    assign weights2[12][11] = 16'b0000000000100001;
    assign weights2[12][12] = 16'b1111111111101111;
    assign weights2[12][13] = 16'b0000000000001100;
    assign weights2[12][14] = 16'b0000000000011011;
    assign weights2[12][15] = 16'b0000000000000100;
    assign weights2[12][16] = 16'b1111111111100100;
    assign weights2[12][17] = 16'b0000000000100111;
    assign weights2[12][18] = 16'b0000000000001000;
    assign weights2[12][19] = 16'b0000000000001001;
    assign weights2[12][20] = 16'b0000000000011111;
    assign weights2[12][21] = 16'b0000000001101011;
    assign weights2[12][22] = 16'b1111111111011010;
    assign weights2[12][23] = 16'b0000000000001010;
    assign weights2[12][24] = 16'b0000000010111111;
    assign weights2[12][25] = 16'b0000000000110101;
    assign weights2[12][26] = 16'b0000000000011110;
    assign weights2[12][27] = 16'b0000000000101011;
    assign weights2[12][28] = 16'b0000000000101010;
    assign weights2[12][29] = 16'b0000000010001110;
    assign weights2[12][30] = 16'b0000000000000000;
    assign weights2[12][31] = 16'b0000000000011011;
    assign weights2[12][32] = 16'b1111111111010100;
    assign weights2[12][33] = 16'b0000000000000001;
    assign weights2[12][34] = 16'b0000000001000000;
    assign weights2[12][35] = 16'b0000000001100101;
    assign weights2[12][36] = 16'b1111111111110110;
    assign weights2[12][37] = 16'b0000000000010111;
    assign weights2[12][38] = 16'b0000000000011011;
    assign weights2[12][39] = 16'b0000000000001110;
    assign weights2[12][40] = 16'b1111111111100010;
    assign weights2[12][41] = 16'b0000000000001001;
    assign weights2[12][42] = 16'b0000000001001100;
    assign weights2[12][43] = 16'b0000000010011011;
    assign weights2[12][44] = 16'b1111111110101011;
    assign weights2[12][45] = 16'b0000000001001111;
    assign weights2[12][46] = 16'b0000000000101111;
    assign weights2[12][47] = 16'b0000000000100101;
    assign weights2[12][48] = 16'b0000000000100100;
    assign weights2[12][49] = 16'b0000000001110111;
    assign weights2[12][50] = 16'b0000000001101101;
    assign weights2[12][51] = 16'b0000000000011001;
    assign weights2[12][52] = 16'b0000000000111011;
    assign weights2[12][53] = 16'b0000000000011000;
    assign weights2[12][54] = 16'b0000000000000000;
    assign weights2[12][55] = 16'b0000000000001000;
    assign weights2[12][56] = 16'b0000000000001100;
    assign weights2[12][57] = 16'b0000000010010111;
    assign weights2[12][58] = 16'b1111111111100011;
    assign weights2[12][59] = 16'b0000000000100000;
    assign weights2[12][60] = 16'b0000000000100000;
    assign weights2[12][61] = 16'b0000000001011111;
    assign weights2[12][62] = 16'b0000000000111001;
    assign weights2[12][63] = 16'b1111111111101101;
    assign weights2[13][0] = 16'b1111111111011100;
    assign weights2[13][1] = 16'b1111111101111111;
    assign weights2[13][2] = 16'b0000000000000111;
    assign weights2[13][3] = 16'b0000000000101001;
    assign weights2[13][4] = 16'b1111111110100011;
    assign weights2[13][5] = 16'b1111111111111100;
    assign weights2[13][6] = 16'b0000000000000000;
    assign weights2[13][7] = 16'b1111111111110110;
    assign weights2[13][8] = 16'b0000000000010000;
    assign weights2[13][9] = 16'b1111111110010010;
    assign weights2[13][10] = 16'b0000000000010111;
    assign weights2[13][11] = 16'b1111111111001110;
    assign weights2[13][12] = 16'b1111111110001011;
    assign weights2[13][13] = 16'b1111111110100100;
    assign weights2[13][14] = 16'b0000000000000110;
    assign weights2[13][15] = 16'b1111111111111101;
    assign weights2[13][16] = 16'b1111111111111110;
    assign weights2[13][17] = 16'b1111111110110111;
    assign weights2[13][18] = 16'b1111111111001011;
    assign weights2[13][19] = 16'b1111111110101101;
    assign weights2[13][20] = 16'b1111111110100011;
    assign weights2[13][21] = 16'b1111111110111111;
    assign weights2[13][22] = 16'b1111111110110111;
    assign weights2[13][23] = 16'b0000000000001001;
    assign weights2[13][24] = 16'b1111111111111111;
    assign weights2[13][25] = 16'b1111111111111110;
    assign weights2[13][26] = 16'b1111111110011100;
    assign weights2[13][27] = 16'b1111111110000100;
    assign weights2[13][28] = 16'b1111111111000101;
    assign weights2[13][29] = 16'b1111111111110111;
    assign weights2[13][30] = 16'b1111111111010110;
    assign weights2[13][31] = 16'b1111111111111111;
    assign weights2[13][32] = 16'b1111111111101111;
    assign weights2[13][33] = 16'b1111111111001001;
    assign weights2[13][34] = 16'b0000000000000111;
    assign weights2[13][35] = 16'b1111111111001000;
    assign weights2[13][36] = 16'b0000000000011101;
    assign weights2[13][37] = 16'b0000000000001100;
    assign weights2[13][38] = 16'b0000000000010111;
    assign weights2[13][39] = 16'b1111111111110111;
    assign weights2[13][40] = 16'b0000000000001011;
    assign weights2[13][41] = 16'b1111111111111111;
    assign weights2[13][42] = 16'b1111111111010101;
    assign weights2[13][43] = 16'b0000000000100110;
    assign weights2[13][44] = 16'b1111111111110010;
    assign weights2[13][45] = 16'b0000000000101011;
    assign weights2[13][46] = 16'b1111111111001010;
    assign weights2[13][47] = 16'b1111111110111001;
    assign weights2[13][48] = 16'b1111111111010010;
    assign weights2[13][49] = 16'b1111111111110100;
    assign weights2[13][50] = 16'b1111111110101001;
    assign weights2[13][51] = 16'b0000000000001101;
    assign weights2[13][52] = 16'b1111111101111011;
    assign weights2[13][53] = 16'b1111111111101001;
    assign weights2[13][54] = 16'b0000000000000000;
    assign weights2[13][55] = 16'b1111111110110101;
    assign weights2[13][56] = 16'b1111111110011101;
    assign weights2[13][57] = 16'b0000000000101011;
    assign weights2[13][58] = 16'b0000000000100110;
    assign weights2[13][59] = 16'b1111111111000101;
    assign weights2[13][60] = 16'b1111111110110111;
    assign weights2[13][61] = 16'b1111111111110101;
    assign weights2[13][62] = 16'b1111111110101101;
    assign weights2[13][63] = 16'b1111111111111010;
    assign weights2[14][0] = 16'b0000000000000111;
    assign weights2[14][1] = 16'b1111111111101000;
    assign weights2[14][2] = 16'b1111111110100011;
    assign weights2[14][3] = 16'b1111111101111000;
    assign weights2[14][4] = 16'b1111111111010010;
    assign weights2[14][5] = 16'b1111111110100010;
    assign weights2[14][6] = 16'b0000000000000000;
    assign weights2[14][7] = 16'b1111111111111100;
    assign weights2[14][8] = 16'b1111111110100110;
    assign weights2[14][9] = 16'b1111111111101100;
    assign weights2[14][10] = 16'b1111111111000100;
    assign weights2[14][11] = 16'b1111111110101010;
    assign weights2[14][12] = 16'b1111111111101010;
    assign weights2[14][13] = 16'b1111111111100100;
    assign weights2[14][14] = 16'b0000000000000110;
    assign weights2[14][15] = 16'b0000000000000010;
    assign weights2[14][16] = 16'b0000000001001101;
    assign weights2[14][17] = 16'b1111111110101100;
    assign weights2[14][18] = 16'b1111111111000011;
    assign weights2[14][19] = 16'b1111111110110001;
    assign weights2[14][20] = 16'b0000000001100011;
    assign weights2[14][21] = 16'b1111111111101100;
    assign weights2[14][22] = 16'b1111111111101110;
    assign weights2[14][23] = 16'b1111111111100110;
    assign weights2[14][24] = 16'b1111111101011011;
    assign weights2[14][25] = 16'b0000000000100011;
    assign weights2[14][26] = 16'b1111111110111111;
    assign weights2[14][27] = 16'b1111111111001110;
    assign weights2[14][28] = 16'b0000000001001100;
    assign weights2[14][29] = 16'b1111111110110010;
    assign weights2[14][30] = 16'b1111111110011101;
    assign weights2[14][31] = 16'b0000000000000111;
    assign weights2[14][32] = 16'b0000000000010100;
    assign weights2[14][33] = 16'b1111111110110011;
    assign weights2[14][34] = 16'b1111111110000111;
    assign weights2[14][35] = 16'b1111111110001100;
    assign weights2[14][36] = 16'b1111111111011001;
    assign weights2[14][37] = 16'b0000000000000010;
    assign weights2[14][38] = 16'b1111111111001000;
    assign weights2[14][39] = 16'b1111111111110011;
    assign weights2[14][40] = 16'b1111111111110111;
    assign weights2[14][41] = 16'b0000000000001101;
    assign weights2[14][42] = 16'b0000000000011111;
    assign weights2[14][43] = 16'b1111111101101100;
    assign weights2[14][44] = 16'b0000000000011100;
    assign weights2[14][45] = 16'b1111111111010010;
    assign weights2[14][46] = 16'b0000000001010000;
    assign weights2[14][47] = 16'b1111111111011101;
    assign weights2[14][48] = 16'b1111111111100011;
    assign weights2[14][49] = 16'b0000000000101010;
    assign weights2[14][50] = 16'b0000000000001100;
    assign weights2[14][51] = 16'b0000000000010110;
    assign weights2[14][52] = 16'b0000000000011111;
    assign weights2[14][53] = 16'b0000000000001011;
    assign weights2[14][54] = 16'b0000000000000000;
    assign weights2[14][55] = 16'b1111111111101101;
    assign weights2[14][56] = 16'b0000000000000011;
    assign weights2[14][57] = 16'b1111111101111110;
    assign weights2[14][58] = 16'b0000000000000010;
    assign weights2[14][59] = 16'b0000000001001011;
    assign weights2[14][60] = 16'b0000000010000010;
    assign weights2[14][61] = 16'b0000000000010110;
    assign weights2[14][62] = 16'b1111111111010000;
    assign weights2[14][63] = 16'b1111111111010110;
    assign weights2[15][0] = 16'b1111111111000101;
    assign weights2[15][1] = 16'b1111111101000011;
    assign weights2[15][2] = 16'b0000000000011101;
    assign weights2[15][3] = 16'b0000000000011110;
    assign weights2[15][4] = 16'b0000000000001000;
    assign weights2[15][5] = 16'b0000000000100000;
    assign weights2[15][6] = 16'b0000000000000000;
    assign weights2[15][7] = 16'b1111111111111010;
    assign weights2[15][8] = 16'b0000000000000011;
    assign weights2[15][9] = 16'b0000000000000001;
    assign weights2[15][10] = 16'b0000000000000101;
    assign weights2[15][11] = 16'b1111111101001010;
    assign weights2[15][12] = 16'b1111111110111111;
    assign weights2[15][13] = 16'b1111111101111001;
    assign weights2[15][14] = 16'b0000000000001001;
    assign weights2[15][15] = 16'b0000000000010101;
    assign weights2[15][16] = 16'b1111111101100111;
    assign weights2[15][17] = 16'b0000000000111001;
    assign weights2[15][18] = 16'b1111111101000101;
    assign weights2[15][19] = 16'b1111111110100110;
    assign weights2[15][20] = 16'b1111111110110111;
    assign weights2[15][21] = 16'b0000000001100000;
    assign weights2[15][22] = 16'b1111111101000111;
    assign weights2[15][23] = 16'b1111111111111111;
    assign weights2[15][24] = 16'b0000000000111001;
    assign weights2[15][25] = 16'b1111111111011010;
    assign weights2[15][26] = 16'b1111111111111010;
    assign weights2[15][27] = 16'b1111111110001101;
    assign weights2[15][28] = 16'b0000000000110000;
    assign weights2[15][29] = 16'b0000000000101111;
    assign weights2[15][30] = 16'b0000000001011101;
    assign weights2[15][31] = 16'b0000000000000010;
    assign weights2[15][32] = 16'b1111111111111100;
    assign weights2[15][33] = 16'b0000000000001011;
    assign weights2[15][34] = 16'b0000000000010011;
    assign weights2[15][35] = 16'b1111111111111001;
    assign weights2[15][36] = 16'b0000000000000101;
    assign weights2[15][37] = 16'b0000000000001010;
    assign weights2[15][38] = 16'b0000000001001010;
    assign weights2[15][39] = 16'b1111111101111100;
    assign weights2[15][40] = 16'b1111111111010111;
    assign weights2[15][41] = 16'b1111111101111011;
    assign weights2[15][42] = 16'b1111111111110010;
    assign weights2[15][43] = 16'b0000000000110101;
    assign weights2[15][44] = 16'b1111111111101101;
    assign weights2[15][45] = 16'b0000000000101000;
    assign weights2[15][46] = 16'b0000000000110011;
    assign weights2[15][47] = 16'b1111111100111100;
    assign weights2[15][48] = 16'b0000000000010010;
    assign weights2[15][49] = 16'b0000000000101010;
    assign weights2[15][50] = 16'b0000000000100110;
    assign weights2[15][51] = 16'b1111111111010110;
    assign weights2[15][52] = 16'b1111111110100000;
    assign weights2[15][53] = 16'b1111111101110010;
    assign weights2[15][54] = 16'b0000000000000000;
    assign weights2[15][55] = 16'b1111111111110110;
    assign weights2[15][56] = 16'b1111111110000011;
    assign weights2[15][57] = 16'b0000000000110110;
    assign weights2[15][58] = 16'b1111111111100010;
    assign weights2[15][59] = 16'b1111111101110001;
    assign weights2[15][60] = 16'b1111111101000010;
    assign weights2[15][61] = 16'b0000000000010111;
    assign weights2[15][62] = 16'b1111111111111000;
    assign weights2[15][63] = 16'b0000000000100110;
    assign weights2[16][0] = 16'b0000000000010010;
    assign weights2[16][1] = 16'b0000000001101100;
    assign weights2[16][2] = 16'b0000000001010010;
    assign weights2[16][3] = 16'b0000000000101111;
    assign weights2[16][4] = 16'b1111111101111010;
    assign weights2[16][5] = 16'b0000000000110000;
    assign weights2[16][6] = 16'b0000000000000000;
    assign weights2[16][7] = 16'b0000000000110101;
    assign weights2[16][8] = 16'b1111111111011110;
    assign weights2[16][9] = 16'b1111111110100000;
    assign weights2[16][10] = 16'b0000000000010011;
    assign weights2[16][11] = 16'b0000000000100110;
    assign weights2[16][12] = 16'b0000000001000110;
    assign weights2[16][13] = 16'b0000000010000000;
    assign weights2[16][14] = 16'b0000000001011011;
    assign weights2[16][15] = 16'b1111111110111011;
    assign weights2[16][16] = 16'b1111111111100110;
    assign weights2[16][17] = 16'b0000000000100110;
    assign weights2[16][18] = 16'b0000000000001111;
    assign weights2[16][19] = 16'b0000000000011011;
    assign weights2[16][20] = 16'b0000000001010001;
    assign weights2[16][21] = 16'b0000000001001010;
    assign weights2[16][22] = 16'b0000000000001100;
    assign weights2[16][23] = 16'b1111111111010000;
    assign weights2[16][24] = 16'b0000000000101011;
    assign weights2[16][25] = 16'b0000000000010110;
    assign weights2[16][26] = 16'b1111111110101011;
    assign weights2[16][27] = 16'b0000000001000101;
    assign weights2[16][28] = 16'b0000000001011111;
    assign weights2[16][29] = 16'b0000000000111000;
    assign weights2[16][30] = 16'b0000000001000111;
    assign weights2[16][31] = 16'b0000000001000110;
    assign weights2[16][32] = 16'b0000000000000101;
    assign weights2[16][33] = 16'b1111111101111101;
    assign weights2[16][34] = 16'b0000000000101000;
    assign weights2[16][35] = 16'b1111111101100101;
    assign weights2[16][36] = 16'b0000000000110111;
    assign weights2[16][37] = 16'b0000000001001111;
    assign weights2[16][38] = 16'b0000000000101001;
    assign weights2[16][39] = 16'b0000000000101001;
    assign weights2[16][40] = 16'b1111111110101111;
    assign weights2[16][41] = 16'b0000000000001101;
    assign weights2[16][42] = 16'b0000000000000100;
    assign weights2[16][43] = 16'b0000000000011101;
    assign weights2[16][44] = 16'b0000000000000111;
    assign weights2[16][45] = 16'b1111111111111111;
    assign weights2[16][46] = 16'b0000000000111010;
    assign weights2[16][47] = 16'b0000000001011000;
    assign weights2[16][48] = 16'b1111111111001101;
    assign weights2[16][49] = 16'b0000000000101001;
    assign weights2[16][50] = 16'b0000000001010101;
    assign weights2[16][51] = 16'b1111111111100001;
    assign weights2[16][52] = 16'b1111111111110000;
    assign weights2[16][53] = 16'b0000000000101000;
    assign weights2[16][54] = 16'b0000000000000000;
    assign weights2[16][55] = 16'b1111111110000110;
    assign weights2[16][56] = 16'b0000000001111001;
    assign weights2[16][57] = 16'b0000000000011011;
    assign weights2[16][58] = 16'b0000000000011001;
    assign weights2[16][59] = 16'b0000000000001011;
    assign weights2[16][60] = 16'b0000000000001101;
    assign weights2[16][61] = 16'b0000000000101000;
    assign weights2[16][62] = 16'b1111111110101110;
    assign weights2[16][63] = 16'b1111111110110011;
    assign weights2[17][0] = 16'b1111111110110110;
    assign weights2[17][1] = 16'b0000000000000100;
    assign weights2[17][2] = 16'b1111111111001011;
    assign weights2[17][3] = 16'b1111111111110100;
    assign weights2[17][4] = 16'b0000000001101111;
    assign weights2[17][5] = 16'b1111111111110100;
    assign weights2[17][6] = 16'b0000000000000000;
    assign weights2[17][7] = 16'b1111111110110110;
    assign weights2[17][8] = 16'b1111111101111100;
    assign weights2[17][9] = 16'b0000000000101110;
    assign weights2[17][10] = 16'b1111111111111010;
    assign weights2[17][11] = 16'b1111111110101110;
    assign weights2[17][12] = 16'b1111111111010010;
    assign weights2[17][13] = 16'b0000000000011011;
    assign weights2[17][14] = 16'b0000000000100000;
    assign weights2[17][15] = 16'b1111111100101001;
    assign weights2[17][16] = 16'b1111111111100110;
    assign weights2[17][17] = 16'b1111111101110110;
    assign weights2[17][18] = 16'b1111111101101110;
    assign weights2[17][19] = 16'b1111111110010100;
    assign weights2[17][20] = 16'b1111111111011001;
    assign weights2[17][21] = 16'b1111111101111110;
    assign weights2[17][22] = 16'b1111111110011110;
    assign weights2[17][23] = 16'b1111111101001111;
    assign weights2[17][24] = 16'b0000000000001010;
    assign weights2[17][25] = 16'b1111111111011011;
    assign weights2[17][26] = 16'b0000000000011110;
    assign weights2[17][27] = 16'b1111111110111000;
    assign weights2[17][28] = 16'b1111111111100111;
    assign weights2[17][29] = 16'b1111111111110111;
    assign weights2[17][30] = 16'b1111111110100111;
    assign weights2[17][31] = 16'b0000000000100000;
    assign weights2[17][32] = 16'b1111111111110011;
    assign weights2[17][33] = 16'b0000000000011100;
    assign weights2[17][34] = 16'b1111111111111001;
    assign weights2[17][35] = 16'b1111111111000000;
    assign weights2[17][36] = 16'b1111111111111100;
    assign weights2[17][37] = 16'b0000000000110100;
    assign weights2[17][38] = 16'b1111111111100001;
    assign weights2[17][39] = 16'b0000000000111000;
    assign weights2[17][40] = 16'b1111111111011001;
    assign weights2[17][41] = 16'b0000000000011000;
    assign weights2[17][42] = 16'b1111111110111101;
    assign weights2[17][43] = 16'b0000000000000101;
    assign weights2[17][44] = 16'b1111111111111100;
    assign weights2[17][45] = 16'b1111111111111110;
    assign weights2[17][46] = 16'b0000000000000000;
    assign weights2[17][47] = 16'b1111111111101101;
    assign weights2[17][48] = 16'b1111111101000000;
    assign weights2[17][49] = 16'b1111111110111010;
    assign weights2[17][50] = 16'b1111111111111010;
    assign weights2[17][51] = 16'b0000000000000100;
    assign weights2[17][52] = 16'b1111111111010000;
    assign weights2[17][53] = 16'b0000000000000111;
    assign weights2[17][54] = 16'b0000000000000000;
    assign weights2[17][55] = 16'b1111111111111000;
    assign weights2[17][56] = 16'b0000000000011000;
    assign weights2[17][57] = 16'b1111111111111100;
    assign weights2[17][58] = 16'b1111111111110101;
    assign weights2[17][59] = 16'b1111111111000101;
    assign weights2[17][60] = 16'b1111111111100010;
    assign weights2[17][61] = 16'b1111111111010011;
    assign weights2[17][62] = 16'b1111111110000000;
    assign weights2[17][63] = 16'b0000000000100000;
    assign weights2[18][0] = 16'b0000000001110100;
    assign weights2[18][1] = 16'b0000000001101101;
    assign weights2[18][2] = 16'b1111111111111010;
    assign weights2[18][3] = 16'b0000000000000011;
    assign weights2[18][4] = 16'b1111111111110110;
    assign weights2[18][5] = 16'b0000000000100111;
    assign weights2[18][6] = 16'b0000000000000000;
    assign weights2[18][7] = 16'b1111111110110001;
    assign weights2[18][8] = 16'b0000000000000101;
    assign weights2[18][9] = 16'b1111111111111100;
    assign weights2[18][10] = 16'b1111111111101100;
    assign weights2[18][11] = 16'b0000000000111110;
    assign weights2[18][12] = 16'b0000000001101011;
    assign weights2[18][13] = 16'b0000000001101110;
    assign weights2[18][14] = 16'b1111111111101011;
    assign weights2[18][15] = 16'b0000000000001001;
    assign weights2[18][16] = 16'b0000000001000101;
    assign weights2[18][17] = 16'b0000000000010101;
    assign weights2[18][18] = 16'b0000000000111110;
    assign weights2[18][19] = 16'b0000000000110001;
    assign weights2[18][20] = 16'b0000000000000011;
    assign weights2[18][21] = 16'b0000000001000110;
    assign weights2[18][22] = 16'b0000000001011101;
    assign weights2[18][23] = 16'b1111111111100001;
    assign weights2[18][24] = 16'b1111111111011110;
    assign weights2[18][25] = 16'b0000000000110000;
    assign weights2[18][26] = 16'b0000000000000011;
    assign weights2[18][27] = 16'b0000000001011011;
    assign weights2[18][28] = 16'b1111111111011010;
    assign weights2[18][29] = 16'b1111111111110001;
    assign weights2[18][30] = 16'b0000000001000011;
    assign weights2[18][31] = 16'b1111111111100110;
    assign weights2[18][32] = 16'b0000000001001010;
    assign weights2[18][33] = 16'b1111111111111101;
    assign weights2[18][34] = 16'b1111111111101110;
    assign weights2[18][35] = 16'b0000000000001110;
    assign weights2[18][36] = 16'b1111111101111011;
    assign weights2[18][37] = 16'b1111111110110111;
    assign weights2[18][38] = 16'b1111111111100110;
    assign weights2[18][39] = 16'b1111111111010000;
    assign weights2[18][40] = 16'b1111111111101001;
    assign weights2[18][41] = 16'b0000000000000101;
    assign weights2[18][42] = 16'b0000000000101001;
    assign weights2[18][43] = 16'b1111111111001011;
    assign weights2[18][44] = 16'b0000000001001001;
    assign weights2[18][45] = 16'b1111111111111101;
    assign weights2[18][46] = 16'b1111111111101101;
    assign weights2[18][47] = 16'b0000000010000101;
    assign weights2[18][48] = 16'b0000000000101010;
    assign weights2[18][49] = 16'b0000000001010110;
    assign weights2[18][50] = 16'b1111111111111010;
    assign weights2[18][51] = 16'b1111111111110111;
    assign weights2[18][52] = 16'b0000000010000011;
    assign weights2[18][53] = 16'b0000000000010101;
    assign weights2[18][54] = 16'b0000000000000000;
    assign weights2[18][55] = 16'b0000000000001111;
    assign weights2[18][56] = 16'b0000000001010000;
    assign weights2[18][57] = 16'b1111111111011110;
    assign weights2[18][58] = 16'b1111111110110111;
    assign weights2[18][59] = 16'b0000000000101110;
    assign weights2[18][60] = 16'b0000000001111101;
    assign weights2[18][61] = 16'b0000000000110001;
    assign weights2[18][62] = 16'b0000000000101101;
    assign weights2[18][63] = 16'b1111111111110000;
    assign weights2[19][0] = 16'b1111111111110011;
    assign weights2[19][1] = 16'b0000000000010100;
    assign weights2[19][2] = 16'b0000000000101110;
    assign weights2[19][3] = 16'b0000000010001001;
    assign weights2[19][4] = 16'b0000000000110101;
    assign weights2[19][5] = 16'b0000000000010011;
    assign weights2[19][6] = 16'b0000000000000000;
    assign weights2[19][7] = 16'b1111111111011000;
    assign weights2[19][8] = 16'b0000000001101001;
    assign weights2[19][9] = 16'b0000000000001001;
    assign weights2[19][10] = 16'b0000000000000010;
    assign weights2[19][11] = 16'b0000000000010011;
    assign weights2[19][12] = 16'b0000000000000011;
    assign weights2[19][13] = 16'b0000000000011010;
    assign weights2[19][14] = 16'b0000000000001001;
    assign weights2[19][15] = 16'b0000000000000010;
    assign weights2[19][16] = 16'b1111111111010100;
    assign weights2[19][17] = 16'b0000000000010101;
    assign weights2[19][18] = 16'b0000000000000010;
    assign weights2[19][19] = 16'b1111111111111011;
    assign weights2[19][20] = 16'b1111111110101011;
    assign weights2[19][21] = 16'b0000000000101110;
    assign weights2[19][22] = 16'b0000000000001111;
    assign weights2[19][23] = 16'b0000000001001110;
    assign weights2[19][24] = 16'b0000000010000101;
    assign weights2[19][25] = 16'b1111111110111110;
    assign weights2[19][26] = 16'b0000000000111010;
    assign weights2[19][27] = 16'b0000000000101001;
    assign weights2[19][28] = 16'b1111111101111101;
    assign weights2[19][29] = 16'b0000000000110011;
    assign weights2[19][30] = 16'b0000000000111010;
    assign weights2[19][31] = 16'b0000000000010000;
    assign weights2[19][32] = 16'b0000000000001000;
    assign weights2[19][33] = 16'b0000000001001000;
    assign weights2[19][34] = 16'b0000000001110110;
    assign weights2[19][35] = 16'b0000000001011101;
    assign weights2[19][36] = 16'b0000000000011010;
    assign weights2[19][37] = 16'b0000000000000111;
    assign weights2[19][38] = 16'b0000000000100101;
    assign weights2[19][39] = 16'b0000000000000100;
    assign weights2[19][40] = 16'b1111111111111101;
    assign weights2[19][41] = 16'b0000000000000000;
    assign weights2[19][42] = 16'b1111111111110000;
    assign weights2[19][43] = 16'b0000000010000101;
    assign weights2[19][44] = 16'b0000000000001000;
    assign weights2[19][45] = 16'b0000000000001111;
    assign weights2[19][46] = 16'b1111111101010011;
    assign weights2[19][47] = 16'b0000000000110010;
    assign weights2[19][48] = 16'b0000000000001100;
    assign weights2[19][49] = 16'b1111111111111100;
    assign weights2[19][50] = 16'b1111111110100101;
    assign weights2[19][51] = 16'b1111111111010011;
    assign weights2[19][52] = 16'b0000000000001010;
    assign weights2[19][53] = 16'b1111111111110110;
    assign weights2[19][54] = 16'b0000000000000000;
    assign weights2[19][55] = 16'b0000000000100111;
    assign weights2[19][56] = 16'b0000000000100110;
    assign weights2[19][57] = 16'b0000000001101101;
    assign weights2[19][58] = 16'b1111111111110011;
    assign weights2[19][59] = 16'b1111111110101111;
    assign weights2[19][60] = 16'b1111111110100110;
    assign weights2[19][61] = 16'b1111111111100000;
    assign weights2[19][62] = 16'b0000000000110000;
    assign weights2[19][63] = 16'b0000000000011011;
    assign weights2[20][0] = 16'b1111111111001000;
    assign weights2[20][1] = 16'b1111111111101111;
    assign weights2[20][2] = 16'b1111111111001011;
    assign weights2[20][3] = 16'b1111111101100011;
    assign weights2[20][4] = 16'b1111111111101011;
    assign weights2[20][5] = 16'b1111111110010111;
    assign weights2[20][6] = 16'b0000000000000000;
    assign weights2[20][7] = 16'b0000000000110110;
    assign weights2[20][8] = 16'b0000000000100110;
    assign weights2[20][9] = 16'b1111111111110011;
    assign weights2[20][10] = 16'b1111111110010001;
    assign weights2[20][11] = 16'b1111111110011110;
    assign weights2[20][12] = 16'b1111111111111011;
    assign weights2[20][13] = 16'b1111111111110011;
    assign weights2[20][14] = 16'b1111111110011001;
    assign weights2[20][15] = 16'b0000000000000010;
    assign weights2[20][16] = 16'b0000000000000000;
    assign weights2[20][17] = 16'b1111111110101110;
    assign weights2[20][18] = 16'b1111111110100001;
    assign weights2[20][19] = 16'b1111111110111011;
    assign weights2[20][20] = 16'b1111111111011110;
    assign weights2[20][21] = 16'b1111111110100001;
    assign weights2[20][22] = 16'b1111111110100000;
    assign weights2[20][23] = 16'b0000000000001111;
    assign weights2[20][24] = 16'b1111111111011011;
    assign weights2[20][25] = 16'b0000000000100101;
    assign weights2[20][26] = 16'b1111111111101100;
    assign weights2[20][27] = 16'b1111111111101111;
    assign weights2[20][28] = 16'b0000000001010101;
    assign weights2[20][29] = 16'b0000000001001011;
    assign weights2[20][30] = 16'b1111111110001110;
    assign weights2[20][31] = 16'b1111111101110010;
    assign weights2[20][32] = 16'b1111111111000000;
    assign weights2[20][33] = 16'b1111111111111000;
    assign weights2[20][34] = 16'b1111111100001011;
    assign weights2[20][35] = 16'b0000000000011010;
    assign weights2[20][36] = 16'b0000000001010000;
    assign weights2[20][37] = 16'b1111111110111010;
    assign weights2[20][38] = 16'b1111111110110010;
    assign weights2[20][39] = 16'b1111111111010010;
    assign weights2[20][40] = 16'b1111111111111000;
    assign weights2[20][41] = 16'b1111111111111111;
    assign weights2[20][42] = 16'b0000000000100110;
    assign weights2[20][43] = 16'b0000000000010111;
    assign weights2[20][44] = 16'b1111111110110100;
    assign weights2[20][45] = 16'b0000000001100001;
    assign weights2[20][46] = 16'b0000000001111001;
    assign weights2[20][47] = 16'b1111111111100110;
    assign weights2[20][48] = 16'b0000000000001100;
    assign weights2[20][49] = 16'b0000000000111000;
    assign weights2[20][50] = 16'b0000000001101111;
    assign weights2[20][51] = 16'b0000000000110100;
    assign weights2[20][52] = 16'b1111111111110001;
    assign weights2[20][53] = 16'b0000000000000011;
    assign weights2[20][54] = 16'b0000000000000000;
    assign weights2[20][55] = 16'b1111111111110001;
    assign weights2[20][56] = 16'b1111111111101011;
    assign weights2[20][57] = 16'b0000000000000101;
    assign weights2[20][58] = 16'b0000000000000001;
    assign weights2[20][59] = 16'b0000000000001010;
    assign weights2[20][60] = 16'b0000000000001100;
    assign weights2[20][61] = 16'b0000000000111010;
    assign weights2[20][62] = 16'b0000000000010001;
    assign weights2[20][63] = 16'b0000000000000011;
    assign weights2[21][0] = 16'b1111111100110100;
    assign weights2[21][1] = 16'b1111111111111011;
    assign weights2[21][2] = 16'b1111111110111111;
    assign weights2[21][3] = 16'b1111111111101011;
    assign weights2[21][4] = 16'b0000000000011100;
    assign weights2[21][5] = 16'b1111111110010111;
    assign weights2[21][6] = 16'b0000000000000000;
    assign weights2[21][7] = 16'b0000000000101011;
    assign weights2[21][8] = 16'b0000000000011110;
    assign weights2[21][9] = 16'b0000000000001100;
    assign weights2[21][10] = 16'b0000000000100111;
    assign weights2[21][11] = 16'b1111111110000100;
    assign weights2[21][12] = 16'b0000000000000110;
    assign weights2[21][13] = 16'b0000000000011100;
    assign weights2[21][14] = 16'b0000000000000001;
    assign weights2[21][15] = 16'b0000000000000101;
    assign weights2[21][16] = 16'b1111111111000100;
    assign weights2[21][17] = 16'b1111111111111000;
    assign weights2[21][18] = 16'b1111111100111111;
    assign weights2[21][19] = 16'b1111111110110011;
    assign weights2[21][20] = 16'b1111111110010111;
    assign weights2[21][21] = 16'b1111111110110011;
    assign weights2[21][22] = 16'b1111111100011111;
    assign weights2[21][23] = 16'b0000000000010101;
    assign weights2[21][24] = 16'b0000000000100010;
    assign weights2[21][25] = 16'b1111111111001110;
    assign weights2[21][26] = 16'b0000000000100110;
    assign weights2[21][27] = 16'b1111111111101001;
    assign weights2[21][28] = 16'b0000000010000111;
    assign weights2[21][29] = 16'b0000000000101001;
    assign weights2[21][30] = 16'b1111111101111000;
    assign weights2[21][31] = 16'b0000000000001101;
    assign weights2[21][32] = 16'b1111111110100100;
    assign weights2[21][33] = 16'b0000000000100000;
    assign weights2[21][34] = 16'b0000000000000001;
    assign weights2[21][35] = 16'b1111111111100010;
    assign weights2[21][36] = 16'b1111111110011101;
    assign weights2[21][37] = 16'b1111111111111010;
    assign weights2[21][38] = 16'b1111111111111010;
    assign weights2[21][39] = 16'b0000000000101110;
    assign weights2[21][40] = 16'b1111111111111010;
    assign weights2[21][41] = 16'b0000000000110101;
    assign weights2[21][42] = 16'b1111111111011111;
    assign weights2[21][43] = 16'b0000000000101110;
    assign weights2[21][44] = 16'b1111111110000110;
    assign weights2[21][45] = 16'b0000000000101011;
    assign weights2[21][46] = 16'b0000000010010001;
    assign weights2[21][47] = 16'b1111111111110001;
    assign weights2[21][48] = 16'b1111111111111001;
    assign weights2[21][49] = 16'b1111111111010100;
    assign weights2[21][50] = 16'b0000000001101001;
    assign weights2[21][51] = 16'b0000000000001011;
    assign weights2[21][52] = 16'b1111111110101100;
    assign weights2[21][53] = 16'b0000000000001110;
    assign weights2[21][54] = 16'b1111111111111111;
    assign weights2[21][55] = 16'b1111111111111101;
    assign weights2[21][56] = 16'b0000000000011000;
    assign weights2[21][57] = 16'b0000000000101010;
    assign weights2[21][58] = 16'b0000000000000101;
    assign weights2[21][59] = 16'b1111111110101101;
    assign weights2[21][60] = 16'b1111111111101101;
    assign weights2[21][61] = 16'b1111111111110100;
    assign weights2[21][62] = 16'b1111111111110000;
    assign weights2[21][63] = 16'b0000000000010011;
    assign weights2[22][0] = 16'b0000000000000100;
    assign weights2[22][1] = 16'b1111111110101110;
    assign weights2[22][2] = 16'b1111111110011011;
    assign weights2[22][3] = 16'b1111111111100000;
    assign weights2[22][4] = 16'b1111111110111001;
    assign weights2[22][5] = 16'b1111111111100011;
    assign weights2[22][6] = 16'b0000000000000000;
    assign weights2[22][7] = 16'b0000000000101010;
    assign weights2[22][8] = 16'b1111111111100110;
    assign weights2[22][9] = 16'b1111111111101010;
    assign weights2[22][10] = 16'b0000000000001110;
    assign weights2[22][11] = 16'b0000000000000000;
    assign weights2[22][12] = 16'b1111111111111011;
    assign weights2[22][13] = 16'b0000000000101010;
    assign weights2[22][14] = 16'b1111111101010111;
    assign weights2[22][15] = 16'b0000000001011101;
    assign weights2[22][16] = 16'b1111111111111000;
    assign weights2[22][17] = 16'b1111111110000100;
    assign weights2[22][18] = 16'b0000000000001010;
    assign weights2[22][19] = 16'b1111111111110100;
    assign weights2[22][20] = 16'b1111111111011011;
    assign weights2[22][21] = 16'b1111111111011011;
    assign weights2[22][22] = 16'b1111111111111111;
    assign weights2[22][23] = 16'b1111111110101000;
    assign weights2[22][24] = 16'b1111111111011011;
    assign weights2[22][25] = 16'b1111111111111101;
    assign weights2[22][26] = 16'b1111111111011000;
    assign weights2[22][27] = 16'b1111111110110100;
    assign weights2[22][28] = 16'b0000000001111111;
    assign weights2[22][29] = 16'b0000000000001110;
    assign weights2[22][30] = 16'b1111111111111000;
    assign weights2[22][31] = 16'b1111111110000110;
    assign weights2[22][32] = 16'b0000000000000111;
    assign weights2[22][33] = 16'b0000000000000100;
    assign weights2[22][34] = 16'b1111111111001101;
    assign weights2[22][35] = 16'b0000000010110110;
    assign weights2[22][36] = 16'b1111111111100001;
    assign weights2[22][37] = 16'b1111111101010011;
    assign weights2[22][38] = 16'b1111111111000001;
    assign weights2[22][39] = 16'b1111111111110010;
    assign weights2[22][40] = 16'b0000000000001111;
    assign weights2[22][41] = 16'b1111111111101111;
    assign weights2[22][42] = 16'b1111111111110011;
    assign weights2[22][43] = 16'b1111111111101010;
    assign weights2[22][44] = 16'b1111111111111111;
    assign weights2[22][45] = 16'b1111111111111100;
    assign weights2[22][46] = 16'b0000000000110001;
    assign weights2[22][47] = 16'b0000000000011010;
    assign weights2[22][48] = 16'b0000000010011110;
    assign weights2[22][49] = 16'b1111111111000011;
    assign weights2[22][50] = 16'b0000000000100000;
    assign weights2[22][51] = 16'b0000000000011000;
    assign weights2[22][52] = 16'b1111111111011000;
    assign weights2[22][53] = 16'b1111111111000011;
    assign weights2[22][54] = 16'b0000000000000000;
    assign weights2[22][55] = 16'b1111111111100001;
    assign weights2[22][56] = 16'b1111111111010100;
    assign weights2[22][57] = 16'b1111111111100110;
    assign weights2[22][58] = 16'b1111111111110101;
    assign weights2[22][59] = 16'b0000000000000101;
    assign weights2[22][60] = 16'b1111111111011111;
    assign weights2[22][61] = 16'b1111111111111001;
    assign weights2[22][62] = 16'b0000000001111100;
    assign weights2[22][63] = 16'b1111111110101111;
    assign weights2[23][0] = 16'b0000000000101011;
    assign weights2[23][1] = 16'b1111111111111001;
    assign weights2[23][2] = 16'b0000000000011010;
    assign weights2[23][3] = 16'b1111111110001010;
    assign weights2[23][4] = 16'b1111111110001111;
    assign weights2[23][5] = 16'b0000000001001100;
    assign weights2[23][6] = 16'b0000000000000000;
    assign weights2[23][7] = 16'b1111111111101010;
    assign weights2[23][8] = 16'b1111111111110101;
    assign weights2[23][9] = 16'b1111111111101100;
    assign weights2[23][10] = 16'b1111111111100100;
    assign weights2[23][11] = 16'b1111111111111011;
    assign weights2[23][12] = 16'b1111111111110110;
    assign weights2[23][13] = 16'b0000000000000000;
    assign weights2[23][14] = 16'b0000000000010100;
    assign weights2[23][15] = 16'b0000000000000011;
    assign weights2[23][16] = 16'b0000000000101110;
    assign weights2[23][17] = 16'b0000000000001100;
    assign weights2[23][18] = 16'b1111111111111001;
    assign weights2[23][19] = 16'b0000000000100110;
    assign weights2[23][20] = 16'b0000000000000111;
    assign weights2[23][21] = 16'b1111111111110001;
    assign weights2[23][22] = 16'b0000000000010011;
    assign weights2[23][23] = 16'b1111111111100010;
    assign weights2[23][24] = 16'b1111111110010101;
    assign weights2[23][25] = 16'b1111111110111111;
    assign weights2[23][26] = 16'b1111111101111011;
    assign weights2[23][27] = 16'b1111111111110001;
    assign weights2[23][28] = 16'b1111111111001111;
    assign weights2[23][29] = 16'b1111111110000011;
    assign weights2[23][30] = 16'b0000000001001001;
    assign weights2[23][31] = 16'b0000000000000110;
    assign weights2[23][32] = 16'b0000000001100111;
    assign weights2[23][33] = 16'b1111111101000110;
    assign weights2[23][34] = 16'b1111111111001100;
    assign weights2[23][35] = 16'b1111111100110101;
    assign weights2[23][36] = 16'b1111111111011110;
    assign weights2[23][37] = 16'b0000000000001000;
    assign weights2[23][38] = 16'b0000000000010100;
    assign weights2[23][39] = 16'b1111111111110111;
    assign weights2[23][40] = 16'b1111111111101111;
    assign weights2[23][41] = 16'b0000000000000010;
    assign weights2[23][42] = 16'b1111111111101011;
    assign weights2[23][43] = 16'b1111111101101110;
    assign weights2[23][44] = 16'b0000000001100110;
    assign weights2[23][45] = 16'b1111111110101010;
    assign weights2[23][46] = 16'b1111111111000101;
    assign weights2[23][47] = 16'b1111111111110001;
    assign weights2[23][48] = 16'b1111111111110101;
    assign weights2[23][49] = 16'b1111111111010011;
    assign weights2[23][50] = 16'b1111111110111001;
    assign weights2[23][51] = 16'b1111111111101000;
    assign weights2[23][52] = 16'b1111111111101010;
    assign weights2[23][53] = 16'b1111111111111111;
    assign weights2[23][54] = 16'b0000000000000000;
    assign weights2[23][55] = 16'b1111111111010010;
    assign weights2[23][56] = 16'b1111111111110111;
    assign weights2[23][57] = 16'b1111111110010000;
    assign weights2[23][58] = 16'b0000000000000000;
    assign weights2[23][59] = 16'b1111111111101101;
    assign weights2[23][60] = 16'b0000000000011100;
    assign weights2[23][61] = 16'b1111111110100101;
    assign weights2[23][62] = 16'b1111111110100110;
    assign weights2[23][63] = 16'b1111111111100101;
    assign weights2[24][0] = 16'b0000000000010100;
    assign weights2[24][1] = 16'b1111111111100111;
    assign weights2[24][2] = 16'b0000000001100001;
    assign weights2[24][3] = 16'b0000000001111001;
    assign weights2[24][4] = 16'b0000000000010001;
    assign weights2[24][5] = 16'b0000000000000111;
    assign weights2[24][6] = 16'b0000000000000000;
    assign weights2[24][7] = 16'b1111111110100001;
    assign weights2[24][8] = 16'b0000000000001101;
    assign weights2[24][9] = 16'b0000000000001111;
    assign weights2[24][10] = 16'b1111111100011011;
    assign weights2[24][11] = 16'b1111111111111101;
    assign weights2[24][12] = 16'b1111111111111000;
    assign weights2[24][13] = 16'b1111111110111001;
    assign weights2[24][14] = 16'b0000000000000101;
    assign weights2[24][15] = 16'b0000000000010001;
    assign weights2[24][16] = 16'b1111111111110111;
    assign weights2[24][17] = 16'b0000000000011110;
    assign weights2[24][18] = 16'b1111111111110000;
    assign weights2[24][19] = 16'b0000000000000100;
    assign weights2[24][20] = 16'b1111111111001000;
    assign weights2[24][21] = 16'b0000000000110010;
    assign weights2[24][22] = 16'b1111111111101110;
    assign weights2[24][23] = 16'b0000000000001000;
    assign weights2[24][24] = 16'b0000000001101011;
    assign weights2[24][25] = 16'b0000000000010110;
    assign weights2[24][26] = 16'b0000000000100110;
    assign weights2[24][27] = 16'b1111111111111101;
    assign weights2[24][28] = 16'b1111111110001101;
    assign weights2[24][29] = 16'b0000000000111101;
    assign weights2[24][30] = 16'b0000000000011111;
    assign weights2[24][31] = 16'b1111111111111000;
    assign weights2[24][32] = 16'b0000000000011111;
    assign weights2[24][33] = 16'b0000000000010101;
    assign weights2[24][34] = 16'b0000000001100110;
    assign weights2[24][35] = 16'b0000000001100111;
    assign weights2[24][36] = 16'b1111111110110101;
    assign weights2[24][37] = 16'b1111111111111000;
    assign weights2[24][38] = 16'b0000000000011110;
    assign weights2[24][39] = 16'b1111111110011100;
    assign weights2[24][40] = 16'b1111111111111011;
    assign weights2[24][41] = 16'b1111111111001000;
    assign weights2[24][42] = 16'b0000000000100111;
    assign weights2[24][43] = 16'b0000000010000001;
    assign weights2[24][44] = 16'b0000000000100001;
    assign weights2[24][45] = 16'b0000000001010000;
    assign weights2[24][46] = 16'b1111111110100000;
    assign weights2[24][47] = 16'b1111111111010111;
    assign weights2[24][48] = 16'b0000000000110111;
    assign weights2[24][49] = 16'b0000000001001100;
    assign weights2[24][50] = 16'b1111111111000101;
    assign weights2[24][51] = 16'b1111111111111011;
    assign weights2[24][52] = 16'b1111111111100110;
    assign weights2[24][53] = 16'b0000000000000011;
    assign weights2[24][54] = 16'b0000000000000000;
    assign weights2[24][55] = 16'b0000000001001001;
    assign weights2[24][56] = 16'b0000000000000000;
    assign weights2[24][57] = 16'b0000000001111111;
    assign weights2[24][58] = 16'b1111111110011110;
    assign weights2[24][59] = 16'b0000000000010100;
    assign weights2[24][60] = 16'b1111111111001001;
    assign weights2[24][61] = 16'b0000000000101101;
    assign weights2[24][62] = 16'b0000000001010011;
    assign weights2[24][63] = 16'b0000000000011110;
    assign weights2[25][0] = 16'b1111111110110000;
    assign weights2[25][1] = 16'b1111111111001111;
    assign weights2[25][2] = 16'b1111111111111111;
    assign weights2[25][3] = 16'b0000000000100110;
    assign weights2[25][4] = 16'b0000000000000100;
    assign weights2[25][5] = 16'b1111111111101101;
    assign weights2[25][6] = 16'b0000000000000000;
    assign weights2[25][7] = 16'b1111111111101010;
    assign weights2[25][8] = 16'b1111111111111110;
    assign weights2[25][9] = 16'b0000000000010010;
    assign weights2[25][10] = 16'b1111111111110110;
    assign weights2[25][11] = 16'b1111111101111111;
    assign weights2[25][12] = 16'b1111111111000011;
    assign weights2[25][13] = 16'b1111111111101000;
    assign weights2[25][14] = 16'b0000000000111100;
    assign weights2[25][15] = 16'b1111111111110101;
    assign weights2[25][16] = 16'b0000000000000110;
    assign weights2[25][17] = 16'b1111111110110100;
    assign weights2[25][18] = 16'b1111111110000010;
    assign weights2[25][19] = 16'b1111111110100010;
    assign weights2[25][20] = 16'b0000000000000100;
    assign weights2[25][21] = 16'b1111111111010010;
    assign weights2[25][22] = 16'b1111111101111100;
    assign weights2[25][23] = 16'b0000000000011100;
    assign weights2[25][24] = 16'b1111111111111111;
    assign weights2[25][25] = 16'b1111111110111100;
    assign weights2[25][26] = 16'b1111111111110110;
    assign weights2[25][27] = 16'b1111111110110001;
    assign weights2[25][28] = 16'b1111111110101111;
    assign weights2[25][29] = 16'b1111111111110010;
    assign weights2[25][30] = 16'b1111111110110101;
    assign weights2[25][31] = 16'b0000000000101100;
    assign weights2[25][32] = 16'b1111111111111000;
    assign weights2[25][33] = 16'b1111111111011011;
    assign weights2[25][34] = 16'b0000000000011110;
    assign weights2[25][35] = 16'b1111111110010111;
    assign weights2[25][36] = 16'b0000000000101000;
    assign weights2[25][37] = 16'b0000000000111011;
    assign weights2[25][38] = 16'b1111111111101111;
    assign weights2[25][39] = 16'b1111111101011110;
    assign weights2[25][40] = 16'b1111111111110011;
    assign weights2[25][41] = 16'b0000000000111010;
    assign weights2[25][42] = 16'b1111111110010111;
    assign weights2[25][43] = 16'b1111111111101001;
    assign weights2[25][44] = 16'b1111111111111001;
    assign weights2[25][45] = 16'b0000000000001011;
    assign weights2[25][46] = 16'b1111111110011000;
    assign weights2[25][47] = 16'b1111111110101010;
    assign weights2[25][48] = 16'b1111111111000110;
    assign weights2[25][49] = 16'b1111111111010111;
    assign weights2[25][50] = 16'b1111111110101001;
    assign weights2[25][51] = 16'b1111111111110010;
    assign weights2[25][52] = 16'b1111111110000011;
    assign weights2[25][53] = 16'b0000000000100101;
    assign weights2[25][54] = 16'b0000000000000000;
    assign weights2[25][55] = 16'b1111111111101001;
    assign weights2[25][56] = 16'b1111111111111100;
    assign weights2[25][57] = 16'b1111111111110011;
    assign weights2[25][58] = 16'b0000000000110001;
    assign weights2[25][59] = 16'b1111111110100101;
    assign weights2[25][60] = 16'b1111111111101001;
    assign weights2[25][61] = 16'b1111111110110110;
    assign weights2[25][62] = 16'b1111111110101011;
    assign weights2[25][63] = 16'b1111111111100010;
    assign weights2[26][0] = 16'b1111111111110010;
    assign weights2[26][1] = 16'b0000000000111001;
    assign weights2[26][2] = 16'b1111111111111111;
    assign weights2[26][3] = 16'b0000000001101111;
    assign weights2[26][4] = 16'b1111111111100000;
    assign weights2[26][5] = 16'b0000000000010011;
    assign weights2[26][6] = 16'b0000000000000000;
    assign weights2[26][7] = 16'b1111111111111001;
    assign weights2[26][8] = 16'b1111111111110111;
    assign weights2[26][9] = 16'b1111111111101100;
    assign weights2[26][10] = 16'b0000000000111111;
    assign weights2[26][11] = 16'b1111111111010001;
    assign weights2[26][12] = 16'b0000000000100101;
    assign weights2[26][13] = 16'b0000000000111000;
    assign weights2[26][14] = 16'b0000000000000111;
    assign weights2[26][15] = 16'b0000000000000011;
    assign weights2[26][16] = 16'b1111111111111100;
    assign weights2[26][17] = 16'b1111111111101000;
    assign weights2[26][18] = 16'b1111111111100100;
    assign weights2[26][19] = 16'b1111111111011011;
    assign weights2[26][20] = 16'b1111111110110101;
    assign weights2[26][21] = 16'b1111111111011000;
    assign weights2[26][22] = 16'b1111111111101101;
    assign weights2[26][23] = 16'b1111111111101001;
    assign weights2[26][24] = 16'b0000000001011101;
    assign weights2[26][25] = 16'b1111111110000001;
    assign weights2[26][26] = 16'b1111111111100011;
    assign weights2[26][27] = 16'b0000000000000010;
    assign weights2[26][28] = 16'b1111111111000100;
    assign weights2[26][29] = 16'b1111111111110100;
    assign weights2[26][30] = 16'b0000000000110010;
    assign weights2[26][31] = 16'b0000000000010001;
    assign weights2[26][32] = 16'b0000000000011110;
    assign weights2[26][33] = 16'b1111111111110100;
    assign weights2[26][34] = 16'b0000000001101110;
    assign weights2[26][35] = 16'b1111111111001001;
    assign weights2[26][36] = 16'b1111111111011000;
    assign weights2[26][37] = 16'b0000000000000100;
    assign weights2[26][38] = 16'b0000000000010111;
    assign weights2[26][39] = 16'b0000000000010011;
    assign weights2[26][40] = 16'b1111111111110110;
    assign weights2[26][41] = 16'b0000000000110011;
    assign weights2[26][42] = 16'b1111111110110001;
    assign weights2[26][43] = 16'b0000000000110010;
    assign weights2[26][44] = 16'b0000000000010111;
    assign weights2[26][45] = 16'b1111111111010000;
    assign weights2[26][46] = 16'b1111111101001011;
    assign weights2[26][47] = 16'b0000000000010111;
    assign weights2[26][48] = 16'b0000000000011011;
    assign weights2[26][49] = 16'b1111111110101101;
    assign weights2[26][50] = 16'b1111111100111110;
    assign weights2[26][51] = 16'b1111111111101100;
    assign weights2[26][52] = 16'b1111111111000000;
    assign weights2[26][53] = 16'b0000000000000000;
    assign weights2[26][54] = 16'b0000000000000000;
    assign weights2[26][55] = 16'b1111111111101110;
    assign weights2[26][56] = 16'b0000000001010100;
    assign weights2[26][57] = 16'b0000000000110010;
    assign weights2[26][58] = 16'b0000000001001011;
    assign weights2[26][59] = 16'b1111111110011001;
    assign weights2[26][60] = 16'b1111111111001011;
    assign weights2[26][61] = 16'b1111111101000110;
    assign weights2[26][62] = 16'b0000000000000101;
    assign weights2[26][63] = 16'b1111111111000000;
    assign weights2[27][0] = 16'b1111111111100110;
    assign weights2[27][1] = 16'b0000000001010010;
    assign weights2[27][2] = 16'b1111111111011000;
    assign weights2[27][3] = 16'b0000000000010011;
    assign weights2[27][4] = 16'b1111111110000001;
    assign weights2[27][5] = 16'b1111111111100101;
    assign weights2[27][6] = 16'b0000000000000000;
    assign weights2[27][7] = 16'b0000000000100111;
    assign weights2[27][8] = 16'b1111111111011110;
    assign weights2[27][9] = 16'b1111111111111011;
    assign weights2[27][10] = 16'b0000000000010011;
    assign weights2[27][11] = 16'b0000000001010100;
    assign weights2[27][12] = 16'b0000000000010101;
    assign weights2[27][13] = 16'b0000000001111001;
    assign weights2[27][14] = 16'b0000000000011110;
    assign weights2[27][15] = 16'b1111111111100110;
    assign weights2[27][16] = 16'b0000000000010001;
    assign weights2[27][17] = 16'b1111111111110111;
    assign weights2[27][18] = 16'b0000000000101100;
    assign weights2[27][19] = 16'b0000000001011101;
    assign weights2[27][20] = 16'b0000000001001101;
    assign weights2[27][21] = 16'b1111111111101000;
    assign weights2[27][22] = 16'b0000000000110010;
    assign weights2[27][23] = 16'b1111111110011000;
    assign weights2[27][24] = 16'b0000000000000111;
    assign weights2[27][25] = 16'b0000000000001010;
    assign weights2[27][26] = 16'b0000000000001101;
    assign weights2[27][27] = 16'b0000000001011010;
    assign weights2[27][28] = 16'b0000000001001111;
    assign weights2[27][29] = 16'b0000000000000011;
    assign weights2[27][30] = 16'b0000000000110100;
    assign weights2[27][31] = 16'b0000000000100011;
    assign weights2[27][32] = 16'b1111111111111100;
    assign weights2[27][33] = 16'b0000000000000001;
    assign weights2[27][34] = 16'b0000000000010011;
    assign weights2[27][35] = 16'b1111111101010000;
    assign weights2[27][36] = 16'b1111111111111111;
    assign weights2[27][37] = 16'b0000000000100100;
    assign weights2[27][38] = 16'b1111111111011101;
    assign weights2[27][39] = 16'b0000000010000110;
    assign weights2[27][40] = 16'b1111111111111110;
    assign weights2[27][41] = 16'b0000000000110111;
    assign weights2[27][42] = 16'b0000000000001000;
    assign weights2[27][43] = 16'b1111111111111101;
    assign weights2[27][44] = 16'b1111111111001010;
    assign weights2[27][45] = 16'b1111111111101100;
    assign weights2[27][46] = 16'b0000000000010111;
    assign weights2[27][47] = 16'b0000000010011101;
    assign weights2[27][48] = 16'b1111111111010111;
    assign weights2[27][49] = 16'b1111111111110110;
    assign weights2[27][50] = 16'b1111111111110111;
    assign weights2[27][51] = 16'b0000000000001101;
    assign weights2[27][52] = 16'b0000000000010101;
    assign weights2[27][53] = 16'b0000000001100001;
    assign weights2[27][54] = 16'b0000000000000000;
    assign weights2[27][55] = 16'b1111111110111100;
    assign weights2[27][56] = 16'b0000000010000010;
    assign weights2[27][57] = 16'b0000000000000101;
    assign weights2[27][58] = 16'b0000000000001010;
    assign weights2[27][59] = 16'b0000000000010100;
    assign weights2[27][60] = 16'b0000000000101010;
    assign weights2[27][61] = 16'b1111111111111010;
    assign weights2[27][62] = 16'b1111111110111111;
    assign weights2[27][63] = 16'b1111111111000110;
    assign weights2[28][0] = 16'b0000000000110101;
    assign weights2[28][1] = 16'b1111111111101110;
    assign weights2[28][2] = 16'b1111111111100111;
    assign weights2[28][3] = 16'b1111111111111011;
    assign weights2[28][4] = 16'b1111111111110010;
    assign weights2[28][5] = 16'b0000000000100100;
    assign weights2[28][6] = 16'b0000000000000000;
    assign weights2[28][7] = 16'b0000000000001101;
    assign weights2[28][8] = 16'b0000000000110101;
    assign weights2[28][9] = 16'b1111111111110110;
    assign weights2[28][10] = 16'b0000000000001000;
    assign weights2[28][11] = 16'b0000000000111111;
    assign weights2[28][12] = 16'b1111111111111011;
    assign weights2[28][13] = 16'b1111111111110000;
    assign weights2[28][14] = 16'b1111111111100100;
    assign weights2[28][15] = 16'b0000000000000101;
    assign weights2[28][16] = 16'b0000000000110000;
    assign weights2[28][17] = 16'b0000000001000001;
    assign weights2[28][18] = 16'b0000000001100111;
    assign weights2[28][19] = 16'b0000000010010101;
    assign weights2[28][20] = 16'b1111111110011100;
    assign weights2[28][21] = 16'b0000000000110111;
    assign weights2[28][22] = 16'b0000000010010010;
    assign weights2[28][23] = 16'b0000000001001010;
    assign weights2[28][24] = 16'b1111111111000111;
    assign weights2[28][25] = 16'b1111111101010010;
    assign weights2[28][26] = 16'b0000000000000001;
    assign weights2[28][27] = 16'b0000000000010001;
    assign weights2[28][28] = 16'b1111111111000101;
    assign weights2[28][29] = 16'b1111111101001110;
    assign weights2[28][30] = 16'b0000000001110101;
    assign weights2[28][31] = 16'b1111111111100001;
    assign weights2[28][32] = 16'b0000000000010000;
    assign weights2[28][33] = 16'b0000000000011101;
    assign weights2[28][34] = 16'b0000000000000101;
    assign weights2[28][35] = 16'b0000000000000000;
    assign weights2[28][36] = 16'b0000000000100111;
    assign weights2[28][37] = 16'b1111111111011100;
    assign weights2[28][38] = 16'b1111111111111101;
    assign weights2[28][39] = 16'b1111111110011110;
    assign weights2[28][40] = 16'b0000000000001011;
    assign weights2[28][41] = 16'b0000000000001111;
    assign weights2[28][42] = 16'b1111111111000011;
    assign weights2[28][43] = 16'b1111111111010111;
    assign weights2[28][44] = 16'b0000000000010000;
    assign weights2[28][45] = 16'b1111111111100010;
    assign weights2[28][46] = 16'b1111111110111001;
    assign weights2[28][47] = 16'b0000000000000010;
    assign weights2[28][48] = 16'b0000000000010000;
    assign weights2[28][49] = 16'b1111111110111110;
    assign weights2[28][50] = 16'b1111111101100000;
    assign weights2[28][51] = 16'b1111111111001101;
    assign weights2[28][52] = 16'b0000000000000101;
    assign weights2[28][53] = 16'b1111111111100010;
    assign weights2[28][54] = 16'b0000000000000000;
    assign weights2[28][55] = 16'b1111111111101001;
    assign weights2[28][56] = 16'b1111111111111100;
    assign weights2[28][57] = 16'b1111111110101000;
    assign weights2[28][58] = 16'b1111111111111100;
    assign weights2[28][59] = 16'b1111111101000010;
    assign weights2[28][60] = 16'b0000000000000111;
    assign weights2[28][61] = 16'b1111111110101011;
    assign weights2[28][62] = 16'b0000000000000100;
    assign weights2[28][63] = 16'b1111111110101011;
    assign weights2[29][0] = 16'b0000000001011111;
    assign weights2[29][1] = 16'b0000000000011101;
    assign weights2[29][2] = 16'b0000000001011000;
    assign weights2[29][3] = 16'b0000000000011011;
    assign weights2[29][4] = 16'b1111111111111111;
    assign weights2[29][5] = 16'b0000000001101101;
    assign weights2[29][6] = 16'b0000000000000000;
    assign weights2[29][7] = 16'b1111111111110101;
    assign weights2[29][8] = 16'b0000000000100011;
    assign weights2[29][9] = 16'b1111111111111011;
    assign weights2[29][10] = 16'b1111111111110010;
    assign weights2[29][11] = 16'b0000000000111010;
    assign weights2[29][12] = 16'b0000000000011010;
    assign weights2[29][13] = 16'b0000000000000100;
    assign weights2[29][14] = 16'b0000000000110110;
    assign weights2[29][15] = 16'b0000000000000000;
    assign weights2[29][16] = 16'b0000000000111000;
    assign weights2[29][17] = 16'b0000000010001110;
    assign weights2[29][18] = 16'b0000000000111110;
    assign weights2[29][19] = 16'b0000000001110011;
    assign weights2[29][20] = 16'b0000000000100100;
    assign weights2[29][21] = 16'b0000000010100100;
    assign weights2[29][22] = 16'b0000000001101010;
    assign weights2[29][23] = 16'b0000000000100100;
    assign weights2[29][24] = 16'b1111111111110100;
    assign weights2[29][25] = 16'b1111111110101101;
    assign weights2[29][26] = 16'b0000000000011010;
    assign weights2[29][27] = 16'b0000000001011000;
    assign weights2[29][28] = 16'b1111111111101001;
    assign weights2[29][29] = 16'b1111111110010000;
    assign weights2[29][30] = 16'b0000000010110100;
    assign weights2[29][31] = 16'b0000000000110011;
    assign weights2[29][32] = 16'b0000000000110010;
    assign weights2[29][33] = 16'b0000000000100110;
    assign weights2[29][34] = 16'b0000000000100010;
    assign weights2[29][35] = 16'b0000000000101010;
    assign weights2[29][36] = 16'b1111111111010011;
    assign weights2[29][37] = 16'b0000000000101100;
    assign weights2[29][38] = 16'b0000000000101110;
    assign weights2[29][39] = 16'b1111111111100100;
    assign weights2[29][40] = 16'b1111111111011011;
    assign weights2[29][41] = 16'b1111111111101111;
    assign weights2[29][42] = 16'b1111111111111000;
    assign weights2[29][43] = 16'b1111111111010110;
    assign weights2[29][44] = 16'b0000000000110111;
    assign weights2[29][45] = 16'b1111111101110100;
    assign weights2[29][46] = 16'b1111111111011011;
    assign weights2[29][47] = 16'b0000000000101101;
    assign weights2[29][48] = 16'b0000000000001010;
    assign weights2[29][49] = 16'b0000000000101001;
    assign weights2[29][50] = 16'b1111111110101111;
    assign weights2[29][51] = 16'b1111111111000000;
    assign weights2[29][52] = 16'b0000000000110000;
    assign weights2[29][53] = 16'b1111111111111111;
    assign weights2[29][54] = 16'b0000000000000000;
    assign weights2[29][55] = 16'b0000000000000010;
    assign weights2[29][56] = 16'b0000000000011010;
    assign weights2[29][57] = 16'b1111111111010001;
    assign weights2[29][58] = 16'b1111111111100011;
    assign weights2[29][59] = 16'b1111111110101111;
    assign weights2[29][60] = 16'b0000000000011101;
    assign weights2[29][61] = 16'b1111111111011000;
    assign weights2[29][62] = 16'b0000000000001010;
    assign weights2[29][63] = 16'b0000000000000001;
    assign weights2[30][0] = 16'b1111111111111001;
    assign weights2[30][1] = 16'b0000000010111100;
    assign weights2[30][2] = 16'b0000000001011010;
    assign weights2[30][3] = 16'b0000000000001101;
    assign weights2[30][4] = 16'b1111111111100011;
    assign weights2[30][5] = 16'b0000000000011111;
    assign weights2[30][6] = 16'b0000000000000000;
    assign weights2[30][7] = 16'b0000000001110001;
    assign weights2[30][8] = 16'b0000000000111010;
    assign weights2[30][9] = 16'b1111111111101101;
    assign weights2[30][10] = 16'b0000000000111011;
    assign weights2[30][11] = 16'b0000000000010100;
    assign weights2[30][12] = 16'b0000000010101101;
    assign weights2[30][13] = 16'b0000000010001001;
    assign weights2[30][14] = 16'b1111111111111010;
    assign weights2[30][15] = 16'b1111111111111010;
    assign weights2[30][16] = 16'b1111111111010001;
    assign weights2[30][17] = 16'b0000000001001110;
    assign weights2[30][18] = 16'b1111111111110110;
    assign weights2[30][19] = 16'b1111111111100011;
    assign weights2[30][20] = 16'b1111111110001100;
    assign weights2[30][21] = 16'b0000000001010011;
    assign weights2[30][22] = 16'b0000000000000001;
    assign weights2[30][23] = 16'b0000000000000111;
    assign weights2[30][24] = 16'b0000000000010110;
    assign weights2[30][25] = 16'b0000000000001011;
    assign weights2[30][26] = 16'b1111111111111110;
    assign weights2[30][27] = 16'b0000000000110101;
    assign weights2[30][28] = 16'b0000000010001001;
    assign weights2[30][29] = 16'b0000000001001000;
    assign weights2[30][30] = 16'b0000000001000010;
    assign weights2[30][31] = 16'b1111111111011110;
    assign weights2[30][32] = 16'b1111111111010111;
    assign weights2[30][33] = 16'b1111111111111001;
    assign weights2[30][34] = 16'b0000000000000010;
    assign weights2[30][35] = 16'b0000000001000001;
    assign weights2[30][36] = 16'b0000000001100101;
    assign weights2[30][37] = 16'b1111111111101101;
    assign weights2[30][38] = 16'b0000000000011101;
    assign weights2[30][39] = 16'b1111111111010010;
    assign weights2[30][40] = 16'b1111111111001001;
    assign weights2[30][41] = 16'b1111111111101000;
    assign weights2[30][42] = 16'b0000000000000101;
    assign weights2[30][43] = 16'b0000000000011001;
    assign weights2[30][44] = 16'b1111111111101010;
    assign weights2[30][45] = 16'b0000000000011111;
    assign weights2[30][46] = 16'b0000000010010010;
    assign weights2[30][47] = 16'b0000000001010010;
    assign weights2[30][48] = 16'b0000000000100101;
    assign weights2[30][49] = 16'b0000000000101011;
    assign weights2[30][50] = 16'b0000000010011110;
    assign weights2[30][51] = 16'b1111111111011000;
    assign weights2[30][52] = 16'b1111111111100100;
    assign weights2[30][53] = 16'b1111111111001101;
    assign weights2[30][54] = 16'b0000000000000000;
    assign weights2[30][55] = 16'b1111111111110000;
    assign weights2[30][56] = 16'b1111111111111100;
    assign weights2[30][57] = 16'b0000000000011110;
    assign weights2[30][58] = 16'b1111111111110001;
    assign weights2[30][59] = 16'b1111111111100111;
    assign weights2[30][60] = 16'b1111111111101110;
    assign weights2[30][61] = 16'b0000000000011010;
    assign weights2[30][62] = 16'b0000000001010100;
    assign weights2[30][63] = 16'b0000000000000101;
    assign weights2[31][0] = 16'b0000000000001001;
    assign weights2[31][1] = 16'b1111111101101111;
    assign weights2[31][2] = 16'b0000000000100110;
    assign weights2[31][3] = 16'b0000000000010011;
    assign weights2[31][4] = 16'b1111111110111101;
    assign weights2[31][5] = 16'b0000000000101110;
    assign weights2[31][6] = 16'b0000000000000000;
    assign weights2[31][7] = 16'b1111111111100110;
    assign weights2[31][8] = 16'b0000000000100111;
    assign weights2[31][9] = 16'b1111111110110100;
    assign weights2[31][10] = 16'b0000000000000110;
    assign weights2[31][11] = 16'b1111111101001001;
    assign weights2[31][12] = 16'b1111111111111111;
    assign weights2[31][13] = 16'b1111111110100000;
    assign weights2[31][14] = 16'b0000000000011111;
    assign weights2[31][15] = 16'b1111111111111001;
    assign weights2[31][16] = 16'b1111111110011111;
    assign weights2[31][17] = 16'b0000000000100001;
    assign weights2[31][18] = 16'b1111111110000101;
    assign weights2[31][19] = 16'b1111111111000100;
    assign weights2[31][20] = 16'b1111111111011100;
    assign weights2[31][21] = 16'b0000000000111101;
    assign weights2[31][22] = 16'b1111111110101100;
    assign weights2[31][23] = 16'b0000000000011001;
    assign weights2[31][24] = 16'b0000000000100100;
    assign weights2[31][25] = 16'b0000000000110101;
    assign weights2[31][26] = 16'b1111111110100101;
    assign weights2[31][27] = 16'b1111111110011010;
    assign weights2[31][28] = 16'b0000000000001001;
    assign weights2[31][29] = 16'b0000000000111001;
    assign weights2[31][30] = 16'b0000000000111100;
    assign weights2[31][31] = 16'b0000000000010010;
    assign weights2[31][32] = 16'b0000000000011111;
    assign weights2[31][33] = 16'b1111111111000101;
    assign weights2[31][34] = 16'b0000000000010110;
    assign weights2[31][35] = 16'b0000000000110101;
    assign weights2[31][36] = 16'b0000000000000100;
    assign weights2[31][37] = 16'b0000000000010100;
    assign weights2[31][38] = 16'b0000000000101101;
    assign weights2[31][39] = 16'b1111111101101100;
    assign weights2[31][40] = 16'b1111111101110011;
    assign weights2[31][41] = 16'b1111111101001110;
    assign weights2[31][42] = 16'b0000000000001001;
    assign weights2[31][43] = 16'b0000000000011111;
    assign weights2[31][44] = 16'b0000000000101110;
    assign weights2[31][45] = 16'b0000000000111001;
    assign weights2[31][46] = 16'b1111111111101100;
    assign weights2[31][47] = 16'b1111111101010111;
    assign weights2[31][48] = 16'b1111111111101110;
    assign weights2[31][49] = 16'b0000000000110110;
    assign weights2[31][50] = 16'b0000000000100100;
    assign weights2[31][51] = 16'b1111111111010001;
    assign weights2[31][52] = 16'b1111111111010100;
    assign weights2[31][53] = 16'b1111111110000111;
    assign weights2[31][54] = 16'b0000000000000000;
    assign weights2[31][55] = 16'b1111111110111010;
    assign weights2[31][56] = 16'b1111111110011101;
    assign weights2[31][57] = 16'b0000000000100101;
    assign weights2[31][58] = 16'b0000000000000111;
    assign weights2[31][59] = 16'b1111111110101100;
    assign weights2[31][60] = 16'b1111111110001000;
    assign weights2[31][61] = 16'b0000000000111001;
    assign weights2[31][62] = 16'b1111111111100111;
    assign weights2[31][63] = 16'b1111111111010000;
    assign biases2[0] = 16'b0000000010000011;
    assign biases2[1] = 16'b0000000001110011;
    assign biases2[2] = 16'b0000000010001011;
    assign biases2[3] = 16'b0000000011010100;
    assign biases2[4] = 16'b0000000010101100;
    assign biases2[5] = 16'b0000000000111101;
    assign biases2[6] = 16'b0000000011111100;
    assign biases2[7] = 16'b0000000011110111;
    assign biases2[8] = 16'b0000000010110001;
    assign biases2[9] = 16'b1111111110001000;
    assign biases2[10] = 16'b0000000000100001;
    assign biases2[11] = 16'b0000000100101101;
    assign biases2[12] = 16'b1111111101101000;
    assign biases2[13] = 16'b0000000110110010;
    assign biases2[14] = 16'b0000000100000101;
    assign biases2[15] = 16'b0000000010011100;
    assign biases2[16] = 16'b0000000000010100;
    assign biases2[17] = 16'b0000000100100011;
    assign biases2[18] = 16'b1111111101111111;
    assign biases2[19] = 16'b1111111110010101;
    assign biases2[20] = 16'b0000000011101001;
    assign biases2[21] = 16'b0000000010101111;
    assign biases2[22] = 16'b0000000011010101;
    assign biases2[23] = 16'b0000000100011011;
    assign biases2[24] = 16'b1111111111010110;
    assign biases2[25] = 16'b0000000101010010;
    assign biases2[26] = 16'b0000000010000000;
    assign biases2[27] = 16'b0000000000000111;
    assign biases2[28] = 16'b0000000001011011;
    assign biases2[29] = 16'b1111111100101010;
    assign biases2[30] = 16'b1111111110011101;
    assign biases2[31] = 16'b0000000001110000;
    assign weights3[0][0] = 16'b0000000001111011;
    assign weights3[0][1] = 16'b1111111110001010;
    assign weights3[0][2] = 16'b0000000000111111;
    assign weights3[0][3] = 16'b0000000010110101;
    assign weights3[0][4] = 16'b1111111101101011;
    assign weights3[0][5] = 16'b0000000000110001;
    assign weights3[0][6] = 16'b0000000010011111;
    assign weights3[0][7] = 16'b0000000000000000;
    assign weights3[0][8] = 16'b1111111101101001;
    assign weights3[0][9] = 16'b1111111101101000;
    assign weights3[0][10] = 16'b1111111101111110;
    assign weights3[0][11] = 16'b1111111111101110;
    assign weights3[0][12] = 16'b0000000000010110;
    assign weights3[0][13] = 16'b0000000000100100;
    assign weights3[0][14] = 16'b0000000001100010;
    assign weights3[0][15] = 16'b1111111111011101;
    assign weights3[0][16] = 16'b1111111101001100;
    assign weights3[0][17] = 16'b1111111110100000;
    assign weights3[0][18] = 16'b0000000001001101;
    assign weights3[0][19] = 16'b1111111110101111;
    assign weights3[0][20] = 16'b0000000001000001;
    assign weights3[0][21] = 16'b1111111101101101;
    assign weights3[0][22] = 16'b0000000001000000;
    assign weights3[0][23] = 16'b0000000000011101;
    assign weights3[0][24] = 16'b0000000001000100;
    assign weights3[0][25] = 16'b1111111110010100;
    assign weights3[0][26] = 16'b1111111110100000;
    assign weights3[0][27] = 16'b1111111110101011;
    assign weights3[0][28] = 16'b1111111110101010;
    assign weights3[0][29] = 16'b1111111110101010;
    assign weights3[0][30] = 16'b1111111101111001;
    assign weights3[0][31] = 16'b0000000000011010;
    assign weights3[1][0] = 16'b1111111110000100;
    assign weights3[1][1] = 16'b1111111110000010;
    assign weights3[1][2] = 16'b0000000000100111;
    assign weights3[1][3] = 16'b1111111110100111;
    assign weights3[1][4] = 16'b0000000000110110;
    assign weights3[1][5] = 16'b0000000000000110;
    assign weights3[1][6] = 16'b1111111100000000;
    assign weights3[1][7] = 16'b0000000001110000;
    assign weights3[1][8] = 16'b1111111111100011;
    assign weights3[1][9] = 16'b0000000000000011;
    assign weights3[1][10] = 16'b1111111111011101;
    assign weights3[1][11] = 16'b1111111110101101;
    assign weights3[1][12] = 16'b0000000001001011;
    assign weights3[1][13] = 16'b0000000001101011;
    assign weights3[1][14] = 16'b1111111101101010;
    assign weights3[1][15] = 16'b0000000010000111;
    assign weights3[1][16] = 16'b0000000001001011;
    assign weights3[1][17] = 16'b1111111100100011;
    assign weights3[1][18] = 16'b0000000000000101;
    assign weights3[1][19] = 16'b0000000000110001;
    assign weights3[1][20] = 16'b0000000000011111;
    assign weights3[1][21] = 16'b1111111101011101;
    assign weights3[1][22] = 16'b1111111101111001;
    assign weights3[1][23] = 16'b0000000000010100;
    assign weights3[1][24] = 16'b0000000000110110;
    assign weights3[1][25] = 16'b0000000001010010;
    assign weights3[1][26] = 16'b0000000001000001;
    assign weights3[1][27] = 16'b1111111101101010;
    assign weights3[1][28] = 16'b0000000000001001;
    assign weights3[1][29] = 16'b0000000001001101;
    assign weights3[1][30] = 16'b0000000001011100;
    assign weights3[1][31] = 16'b0000000011000111;
    assign weights3[2][0] = 16'b0000000001001011;
    assign weights3[2][1] = 16'b1111111110001110;
    assign weights3[2][2] = 16'b0000000000101000;
    assign weights3[2][3] = 16'b1111111101101011;
    assign weights3[2][4] = 16'b1111111110011001;
    assign weights3[2][5] = 16'b0000000000011101;
    assign weights3[2][6] = 16'b1111111111011101;
    assign weights3[2][7] = 16'b1111111111010010;
    assign weights3[2][8] = 16'b1111111110101100;
    assign weights3[2][9] = 16'b0000000000110010;
    assign weights3[2][10] = 16'b0000000000110101;
    assign weights3[2][11] = 16'b0000000001111000;
    assign weights3[2][12] = 16'b0000000000001100;
    assign weights3[2][13] = 16'b1111111101011010;
    assign weights3[2][14] = 16'b1111111110111110;
    assign weights3[2][15] = 16'b1111111101111110;
    assign weights3[2][16] = 16'b1111111110100000;
    assign weights3[2][17] = 16'b0000000000010111;
    assign weights3[2][18] = 16'b0000000001000000;
    assign weights3[2][19] = 16'b0000000000111000;
    assign weights3[2][20] = 16'b1111111110001110;
    assign weights3[2][21] = 16'b1111111110110010;
    assign weights3[2][22] = 16'b1111111111111100;
    assign weights3[2][23] = 16'b0000000000000001;
    assign weights3[2][24] = 16'b0000000000110110;
    assign weights3[2][25] = 16'b1111111101011101;
    assign weights3[2][26] = 16'b1111111101100110;
    assign weights3[2][27] = 16'b1111111111111010;
    assign weights3[2][28] = 16'b0000000001001101;
    assign weights3[2][29] = 16'b0000000001010110;
    assign weights3[2][30] = 16'b0000000000000101;
    assign weights3[2][31] = 16'b1111111110011001;
    assign weights3[3][0] = 16'b1111111111000010;
    assign weights3[3][1] = 16'b0000000001000101;
    assign weights3[3][2] = 16'b0000000000110010;
    assign weights3[3][3] = 16'b1111111101111100;
    assign weights3[3][4] = 16'b1111111110110110;
    assign weights3[3][5] = 16'b1111111110101100;
    assign weights3[3][6] = 16'b1111111110111011;
    assign weights3[3][7] = 16'b1111111110111111;
    assign weights3[3][8] = 16'b0000000000110011;
    assign weights3[3][9] = 16'b1111111110111101;
    assign weights3[3][10] = 16'b0000000000110000;
    assign weights3[3][11] = 16'b1111111111011001;
    assign weights3[3][12] = 16'b1111111110110100;
    assign weights3[3][13] = 16'b1111111101101001;
    assign weights3[3][14] = 16'b1111111111011100;
    assign weights3[3][15] = 16'b1111111101100011;
    assign weights3[3][16] = 16'b0000000001000110;
    assign weights3[3][17] = 16'b1111111110101010;
    assign weights3[3][18] = 16'b0000000000111111;
    assign weights3[3][19] = 16'b0000000000010011;
    assign weights3[3][20] = 16'b1111111101101111;
    assign weights3[3][21] = 16'b1111111110011111;
    assign weights3[3][22] = 16'b0000000000110110;
    assign weights3[3][23] = 16'b0000000001000100;
    assign weights3[3][24] = 16'b1111111111001011;
    assign weights3[3][25] = 16'b1111111110101001;
    assign weights3[3][26] = 16'b0000000000111001;
    assign weights3[3][27] = 16'b0000000000110011;
    assign weights3[3][28] = 16'b0000000001001011;
    assign weights3[3][29] = 16'b0000000001000011;
    assign weights3[3][30] = 16'b0000000000100111;
    assign weights3[3][31] = 16'b1111111110011101;
    assign weights3[4][0] = 16'b1111111111011101;
    assign weights3[4][1] = 16'b1111111110101010;
    assign weights3[4][2] = 16'b1111111100011000;
    assign weights3[4][3] = 16'b1111111111101100;
    assign weights3[4][4] = 16'b0000000001010011;
    assign weights3[4][5] = 16'b0000000001000001;
    assign weights3[4][6] = 16'b0000000001100101;
    assign weights3[4][7] = 16'b1111111110010100;
    assign weights3[4][8] = 16'b1111111110000100;
    assign weights3[4][9] = 16'b0000000000011110;
    assign weights3[4][10] = 16'b1111111110100101;
    assign weights3[4][11] = 16'b1111111111010110;
    assign weights3[4][12] = 16'b0000000001000001;
    assign weights3[4][13] = 16'b0000000000111000;
    assign weights3[4][14] = 16'b1111111101111000;
    assign weights3[4][15] = 16'b1111111111111101;
    assign weights3[4][16] = 16'b0000000000011001;
    assign weights3[4][17] = 16'b0000000001101110;
    assign weights3[4][18] = 16'b1111111101110110;
    assign weights3[4][19] = 16'b0000000000111010;
    assign weights3[4][20] = 16'b1111111111010010;
    assign weights3[4][21] = 16'b0000000001000001;
    assign weights3[4][22] = 16'b1111111110001111;
    assign weights3[4][23] = 16'b1111111110001011;
    assign weights3[4][24] = 16'b0000000000111001;
    assign weights3[4][25] = 16'b0000000001011011;
    assign weights3[4][26] = 16'b0000000001001110;
    assign weights3[4][27] = 16'b0000000000111000;
    assign weights3[4][28] = 16'b1111111110000110;
    assign weights3[4][29] = 16'b1111111110100111;
    assign weights3[4][30] = 16'b1111111101011111;
    assign weights3[4][31] = 16'b1111111101011101;
    assign weights3[5][0] = 16'b1111111110111101;
    assign weights3[5][1] = 16'b0000000001001010;
    assign weights3[5][2] = 16'b1111111111111110;
    assign weights3[5][3] = 16'b1111111110000100;
    assign weights3[5][4] = 16'b1111111110100011;
    assign weights3[5][5] = 16'b1111111110111010;
    assign weights3[5][6] = 16'b1111111110110010;
    assign weights3[5][7] = 16'b1111111111010110;
    assign weights3[5][8] = 16'b0000000001010100;
    assign weights3[5][9] = 16'b1111111111110111;
    assign weights3[5][10] = 16'b0000000000101111;
    assign weights3[5][11] = 16'b1111111110110110;
    assign weights3[5][12] = 16'b0000000001000101;
    assign weights3[5][13] = 16'b1111111101110110;
    assign weights3[5][14] = 16'b0000000000111111;
    assign weights3[5][15] = 16'b1111111111000110;
    assign weights3[5][16] = 16'b0000000000111111;
    assign weights3[5][17] = 16'b1111111110101111;
    assign weights3[5][18] = 16'b0000000000101011;
    assign weights3[5][19] = 16'b1111111111100001;
    assign weights3[5][20] = 16'b0000000001010010;
    assign weights3[5][21] = 16'b0000000001001001;
    assign weights3[5][22] = 16'b0000000000110001;
    assign weights3[5][23] = 16'b1111111101000100;
    assign weights3[5][24] = 16'b1111111110101101;
    assign weights3[5][25] = 16'b1111111110100000;
    assign weights3[5][26] = 16'b1111111111001011;
    assign weights3[5][27] = 16'b0000000000101111;
    assign weights3[5][28] = 16'b1111111110101010;
    assign weights3[5][29] = 16'b1111111110011000;
    assign weights3[5][30] = 16'b0000000000110100;
    assign weights3[5][31] = 16'b1111111110110111;
    assign weights3[6][0] = 16'b0000000001011101;
    assign weights3[6][1] = 16'b1111111111110000;
    assign weights3[6][2] = 16'b1111111110011011;
    assign weights3[6][3] = 16'b0000000001110011;
    assign weights3[6][4] = 16'b1111111110001110;
    assign weights3[6][5] = 16'b1111111100110001;
    assign weights3[6][6] = 16'b0000000010000001;
    assign weights3[6][7] = 16'b1111111110001011;
    assign weights3[6][8] = 16'b0000000001001001;
    assign weights3[6][9] = 16'b0000000000101100;
    assign weights3[6][10] = 16'b1111111100100100;
    assign weights3[6][11] = 16'b0000000001001001;
    assign weights3[6][12] = 16'b0000000001000001;
    assign weights3[6][13] = 16'b1111111111011100;
    assign weights3[6][14] = 16'b1111111110111110;
    assign weights3[6][15] = 16'b0000000010101000;
    assign weights3[6][16] = 16'b1111111101111100;
    assign weights3[6][17] = 16'b0000000000111101;
    assign weights3[6][18] = 16'b1111111101001111;
    assign weights3[6][19] = 16'b0000000000101110;
    assign weights3[6][20] = 16'b0000000001100010;
    assign weights3[6][21] = 16'b0000000001011111;
    assign weights3[6][22] = 16'b0000000000101001;
    assign weights3[6][23] = 16'b1111111100011010;
    assign weights3[6][24] = 16'b0000000000110000;
    assign weights3[6][25] = 16'b1111111110000110;
    assign weights3[6][26] = 16'b1111111111101001;
    assign weights3[6][27] = 16'b1111111101010101;
    assign weights3[6][28] = 16'b1111111110001001;
    assign weights3[6][29] = 16'b1111111111001101;
    assign weights3[6][30] = 16'b0000000000101111;
    assign weights3[6][31] = 16'b0000000000010001;
    assign weights3[7][0] = 16'b1111111101110011;
    assign weights3[7][1] = 16'b1111111101100001;
    assign weights3[7][2] = 16'b0000000000110011;
    assign weights3[7][3] = 16'b1111111110101111;
    assign weights3[7][4] = 16'b0000000001100100;
    assign weights3[7][5] = 16'b0000000001001111;
    assign weights3[7][6] = 16'b1111111110000001;
    assign weights3[7][7] = 16'b0000000010000010;
    assign weights3[7][8] = 16'b1111111101111111;
    assign weights3[7][9] = 16'b0000000000101100;
    assign weights3[7][10] = 16'b0000000000101111;
    assign weights3[7][11] = 16'b1111111111011100;
    assign weights3[7][12] = 16'b0000000001000000;
    assign weights3[7][13] = 16'b1111111110101011;
    assign weights3[7][14] = 16'b0000000001010000;
    assign weights3[7][15] = 16'b1111111100111100;
    assign weights3[7][16] = 16'b0000000001010101;
    assign weights3[7][17] = 16'b1111111111010111;
    assign weights3[7][18] = 16'b0000000000111000;
    assign weights3[7][19] = 16'b1111111110101111;
    assign weights3[7][20] = 16'b1111111110001100;
    assign weights3[7][21] = 16'b1111111111010000;
    assign weights3[7][22] = 16'b1111111100111111;
    assign weights3[7][23] = 16'b0000000001000110;
    assign weights3[7][24] = 16'b1111111110101000;
    assign weights3[7][25] = 16'b1111111111001000;
    assign weights3[7][26] = 16'b1111111110001110;
    assign weights3[7][27] = 16'b0000000001000010;
    assign weights3[7][28] = 16'b0000000000110010;
    assign weights3[7][29] = 16'b0000000001001111;
    assign weights3[7][30] = 16'b1111111110001111;
    assign weights3[7][31] = 16'b1111111110111111;
    assign weights3[8][0] = 16'b1111111111101110;
    assign weights3[8][1] = 16'b0000000000100110;
    assign weights3[8][2] = 16'b0000000000101110;
    assign weights3[8][3] = 16'b1111111101100001;
    assign weights3[8][4] = 16'b1111111110011111;
    assign weights3[8][5] = 16'b1111111110100000;
    assign weights3[8][6] = 16'b1111111101111011;
    assign weights3[8][7] = 16'b0000000010010011;
    assign weights3[8][8] = 16'b0000000001000011;
    assign weights3[8][9] = 16'b1111111110101001;
    assign weights3[8][10] = 16'b1111111111111100;
    assign weights3[8][11] = 16'b0000000001101101;
    assign weights3[8][12] = 16'b1111111111010001;
    assign weights3[8][13] = 16'b0000000001100000;
    assign weights3[8][14] = 16'b0000000000111011;
    assign weights3[8][15] = 16'b1111111111001011;
    assign weights3[8][16] = 16'b1111111110111110;
    assign weights3[8][17] = 16'b1111111101110000;
    assign weights3[8][18] = 16'b1111111111000101;
    assign weights3[8][19] = 16'b1111111111100011;
    assign weights3[8][20] = 16'b0000000000111010;
    assign weights3[8][21] = 16'b0000000000011101;
    assign weights3[8][22] = 16'b0000000000010110;
    assign weights3[8][23] = 16'b0000000000100110;
    assign weights3[8][24] = 16'b1111111111001010;
    assign weights3[8][25] = 16'b0000000001101000;
    assign weights3[8][26] = 16'b0000000000010010;
    assign weights3[8][27] = 16'b1111111111001110;
    assign weights3[8][28] = 16'b0000000000110011;
    assign weights3[8][29] = 16'b1111111111001011;
    assign weights3[8][30] = 16'b1111111111001111;
    assign weights3[8][31] = 16'b0000000000010110;
    assign weights3[9][0] = 16'b1111111111101101;
    assign weights3[9][1] = 16'b0000000000111111;
    assign weights3[9][2] = 16'b1111111110010010;
    assign weights3[9][3] = 16'b0000000000001110;
    assign weights3[9][4] = 16'b0000000001010011;
    assign weights3[9][5] = 16'b0000000001000001;
    assign weights3[9][6] = 16'b0000000001101111;
    assign weights3[9][7] = 16'b1111111111001111;
    assign weights3[9][8] = 16'b1111111111001010;
    assign weights3[9][9] = 16'b1111111111001000;
    assign weights3[9][10] = 16'b0000000000100000;
    assign weights3[9][11] = 16'b1111111111000110;
    assign weights3[9][12] = 16'b1111111101110110;
    assign weights3[9][13] = 16'b0000000000010011;
    assign weights3[9][14] = 16'b0000000001001001;
    assign weights3[9][15] = 16'b1111111110001010;
    assign weights3[9][16] = 16'b0000000000111101;
    assign weights3[9][17] = 16'b0000000001110010;
    assign weights3[9][18] = 16'b0000000000000110;
    assign weights3[9][19] = 16'b1111111101100110;
    assign weights3[9][20] = 16'b1111111110111001;
    assign weights3[9][21] = 16'b0000000000001010;
    assign weights3[9][22] = 16'b1111111110000010;
    assign weights3[9][23] = 16'b0000000001100010;
    assign weights3[9][24] = 16'b1111111101110010;
    assign weights3[9][25] = 16'b0000000001000110;
    assign weights3[9][26] = 16'b0000000000011011;
    assign weights3[9][27] = 16'b0000000000101011;
    assign weights3[9][28] = 16'b1111111101011110;
    assign weights3[9][29] = 16'b1111111111011111;
    assign weights3[9][30] = 16'b1111111111011101;
    assign weights3[9][31] = 16'b1111111101111110;
    assign biases3[0] = 16'b0000000000000100;
    assign biases3[1] = 16'b1111111011110110;
    assign biases3[2] = 16'b0000000000011001;
    assign biases3[3] = 16'b1111111111110100;
    assign biases3[4] = 16'b0000000001000000;
    assign biases3[5] = 16'b0000000000110111;
    assign biases3[6] = 16'b1111111110001101;
    assign biases3[7] = 16'b1111111101100110;
    assign biases3[8] = 16'b0000000011001010;
    assign biases3[9] = 16'b0000000010001111;


endmodule
