//////////////////////////////////////////////////////////////////////////////////
// AXI4 Lite Slave Example
// By:
//        Ali Jahanian
// 
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module axi4_lite_slave #(
    parameter ADDRESS = 32,
    parameter DATA_WIDTH = 32
    )
    (
        // Global Signals
        input                           ACLK, // # of used = 1
        input                           ARESETN, // # of used = 1

        // Read Address Channel INPUTS
        input           [ADDRESS-1:0]   S_ARADDR, // # of used = 4
        input                           S_ARVALID, // # of used = 2

        // Read Data Channel INPUTS
        input                           S_RREADY, // # of used = 1

        // Write Address Channel INPUTS
        /* verilator lint_off UNUSED */
        input           [ADDRESS-1:0]   S_AWADDR, // # of used = 4
        input                           S_AWVALID, // # of used = 2

        // Write Data  Channel INPUTS
        input          [DATA_WIDTH-1:0] S_WDATA, // # of used = 2
        input          [3:0]            S_WSTRB, // # of used = 0
        input                           S_WVALID, // # of used = 1

        // Write Response Channel INPUTS
        input                           S_BREADY, // # of used = 1

        // Read Address Channel OUTPUTS
        output                     S_ARREADY, // # of used = 2

        // Read Data Channel OUTPUTS
        output [DATA_WIDTH-1:0]    S_RDATA, // # of used = 1
        output          [1:0]      S_RRESP, // # of used = 1
        output                     S_RVALID, // # of used = 2

        // Write Address Channel OUTPUTS
        output                     S_AWREADY, // # of used = 2
        output                     S_WREADY, // # of used = 2
        
        // Write Response Channel OUTPUTS
        output          [1:0]      S_BRESP, // # of used = 1
        output                     S_BVALID // # of used = 2
    );

    localparam REG_NUM       = 32;
    localparam IDLE          = 0;
    localparam WRITE_CHANNEL = 1;
    localparam WRESP_CHANNEL = 2;
    localparam RADDR_CHANNEL = 3;
    localparam RDATA_CHANNEL = 4;
    localparam MY_STATE      = 5;

    reg start;
    wire clk;
    reg rst;
    reg [783:0] in_features;
    reg [783:0] not_reversed_in_features;
    wire [3:0] prediction;
    wire done;

    NeuralNetwork my_NeuralNetwork (clk, rst, start, in_features, prediction, done);

    assign clk = ACLK;
   
    reg  [2:0] state, next_state;
    reg  [ADDRESS-1:0] read_addr;
    wire [ADDRESS-1:0] S_ARADDR_T;
    wire [ADDRESS-1:0] S_AWADDR_T;
    reg  [DATA_WIDTH-1:0] register [0:REG_NUM-1]; // 32 ta register 32bits
    
    // Address Read
    assign S_ARREADY = (state == RADDR_CHANNEL) ? 1 : 0;
    
    // Read
    assign S_RVALID = (state == RDATA_CHANNEL) ? 1 : 0;
    assign S_RDATA  = (state == RDATA_CHANNEL) ? register[read_addr] : 0;
    assign S_RRESP  = (state == RDATA_CHANNEL) ? 2'b00 : 0;

    // Address Write
    assign S_AWREADY = (state == WRITE_CHANNEL) ? 1 : 0;

    // Write
    assign S_WREADY = (state == WRITE_CHANNEL) ? 1 : 0;

    // Response
    assign S_BVALID = (state == WRESP_CHANNEL) ? 1 : 0;
    assign S_BRESP  = (state == WRESP_CHANNEL )? 0:0;

    assign S_ARADDR_T = S_ARADDR[ADDRESS-1:2]; // Read address 
    assign S_AWADDR_T = S_AWADDR[ADDRESS-1:2]; // Write address 
    
    always @(posedge ACLK) begin
        // Reset the register array
        if (~ARESETN) begin
            state <= IDLE;
        end
        else begin
            state <= next_state;
            if (state == WRITE_CHANNEL) begin
                register[S_AWADDR_T] <= S_WDATA;
            end
            else if (state == RADDR_CHANNEL) begin
                read_addr <= S_ARADDR_T;
            end
            else if (state == IDLE) begin
                start <= 0;
                rst <= 1;
            end
            else if (state == MY_STATE) begin
                start <= 1;
                rst <= 0;
                in_features = {register[23], register[22], register[21], register[20], register[19], register[18], register[17], register[16], register[15], register[14], register[13], register[12], register[11], register[10], register[9], register[8], register[7], register[6], register[5], register[4], register[3], register[2], register[1], register[0]};
                // in_features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000011111100000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000000000000000000101111111000000000000000000010100000111000000000000000001110000000110000000000000000110000000001000000000000000011000000000100000000000000000100000000010000000000000000010000000001000000000000000000110000001000000000000000000001111111000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                register[24] <= {28'h0000000, prediction};
            end
        end
    end

    // State machine
    always @(*) begin
        next_state = state;
        case (state)
            IDLE: begin
                if (S_AWVALID) begin
                    next_state = WRITE_CHANNEL;
                end 
                else if (S_ARVALID) begin
                    next_state = RADDR_CHANNEL;
                end 
                else begin
                    next_state = IDLE;
                end
            end

            RADDR_CHANNEL: begin
                if (S_ARVALID && S_ARREADY && S_ARADDR_T == 24)
                    next_state = MY_STATE;
                else if (S_ARVALID && S_ARREADY)
                    next_state = RDATA_CHANNEL;
            end

            MY_STATE: begin
                if (done)
                    next_state = RDATA_CHANNEL;
            end

            RDATA_CHANNEL: begin
                if (S_RVALID && S_RREADY)
                    next_state = IDLE;
            end

            WRITE_CHANNEL: begin
                if (S_AWVALID && S_AWREADY && S_WREADY && S_WVALID)
                    next_state = WRESP_CHANNEL;
            end

            WRESP_CHANNEL: begin
                if (S_BVALID && S_BREADY) 
                    next_state = IDLE;
            end

            default: begin
                next_state = IDLE;
            end 
        endcase
    end
endmodule

module NeuralNetwork (
    input clk,
    input rst,
    input start,
    input [783:0] in_features, // 784 input features
    output reg [3:0] prediction, // 10 output classes (ArgMax index)
    output reg done
);

    // register to hold the input features
    reg [783:0] features;

    // state machine
    localparam IDLE = 0, COMPUTE = 1;
    reg state;
    reg [2:0] count_clocks; 

    // Define the parameters for layer sizes
    parameter INPUT_SIZE = 784;
    parameter HIDDEN1_SIZE = 64;
    parameter HIDDEN2_SIZE = 32;
    parameter OUTPUT_SIZE = 10;

    // Define memory for weights and biases (assumed preloaded)
    wire signed [15:0] weights1;
    wire signed [15:0] biases1 [0:63];
    
    wire signed [15:0] weights2 [0:2047];
    wire signed [15:0] biases2 [0:31];
    
    wire signed [15:0] weights3 [0:319];
    wire signed [15:0] biases3 [0:9];

    // Define address registers for weights and biases
    reg [15:0] weights1_addr;
    // reg [15:0] weights2_addr;
    // reg [15:0] weights3_addr;

    // Instantiate the BRAM for weights1
    mem_weights1 mem_weights1(clk, weights1_addr, weights1);

    // Layer Outputs
    reg signed [15:0] hidden1 [0:HIDDEN1_SIZE-1];
    reg signed [15:0] hidden2 [0:HIDDEN2_SIZE-1];
    reg signed [15:0] output_layer [0:OUTPUT_SIZE-1];
    
    // ReLU activation function
    function signed [15:0] relu;
        input signed [15:0] x;
        begin
            relu = (x > 0) ? x : 0;
        end
    endfunction

    // Define the loop variables
    integer i, j, k;
    reg [5:0] i_neuron;

    // ============================================
    // combinational Computation of the neurons
    // ============================================

    // layer 1
    reg signed [15:0] new_hidden1 [0:HIDDEN1_SIZE-1];
    reg signed [15:0] neuron_out1 [0:HIDDEN1_SIZE-1];

    always @(*) begin
        for (i = 0; i < HIDDEN1_SIZE; i = i + 1) begin
            new_hidden1[i] = relu(neuron_out1[i] + biases1[i]); 
        end
    end

    always @(posedge clk) begin
        neuron_out1[i_neuron] = neuron_out1[i_neuron] + (features[k] == 1 ? weights1 : 0); 
    end

    // layer 2
    reg signed [15:0] new_hidden2 [0:HIDDEN2_SIZE-1];
    reg signed [31:0] multiplier_out2 [0:HIDDEN2_SIZE-1][0:HIDDEN1_SIZE-1];
    reg signed [15:0] shift_out2 [0:HIDDEN2_SIZE-1][0:HIDDEN1_SIZE-1];
    always @(*) begin
        for (i = 0; i < HIDDEN2_SIZE; i = i + 1) begin
            new_hidden2[i] = biases2[i];
            for (j = 0; j < HIDDEN1_SIZE; j = j + 1) begin
                multiplier_out2[i][j] = hidden1[j] * weights2[i*HIDDEN1_SIZE+j];
                shift_out2[i][j] = multiplier_out2[i][j] >> 8;
                new_hidden2[i] = new_hidden2[i] + shift_out2[i][j];
            end
            new_hidden2[i] = relu(new_hidden2[i]);
        end
    end

    // Output Layer computation
    reg signed [15:0] new_output_layer [0:OUTPUT_SIZE-1];
    reg signed [31:0] multiplier_out3 [0:OUTPUT_SIZE-1][0:HIDDEN2_SIZE-1];
    reg signed [15:0] shift_out3 [0:OUTPUT_SIZE-1][0:HIDDEN2_SIZE-1];
    always @(*) begin
        for (i = 0; i < OUTPUT_SIZE; i = i + 1) begin
            new_output_layer[i] = biases3[i];
            for (j = 0; j < HIDDEN2_SIZE; j = j + 1) begin
                multiplier_out3[i][j] = hidden2[j] * weights3[i*HIDDEN2_SIZE+j];
                shift_out3[i][j] = multiplier_out3[i][j] >> 8;
                new_output_layer[i] = new_output_layer[i] + shift_out3[i][j];
            end
        end
    end

    // ArgMax operation
    reg [3:0] new_prediction;
    always @(*) begin
        new_prediction = 0;
        for (i = 1; i < OUTPUT_SIZE; i = i + 1) begin
            if (output_layer[i] > output_layer[new_prediction]) begin
                new_prediction = i;
            end
        end
    end
    

    // ============================================
    // Sequential update of the neurons
    // ============================================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            done <= 0;
            count_clocks <= 0;
            prediction <= 0;
            weights1_addr <= 0;
            k <= 0;
            i_neuron <= 0;
            for (i = 0; i < INPUT_SIZE; i = i + 1) begin
                features[i] <= 0;
            end
        end 
        else if (state == IDLE) begin
            if (start) begin
                // Load the input features
                for (i = 0; i < INPUT_SIZE; i = i + 1) begin
                    features[i] <= in_features[i];
                end
                state <= COMPUTE;
                done <= 0;
                count_clocks <= 0;
                weights1_addr <= 0;
                k <= 0;
                i_neuron <= 0;
            end
        end 
        else begin
            // Layer 1 computation
            for (i = 0; i < HIDDEN1_SIZE; i = i + 1) begin
                hidden1[i] <= new_hidden1[i];
            end

            // Layer 2 computation
            for (i = 0; i < HIDDEN2_SIZE; i = i + 1) begin
                hidden2[i] <= new_hidden2[i];
            end

            // Output Layer computation
            for (i = 0; i < OUTPUT_SIZE; i = i + 1) begin
                output_layer[i] <= new_output_layer[i];
            end

            // ArgMax operation
            prediction <= new_prediction;

            // Update state or increment the clock counter
            if (count_clocks >= 3) begin
                state <= IDLE;
                done <= 1;
            end
            else begin
                count_clocks <= count_clocks + 1;
            end

            // Update the weights1 address
            if (weights1_addr >= 50175) begin
                weights1_addr <= 0;
            end
            else begin
                weights1_addr <= weights1_addr + 1;
            end
            if (k >= INPUT_SIZE - 1) begin
                k <= 0;
                i_neuron <= i_neuron + 1;
            end
            else begin
                k <= k + 1;
            end
        end
    end
    
    assign biases1[0] = 16'b0000000001110011;
    assign biases1[1] = 16'b0000000000100101;
    assign biases1[2] = 16'b0000000001000000;
    assign biases1[3] = 16'b0000000001010010;
    assign biases1[4] = 16'b1111111111100000;
    assign biases1[5] = 16'b0000000001000110;
    assign biases1[6] = 16'b0000000000000000;
    assign biases1[7] = 16'b0000000001010000;
    assign biases1[8] = 16'b1111111101110101;
    assign biases1[9] = 16'b1111111110010110;
    assign biases1[10] = 16'b1111111111001111;
    assign biases1[11] = 16'b0000000000011100;
    assign biases1[12] = 16'b0000000001000100;
    assign biases1[13] = 16'b0000000000011010;
    assign biases1[14] = 16'b1111111111111001;
    assign biases1[15] = 16'b1111111110010111;
    assign biases1[16] = 16'b1111111110010011;
    assign biases1[17] = 16'b0000000100011101;
    assign biases1[18] = 16'b0000000000011001;
    assign biases1[19] = 16'b1111111111111010;
    assign biases1[20] = 16'b0000000001001100;
    assign biases1[21] = 16'b0000000100001110;
    assign biases1[22] = 16'b0000000001000101;
    assign biases1[23] = 16'b1111111110100000;
    assign biases1[24] = 16'b0000000001001101;
    assign biases1[25] = 16'b0000000000011000;
    assign biases1[26] = 16'b1111111111101101;
    assign biases1[27] = 16'b0000000001001010;
    assign biases1[28] = 16'b0000000010000110;
    assign biases1[29] = 16'b0000000010011001;
    assign biases1[30] = 16'b0000000000010111;
    assign biases1[31] = 16'b0000000000100101;
    assign biases1[32] = 16'b1111111111110100;
    assign biases1[33] = 16'b1111111111101000;
    assign biases1[34] = 16'b0000000010011111;
    assign biases1[35] = 16'b0000000000110111;
    assign biases1[36] = 16'b0000000000001001;
    assign biases1[37] = 16'b0000000000101001;
    assign biases1[38] = 16'b0000000000011000;
    assign biases1[39] = 16'b0000000010011101;
    assign biases1[40] = 16'b1111111001101000;
    assign biases1[41] = 16'b1111111101011000;
    assign biases1[42] = 16'b0000000010010111;
    assign biases1[43] = 16'b0000000000000001;
    assign biases1[44] = 16'b0000000000011001;
    assign biases1[45] = 16'b1111111110001111;
    assign biases1[46] = 16'b0000000001000110;
    assign biases1[47] = 16'b0000000000101110;
    assign biases1[48] = 16'b0000000000110100;
    assign biases1[49] = 16'b0000000100010011;
    assign biases1[50] = 16'b0000000010000101;
    assign biases1[51] = 16'b1111111111111000;
    assign biases1[52] = 16'b0000000010010001;
    assign biases1[53] = 16'b1111111111110110;
    assign biases1[54] = 16'b0000000000000000;
    assign biases1[55] = 16'b0000000000000010;
    assign biases1[56] = 16'b0000000001000000;
    assign biases1[57] = 16'b0000000001001100;
    assign biases1[58] = 16'b1111111110100001;
    assign biases1[59] = 16'b0000000010010101;
    assign biases1[60] = 16'b1111111111100010;
    assign biases1[61] = 16'b0000000010100000;
    assign biases1[62] = 16'b0000000000001000;
    assign biases1[63] = 16'b1111111111101010;
    assign weights2[0] = 16'b0000000000000001;
    assign weights2[1] = 16'b1111111101101100;
    assign weights2[2] = 16'b0000000000000100;
    assign weights2[3] = 16'b1111111111001101;
    assign weights2[4] = 16'b0000000000001001;
    assign weights2[5] = 16'b1111111111110101;
    assign weights2[6] = 16'b0000000000000000;
    assign weights2[7] = 16'b1111111111110101;
    assign weights2[8] = 16'b0000000000100011;
    assign weights2[9] = 16'b0000000000010001;
    assign weights2[10] = 16'b1111111110001011;
    assign weights2[11] = 16'b0000000000001000;
    assign weights2[12] = 16'b1111111111010001;
    assign weights2[13] = 16'b1111111100110001;
    assign weights2[14] = 16'b1111111110101110;
    assign weights2[15] = 16'b0000000000011101;
    assign weights2[16] = 16'b0000000000010111;
    assign weights2[17] = 16'b0000000000110010;
    assign weights2[18] = 16'b1111111111111001;
    assign weights2[19] = 16'b1111111111110011;
    assign weights2[20] = 16'b1111111110100001;
    assign weights2[21] = 16'b0000000000011000;
    assign weights2[22] = 16'b0000000000000011;
    assign weights2[23] = 16'b0000000000001010;
    assign weights2[24] = 16'b1111111110111010;
    assign weights2[25] = 16'b0000000000000101;
    assign weights2[26] = 16'b0000000000001111;
    assign weights2[27] = 16'b1111111111010001;
    assign weights2[28] = 16'b1111111111100111;
    assign weights2[29] = 16'b0000000000000100;
    assign weights2[30] = 16'b0000000000000111;
    assign weights2[31] = 16'b1111111110011001;
    assign weights2[32] = 16'b0000000000011001;
    assign weights2[33] = 16'b0000000001000110;
    assign weights2[34] = 16'b1111111110100111;
    assign weights2[35] = 16'b1111111111100010;
    assign weights2[36] = 16'b1111111111010101;
    assign weights2[37] = 16'b1111111110011101;
    assign weights2[38] = 16'b1111111111100100;
    assign weights2[39] = 16'b1111111110011010;
    assign weights2[40] = 16'b0000000000001000;
    assign weights2[41] = 16'b1111111101100100;
    assign weights2[42] = 16'b0000000000011101;
    assign weights2[43] = 16'b1111111111001101;
    assign weights2[44] = 16'b0000000000100011;
    assign weights2[45] = 16'b0000000000101101;
    assign weights2[46] = 16'b1111111111111010;
    assign weights2[47] = 16'b1111111111110100;
    assign weights2[48] = 16'b0000000000101011;
    assign weights2[49] = 16'b0000000000100001;
    assign weights2[50] = 16'b1111111111011100;
    assign weights2[51] = 16'b0000000000001010;
    assign weights2[52] = 16'b0000000000101111;
    assign weights2[53] = 16'b1111111100100011;
    assign weights2[54] = 16'b0000000000000000;
    assign weights2[55] = 16'b0000000000010101;
    assign weights2[56] = 16'b1111111100010100;
    assign weights2[57] = 16'b1111111111101100;
    assign weights2[58] = 16'b1111111101010011;
    assign weights2[59] = 16'b1111111111111000;
    assign weights2[60] = 16'b0000000000001000;
    assign weights2[61] = 16'b0000000000011010;
    assign weights2[62] = 16'b0000000000001111;
    assign weights2[63] = 16'b1111111110001111;
    assign weights2[64] = 16'b1111111111110101;
    assign weights2[65] = 16'b0000000001100001;
    assign weights2[66] = 16'b1111111111001110;
    assign weights2[67] = 16'b1111111101111111;
    assign weights2[68] = 16'b1111111110010110;
    assign weights2[69] = 16'b0000000000001110;
    assign weights2[70] = 16'b0000000000000000;
    assign weights2[71] = 16'b0000000001110100;
    assign weights2[72] = 16'b0000000000011010;
    assign weights2[73] = 16'b1111111110110001;
    assign weights2[74] = 16'b0000000000100100;
    assign weights2[75] = 16'b1111111111111110;
    assign weights2[76] = 16'b0000000001101100;
    assign weights2[77] = 16'b0000000001111000;
    assign weights2[78] = 16'b1111111111110100;
    assign weights2[79] = 16'b0000000000001000;
    assign weights2[80] = 16'b0000000000001000;
    assign weights2[81] = 16'b1111111110110110;
    assign weights2[82] = 16'b1111111111110001;
    assign weights2[83] = 16'b1111111111010111;
    assign weights2[84] = 16'b1111111110010000;
    assign weights2[85] = 16'b1111111111010110;
    assign weights2[86] = 16'b1111111111100101;
    assign weights2[87] = 16'b1111111110110111;
    assign weights2[88] = 16'b1111111110000001;
    assign weights2[89] = 16'b1111111111110001;
    assign weights2[90] = 16'b1111111110011011;
    assign weights2[91] = 16'b0000000000100100;
    assign weights2[92] = 16'b0000000010010011;
    assign weights2[93] = 16'b1111111111100001;
    assign weights2[94] = 16'b1111111111110001;
    assign weights2[95] = 16'b1111111111111101;
    assign weights2[96] = 16'b1111111111100101;
    assign weights2[97] = 16'b1111111101111111;
    assign weights2[98] = 16'b1111111110000111;
    assign weights2[99] = 16'b1111111110110101;
    assign weights2[100] = 16'b0000000001001110;
    assign weights2[101] = 16'b1111111111110010;
    assign weights2[102] = 16'b1111111111011011;
    assign weights2[103] = 16'b0000000000010010;
    assign weights2[104] = 16'b0000000000000000;
    assign weights2[105] = 16'b0000000000110001;
    assign weights2[106] = 16'b1111111111001100;
    assign weights2[107] = 16'b1111111101010110;
    assign weights2[108] = 16'b0000000000001000;
    assign weights2[109] = 16'b1111111111011101;
    assign weights2[110] = 16'b0000000001101101;
    assign weights2[111] = 16'b0000000001001000;
    assign weights2[112] = 16'b0000000000101100;
    assign weights2[113] = 16'b1111111110111011;
    assign weights2[114] = 16'b0000000001010011;
    assign weights2[115] = 16'b0000000000000011;
    assign weights2[116] = 16'b1111111111000011;
    assign weights2[117] = 16'b0000000000010110;
    assign weights2[118] = 16'b0000000000000000;
    assign weights2[119] = 16'b1111111110111100;
    assign weights2[120] = 16'b0000000001101100;
    assign weights2[121] = 16'b1111111110101000;
    assign weights2[122] = 16'b0000000000011111;
    assign weights2[123] = 16'b1111111111011111;
    assign weights2[124] = 16'b1111111111110010;
    assign weights2[125] = 16'b1111111111011100;
    assign weights2[126] = 16'b0000000000101111;
    assign weights2[127] = 16'b1111111110111110;
    assign weights2[128] = 16'b0000000001111111;
    assign weights2[129] = 16'b1111111110100010;
    assign weights2[130] = 16'b0000000000011100;
    assign weights2[131] = 16'b0000000000000110;
    assign weights2[132] = 16'b1111111101110100;
    assign weights2[133] = 16'b0000000000001100;
    assign weights2[134] = 16'b0000000000000000;
    assign weights2[135] = 16'b1111111111110001;
    assign weights2[136] = 16'b0000000001001000;
    assign weights2[137] = 16'b1111111110101000;
    assign weights2[138] = 16'b1111111111011001;
    assign weights2[139] = 16'b1111111111100011;
    assign weights2[140] = 16'b1111111111110100;
    assign weights2[141] = 16'b1111111110011011;
    assign weights2[142] = 16'b0000000000000101;
    assign weights2[143] = 16'b0000000000101010;
    assign weights2[144] = 16'b0000000000111101;
    assign weights2[145] = 16'b0000000001011100;
    assign weights2[146] = 16'b0000000000011010;
    assign weights2[147] = 16'b0000000010000000;
    assign weights2[148] = 16'b0000000000010000;
    assign weights2[149] = 16'b0000000000111001;
    assign weights2[150] = 16'b0000000001111111;
    assign weights2[151] = 16'b0000000001010001;
    assign weights2[152] = 16'b1111111111111011;
    assign weights2[153] = 16'b0000000000010110;
    assign weights2[154] = 16'b1111111101101000;
    assign weights2[155] = 16'b0000000000111110;
    assign weights2[156] = 16'b1111111110100100;
    assign weights2[157] = 16'b1111111111111011;
    assign weights2[158] = 16'b0000000001110101;
    assign weights2[159] = 16'b1111111111111101;
    assign weights2[160] = 16'b0000000000010111;
    assign weights2[161] = 16'b1111111110010000;
    assign weights2[162] = 16'b1111111111111110;
    assign weights2[163] = 16'b1111111111011100;
    assign weights2[164] = 16'b1111111111111010;
    assign weights2[165] = 16'b1111111111111101;
    assign weights2[166] = 16'b0000000000100000;
    assign weights2[167] = 16'b1111111111001010;
    assign weights2[168] = 16'b0000000000000000;
    assign weights2[169] = 16'b1111111111101001;
    assign weights2[170] = 16'b0000000000100111;
    assign weights2[171] = 16'b0000000000000011;
    assign weights2[172] = 16'b0000000000100001;
    assign weights2[173] = 16'b0000000000000010;
    assign weights2[174] = 16'b1111111110110000;
    assign weights2[175] = 16'b1111111111011011;
    assign weights2[176] = 16'b0000000001000110;
    assign weights2[177] = 16'b0000000000110001;
    assign weights2[178] = 16'b1111111111111011;
    assign weights2[179] = 16'b1111111111111100;
    assign weights2[180] = 16'b0000000001000101;
    assign weights2[181] = 16'b1111111111011101;
    assign weights2[182] = 16'b0000000000000000;
    assign weights2[183] = 16'b1111111111001000;
    assign weights2[184] = 16'b1111111111010001;
    assign weights2[185] = 16'b1111111111111010;
    assign weights2[186] = 16'b1111111111101111;
    assign weights2[187] = 16'b0000000000000000;
    assign weights2[188] = 16'b0000000000001001;
    assign weights2[189] = 16'b0000000000011001;
    assign weights2[190] = 16'b0000000000110001;
    assign weights2[191] = 16'b1111111101010000;
    assign weights2[192] = 16'b1111111111111111;
    assign weights2[193] = 16'b1111111101111101;
    assign weights2[194] = 16'b1111111111111011;
    assign weights2[195] = 16'b1111111111100101;
    assign weights2[196] = 16'b1111111111100100;
    assign weights2[197] = 16'b1111111111001011;
    assign weights2[198] = 16'b0000000000000000;
    assign weights2[199] = 16'b1111111100011010;
    assign weights2[200] = 16'b1111111111010111;
    assign weights2[201] = 16'b1111111111111111;
    assign weights2[202] = 16'b1111111110011101;
    assign weights2[203] = 16'b1111111101011010;
    assign weights2[204] = 16'b1111111111111111;
    assign weights2[205] = 16'b1111111110000011;
    assign weights2[206] = 16'b1111111101110010;
    assign weights2[207] = 16'b0000000000001000;
    assign weights2[208] = 16'b1111111111111100;
    assign weights2[209] = 16'b1111111110001111;
    assign weights2[210] = 16'b1111111110001000;
    assign weights2[211] = 16'b1111111101111010;
    assign weights2[212] = 16'b1111111111111111;
    assign weights2[213] = 16'b1111111110101100;
    assign weights2[214] = 16'b1111111110111001;
    assign weights2[215] = 16'b1111111110010111;
    assign weights2[216] = 16'b0000000000011110;
    assign weights2[217] = 16'b0000000000001001;
    assign weights2[218] = 16'b1111111111110011;
    assign weights2[219] = 16'b1111111101010011;
    assign weights2[220] = 16'b0000000000001111;
    assign weights2[221] = 16'b0000000000010100;
    assign weights2[222] = 16'b1111111111110000;
    assign weights2[223] = 16'b1111111110010100;
    assign weights2[224] = 16'b0000000000011000;
    assign weights2[225] = 16'b1111111111111110;
    assign weights2[226] = 16'b1111111111110100;
    assign weights2[227] = 16'b1111111111111001;
    assign weights2[228] = 16'b1111111100111110;
    assign weights2[229] = 16'b1111111101111010;
    assign weights2[230] = 16'b1111111111110110;
    assign weights2[231] = 16'b1111111101111110;
    assign weights2[232] = 16'b1111111111111010;
    assign weights2[233] = 16'b1111111101111000;
    assign weights2[234] = 16'b0000000000101111;
    assign weights2[235] = 16'b0000000000100100;
    assign weights2[236] = 16'b0000000000001010;
    assign weights2[237] = 16'b0000000000010111;
    assign weights2[238] = 16'b0000000000101011;
    assign weights2[239] = 16'b1111111101111110;
    assign weights2[240] = 16'b0000000000011010;
    assign weights2[241] = 16'b0000000000100001;
    assign weights2[242] = 16'b0000000000001011;
    assign weights2[243] = 16'b0000000000010100;
    assign weights2[244] = 16'b0000000000100011;
    assign weights2[245] = 16'b1111111101100111;
    assign weights2[246] = 16'b0000000000000000;
    assign weights2[247] = 16'b0000000000010100;
    assign weights2[248] = 16'b1111111110111101;
    assign weights2[249] = 16'b0000000000110100;
    assign weights2[250] = 16'b1111111101101010;
    assign weights2[251] = 16'b0000000000011111;
    assign weights2[252] = 16'b1111111111111110;
    assign weights2[253] = 16'b0000000000011110;
    assign weights2[254] = 16'b0000000000001010;
    assign weights2[255] = 16'b1111111110001111;
    assign weights2[256] = 16'b1111111111101001;
    assign weights2[257] = 16'b1111111110011101;
    assign weights2[258] = 16'b0000000000111010;
    assign weights2[259] = 16'b0000000000100111;
    assign weights2[260] = 16'b0000000000010110;
    assign weights2[261] = 16'b0000000000011111;
    assign weights2[262] = 16'b0000000000000000;
    assign weights2[263] = 16'b1111111110000100;
    assign weights2[264] = 16'b1111111110100101;
    assign weights2[265] = 16'b0000000000000000;
    assign weights2[266] = 16'b0000000000000011;
    assign weights2[267] = 16'b0000000000001111;
    assign weights2[268] = 16'b1111111101011011;
    assign weights2[269] = 16'b1111111111000000;
    assign weights2[270] = 16'b0000000001101110;
    assign weights2[271] = 16'b1111111100111101;
    assign weights2[272] = 16'b1111111111110011;
    assign weights2[273] = 16'b0000000000011110;
    assign weights2[274] = 16'b1111111111111111;
    assign weights2[275] = 16'b0000000000010111;
    assign weights2[276] = 16'b0000000000110110;
    assign weights2[277] = 16'b0000000001000010;
    assign weights2[278] = 16'b0000000000000101;
    assign weights2[279] = 16'b1111111110111101;
    assign weights2[280] = 16'b0000000000110000;
    assign weights2[281] = 16'b0000000000001001;
    assign weights2[282] = 16'b1111111111111010;
    assign weights2[283] = 16'b1111111111100101;
    assign weights2[284] = 16'b1111111111111001;
    assign weights2[285] = 16'b0000000000000100;
    assign weights2[286] = 16'b0000000000100011;
    assign weights2[287] = 16'b0000000001011011;
    assign weights2[288] = 16'b0000000000001000;
    assign weights2[289] = 16'b1111111111011000;
    assign weights2[290] = 16'b0000000000101010;
    assign weights2[291] = 16'b1111111110001100;
    assign weights2[292] = 16'b1111111110101010;
    assign weights2[293] = 16'b0000000001100101;
    assign weights2[294] = 16'b0000000000100001;
    assign weights2[295] = 16'b0000000000101100;
    assign weights2[296] = 16'b1111111111001001;
    assign weights2[297] = 16'b0000000000011000;
    assign weights2[298] = 16'b0000000000110001;
    assign weights2[299] = 16'b0000000000101011;
    assign weights2[300] = 16'b0000000000000111;
    assign weights2[301] = 16'b1111111111100110;
    assign weights2[302] = 16'b0000000000010000;
    assign weights2[303] = 16'b1111111111010011;
    assign weights2[304] = 16'b1111111100000001;
    assign weights2[305] = 16'b0000000001000011;
    assign weights2[306] = 16'b0000000000000010;
    assign weights2[307] = 16'b0000000000000001;
    assign weights2[308] = 16'b1111111111101101;
    assign weights2[309] = 16'b0000000000111101;
    assign weights2[310] = 16'b0000000000000000;
    assign weights2[311] = 16'b1111111110001001;
    assign weights2[312] = 16'b0000000000010001;
    assign weights2[313] = 16'b0000000000101011;
    assign weights2[314] = 16'b0000000000101001;
    assign weights2[315] = 16'b0000000000000111;
    assign weights2[316] = 16'b1111111111111011;
    assign weights2[317] = 16'b0000000000011111;
    assign weights2[318] = 16'b1111111011111000;
    assign weights2[319] = 16'b1111111111111011;
    assign weights2[320] = 16'b0000000000001111;
    assign weights2[321] = 16'b1111111110101001;
    assign weights2[322] = 16'b0000000001000010;
    assign weights2[323] = 16'b0000000000110100;
    assign weights2[324] = 16'b0000000000110101;
    assign weights2[325] = 16'b0000000000010000;
    assign weights2[326] = 16'b0000000000000000;
    assign weights2[327] = 16'b1111111100001010;
    assign weights2[328] = 16'b1111111111001010;
    assign weights2[329] = 16'b0000000000001110;
    assign weights2[330] = 16'b1111111110110001;
    assign weights2[331] = 16'b0000000000010010;
    assign weights2[332] = 16'b1111111110000001;
    assign weights2[333] = 16'b1111111110101101;
    assign weights2[334] = 16'b0000000001110000;
    assign weights2[335] = 16'b1111111101101011;
    assign weights2[336] = 16'b0000000000100001;
    assign weights2[337] = 16'b1111111111110001;
    assign weights2[338] = 16'b0000000000001001;
    assign weights2[339] = 16'b0000000000100010;
    assign weights2[340] = 16'b0000000000101110;
    assign weights2[341] = 16'b0000000000111011;
    assign weights2[342] = 16'b0000000000100000;
    assign weights2[343] = 16'b1111111110100100;
    assign weights2[344] = 16'b0000000000000001;
    assign weights2[345] = 16'b0000000000010101;
    assign weights2[346] = 16'b0000000000010100;
    assign weights2[347] = 16'b1111111111011100;
    assign weights2[348] = 16'b1111111100010110;
    assign weights2[349] = 16'b1111111111011111;
    assign weights2[350] = 16'b1111111111110101;
    assign weights2[351] = 16'b0000000001011110;
    assign weights2[352] = 16'b0000000000110110;
    assign weights2[353] = 16'b0000000000001100;
    assign weights2[354] = 16'b0000000000010010;
    assign weights2[355] = 16'b1111111111101011;
    assign weights2[356] = 16'b1111111100110001;
    assign weights2[357] = 16'b0000000001110101;
    assign weights2[358] = 16'b1111111111101000;
    assign weights2[359] = 16'b0000000000010110;
    assign weights2[360] = 16'b1111111111101110;
    assign weights2[361] = 16'b0000000000000101;
    assign weights2[362] = 16'b0000000001101000;
    assign weights2[363] = 16'b1111111111110000;
    assign weights2[364] = 16'b0000000000101100;
    assign weights2[365] = 16'b0000000000000000;
    assign weights2[366] = 16'b1111111101101101;
    assign weights2[367] = 16'b1111111111011110;
    assign weights2[368] = 16'b1111111111001110;
    assign weights2[369] = 16'b0000000001011011;
    assign weights2[370] = 16'b1111111110101110;
    assign weights2[371] = 16'b0000000000000101;
    assign weights2[372] = 16'b0000000000110010;
    assign weights2[373] = 16'b0000000000110100;
    assign weights2[374] = 16'b0000000000000000;
    assign weights2[375] = 16'b1111111111111100;
    assign weights2[376] = 16'b0000000000011010;
    assign weights2[377] = 16'b1111111111111111;
    assign weights2[378] = 16'b1111111111111101;
    assign weights2[379] = 16'b0000000000010100;
    assign weights2[380] = 16'b0000000000101101;
    assign weights2[381] = 16'b0000000001000110;
    assign weights2[382] = 16'b1111111111100100;
    assign weights2[383] = 16'b0000000000001101;
    assign weights2[384] = 16'b0000000000000110;
    assign weights2[385] = 16'b0000000001000101;
    assign weights2[386] = 16'b1111111111000010;
    assign weights2[387] = 16'b0000000000000100;
    assign weights2[388] = 16'b1111111111110001;
    assign weights2[389] = 16'b1111111111010001;
    assign weights2[390] = 16'b0000000000000000;
    assign weights2[391] = 16'b1111111100101010;
    assign weights2[392] = 16'b1111111101111110;
    assign weights2[393] = 16'b0000000000100101;
    assign weights2[394] = 16'b1111111110011010;
    assign weights2[395] = 16'b1111111100010100;
    assign weights2[396] = 16'b0000000000111010;
    assign weights2[397] = 16'b0000000000111101;
    assign weights2[398] = 16'b1111111111111111;
    assign weights2[399] = 16'b1111111110111000;
    assign weights2[400] = 16'b0000000000001111;
    assign weights2[401] = 16'b1111111100111010;
    assign weights2[402] = 16'b1111111101000111;
    assign weights2[403] = 16'b1111111101000011;
    assign weights2[404] = 16'b1111111111011001;
    assign weights2[405] = 16'b1111111101101010;
    assign weights2[406] = 16'b1111111110011010;
    assign weights2[407] = 16'b1111111101010000;
    assign weights2[408] = 16'b0000000000000101;
    assign weights2[409] = 16'b1111111111110011;
    assign weights2[410] = 16'b1111111111011010;
    assign weights2[411] = 16'b1111111111000001;
    assign weights2[412] = 16'b1111111101101110;
    assign weights2[413] = 16'b0000000000000111;
    assign weights2[414] = 16'b1111111110011111;
    assign weights2[415] = 16'b1111111111111100;
    assign weights2[416] = 16'b0000000000101010;
    assign weights2[417] = 16'b1111111111110001;
    assign weights2[418] = 16'b1111111111111001;
    assign weights2[419] = 16'b1111111111111100;
    assign weights2[420] = 16'b1111111110000001;
    assign weights2[421] = 16'b0000000000000001;
    assign weights2[422] = 16'b1111111111011000;
    assign weights2[423] = 16'b1111111110011100;
    assign weights2[424] = 16'b1111111111101100;
    assign weights2[425] = 16'b1111111111110011;
    assign weights2[426] = 16'b1111111111010111;
    assign weights2[427] = 16'b0000000000010010;
    assign weights2[428] = 16'b0000000000011100;
    assign weights2[429] = 16'b0000000000011001;
    assign weights2[430] = 16'b1111111111101000;
    assign weights2[431] = 16'b1111111110100111;
    assign weights2[432] = 16'b1111111111110011;
    assign weights2[433] = 16'b1111111110100110;
    assign weights2[434] = 16'b1111111111110101;
    assign weights2[435] = 16'b0000000000001111;
    assign weights2[436] = 16'b1111111110100001;
    assign weights2[437] = 16'b0000000000001100;
    assign weights2[438] = 16'b0000000000000000;
    assign weights2[439] = 16'b0000000001000000;
    assign weights2[440] = 16'b0000000000101010;
    assign weights2[441] = 16'b0000000000001100;
    assign weights2[442] = 16'b1111111101110101;
    assign weights2[443] = 16'b0000000000010110;
    assign weights2[444] = 16'b1111111111110011;
    assign weights2[445] = 16'b1111111111111010;
    assign weights2[446] = 16'b0000000000001100;
    assign weights2[447] = 16'b0000000000101000;
    assign weights2[448] = 16'b0000000000010101;
    assign weights2[449] = 16'b1111111101011000;
    assign weights2[450] = 16'b0000000000011000;
    assign weights2[451] = 16'b1111111111111111;
    assign weights2[452] = 16'b1111111100000011;
    assign weights2[453] = 16'b1111111111101010;
    assign weights2[454] = 16'b0000000000000000;
    assign weights2[455] = 16'b1111111111011111;
    assign weights2[456] = 16'b0000000001000001;
    assign weights2[457] = 16'b1111111100110111;
    assign weights2[458] = 16'b0000000000001011;
    assign weights2[459] = 16'b1111111111100010;
    assign weights2[460] = 16'b1111111101000110;
    assign weights2[461] = 16'b1111111101101110;
    assign weights2[462] = 16'b0000000000010010;
    assign weights2[463] = 16'b1111111111100001;
    assign weights2[464] = 16'b0000000000011101;
    assign weights2[465] = 16'b0000000000110000;
    assign weights2[466] = 16'b0000000000001101;
    assign weights2[467] = 16'b0000000000000111;
    assign weights2[468] = 16'b1111111111110001;
    assign weights2[469] = 16'b0000000000101110;
    assign weights2[470] = 16'b0000000000100101;
    assign weights2[471] = 16'b0000000001000000;
    assign weights2[472] = 16'b0000000000001011;
    assign weights2[473] = 16'b0000000000001111;
    assign weights2[474] = 16'b1111111100111101;
    assign weights2[475] = 16'b1111111111001101;
    assign weights2[476] = 16'b1111111110110101;
    assign weights2[477] = 16'b1111111111111111;
    assign weights2[478] = 16'b1111111111111111;
    assign weights2[479] = 16'b0000000000001001;
    assign weights2[480] = 16'b1111111111111010;
    assign weights2[481] = 16'b1111111110010110;
    assign weights2[482] = 16'b0000000000000000;
    assign weights2[483] = 16'b1111111110101110;
    assign weights2[484] = 16'b0000000000010001;
    assign weights2[485] = 16'b0000000000010110;
    assign weights2[486] = 16'b0000000000100001;
    assign weights2[487] = 16'b1111111111100100;
    assign weights2[488] = 16'b1111111111110011;
    assign weights2[489] = 16'b1111111111101110;
    assign weights2[490] = 16'b0000000000100110;
    assign weights2[491] = 16'b0000000000001100;
    assign weights2[492] = 16'b1111111111110001;
    assign weights2[493] = 16'b0000000000000110;
    assign weights2[494] = 16'b1111111111110010;
    assign weights2[495] = 16'b1111111110000111;
    assign weights2[496] = 16'b1111111111001101;
    assign weights2[497] = 16'b0000000000100000;
    assign weights2[498] = 16'b0000000000011110;
    assign weights2[499] = 16'b0000000000000100;
    assign weights2[500] = 16'b0000000000010000;
    assign weights2[501] = 16'b1111111111111001;
    assign weights2[502] = 16'b0000000000000000;
    assign weights2[503] = 16'b1111111100011111;
    assign weights2[504] = 16'b1111111110100111;
    assign weights2[505] = 16'b0000000000001011;
    assign weights2[506] = 16'b0000000000001110;
    assign weights2[507] = 16'b0000000000010010;
    assign weights2[508] = 16'b0000000000100001;
    assign weights2[509] = 16'b0000000000011010;
    assign weights2[510] = 16'b1111111111001110;
    assign weights2[511] = 16'b1111111110011000;
    assign weights2[512] = 16'b1111111111000101;
    assign weights2[513] = 16'b0000000000011101;
    assign weights2[514] = 16'b1111111111011000;
    assign weights2[515] = 16'b1111111111000011;
    assign weights2[516] = 16'b1111111111010101;
    assign weights2[517] = 16'b1111111111001111;
    assign weights2[518] = 16'b0000000000000000;
    assign weights2[519] = 16'b0000000010110011;
    assign weights2[520] = 16'b0000000000111001;
    assign weights2[521] = 16'b1111111111110010;
    assign weights2[522] = 16'b0000000001011111;
    assign weights2[523] = 16'b0000000000000010;
    assign weights2[524] = 16'b0000000000101111;
    assign weights2[525] = 16'b0000000000011110;
    assign weights2[526] = 16'b1111111110011111;
    assign weights2[527] = 16'b0000000000001100;
    assign weights2[528] = 16'b1111111111111111;
    assign weights2[529] = 16'b0000000000011111;
    assign weights2[530] = 16'b0000000000000011;
    assign weights2[531] = 16'b0000000000010000;
    assign weights2[532] = 16'b1111111101111111;
    assign weights2[533] = 16'b1111111111011011;
    assign weights2[534] = 16'b0000000000001000;
    assign weights2[535] = 16'b0000000000010111;
    assign weights2[536] = 16'b0000000000010010;
    assign weights2[537] = 16'b1111111111011000;
    assign weights2[538] = 16'b1111111111101000;
    assign weights2[539] = 16'b0000000000011011;
    assign weights2[540] = 16'b0000000010011100;
    assign weights2[541] = 16'b0000000000011100;
    assign weights2[542] = 16'b0000000000001000;
    assign weights2[543] = 16'b1111111111000001;
    assign weights2[544] = 16'b1111111110101111;
    assign weights2[545] = 16'b0000000000010100;
    assign weights2[546] = 16'b1111111110110010;
    assign weights2[547] = 16'b1111111111110100;
    assign weights2[548] = 16'b0000000001000100;
    assign weights2[549] = 16'b1111111101100110;
    assign weights2[550] = 16'b1111111111111010;
    assign weights2[551] = 16'b1111111110101100;
    assign weights2[552] = 16'b0000000000000000;
    assign weights2[553] = 16'b0000000000101111;
    assign weights2[554] = 16'b1111111110101011;
    assign weights2[555] = 16'b0000000000010100;
    assign weights2[556] = 16'b1111111111001000;
    assign weights2[557] = 16'b0000000000000101;
    assign weights2[558] = 16'b0000000010001111;
    assign weights2[559] = 16'b0000000000001011;
    assign weights2[560] = 16'b0000000000010010;
    assign weights2[561] = 16'b1111111111000000;
    assign weights2[562] = 16'b0000000010011100;
    assign weights2[563] = 16'b1111111111110010;
    assign weights2[564] = 16'b1111111110101110;
    assign weights2[565] = 16'b1111111110110111;
    assign weights2[566] = 16'b1111111111111111;
    assign weights2[567] = 16'b1111111111001011;
    assign weights2[568] = 16'b0000000000000010;
    assign weights2[569] = 16'b0000000000001011;
    assign weights2[570] = 16'b0000000000011110;
    assign weights2[571] = 16'b1111111111001000;
    assign weights2[572] = 16'b1111111111100100;
    assign weights2[573] = 16'b1111111111011011;
    assign weights2[574] = 16'b0000000000010101;
    assign weights2[575] = 16'b1111111101000011;
    assign weights2[576] = 16'b0000000000001100;
    assign weights2[577] = 16'b1111111110010101;
    assign weights2[578] = 16'b0000000001001001;
    assign weights2[579] = 16'b0000000000111010;
    assign weights2[580] = 16'b0000000000110111;
    assign weights2[581] = 16'b0000000000010110;
    assign weights2[582] = 16'b0000000000000000;
    assign weights2[583] = 16'b0000000000111000;
    assign weights2[584] = 16'b0000000000100111;
    assign weights2[585] = 16'b0000000000010111;
    assign weights2[586] = 16'b1111111111100011;
    assign weights2[587] = 16'b0000000001001001;
    assign weights2[588] = 16'b1111111110001001;
    assign weights2[589] = 16'b1111111110101111;
    assign weights2[590] = 16'b0000000000101010;
    assign weights2[591] = 16'b1111111111100111;
    assign weights2[592] = 16'b1111111111111011;
    assign weights2[593] = 16'b0000000010001011;
    assign weights2[594] = 16'b0000000000110111;
    assign weights2[595] = 16'b0000000000111110;
    assign weights2[596] = 16'b1111111101011110;
    assign weights2[597] = 16'b0000000001111100;
    assign weights2[598] = 16'b0000000001001110;
    assign weights2[599] = 16'b0000000000101111;
    assign weights2[600] = 16'b0000000000101001;
    assign weights2[601] = 16'b1111111111111101;
    assign weights2[602] = 16'b0000000001001001;
    assign weights2[603] = 16'b0000000000000010;
    assign weights2[604] = 16'b0000000000010111;
    assign weights2[605] = 16'b1111111111111001;
    assign weights2[606] = 16'b0000000000101011;
    assign weights2[607] = 16'b0000000000100100;
    assign weights2[608] = 16'b1111111111111110;
    assign weights2[609] = 16'b0000000010100010;
    assign weights2[610] = 16'b0000000000011000;
    assign weights2[611] = 16'b1111111111000001;
    assign weights2[612] = 16'b0000000000001100;
    assign weights2[613] = 16'b0000000000110000;
    assign weights2[614] = 16'b0000000000110100;
    assign weights2[615] = 16'b0000000000110011;
    assign weights2[616] = 16'b1111111111011001;
    assign weights2[617] = 16'b1111111111001110;
    assign weights2[618] = 16'b0000000000100100;
    assign weights2[619] = 16'b0000000000111110;
    assign weights2[620] = 16'b0000000000000010;
    assign weights2[621] = 16'b0000000000001101;
    assign weights2[622] = 16'b0000000000001010;
    assign weights2[623] = 16'b0000000000000001;
    assign weights2[624] = 16'b1111111111101001;
    assign weights2[625] = 16'b0000000000011001;
    assign weights2[626] = 16'b0000000000001011;
    assign weights2[627] = 16'b1111111111010001;
    assign weights2[628] = 16'b0000000001001001;
    assign weights2[629] = 16'b0000000000110010;
    assign weights2[630] = 16'b0000000000000000;
    assign weights2[631] = 16'b0000000000101111;
    assign weights2[632] = 16'b1111111110111001;
    assign weights2[633] = 16'b0000000000100001;
    assign weights2[634] = 16'b1111111111001111;
    assign weights2[635] = 16'b0000000000000111;
    assign weights2[636] = 16'b1111111111100010;
    assign weights2[637] = 16'b0000000000011001;
    assign weights2[638] = 16'b1111111111110111;
    assign weights2[639] = 16'b0000000001000111;
    assign weights2[640] = 16'b0000000000011011;
    assign weights2[641] = 16'b0000000001101000;
    assign weights2[642] = 16'b1111111111010110;
    assign weights2[643] = 16'b1111111110010100;
    assign weights2[644] = 16'b1111111111110011;
    assign weights2[645] = 16'b0000000000001001;
    assign weights2[646] = 16'b0000000000000000;
    assign weights2[647] = 16'b0000000000010011;
    assign weights2[648] = 16'b0000000000011011;
    assign weights2[649] = 16'b0000000000001000;
    assign weights2[650] = 16'b0000000000010100;
    assign weights2[651] = 16'b0000000001111100;
    assign weights2[652] = 16'b0000000001000001;
    assign weights2[653] = 16'b0000000001101101;
    assign weights2[654] = 16'b0000000000111000;
    assign weights2[655] = 16'b1111111111111101;
    assign weights2[656] = 16'b0000000000110101;
    assign weights2[657] = 16'b0000000000111110;
    assign weights2[658] = 16'b0000000001110101;
    assign weights2[659] = 16'b0000000001010111;
    assign weights2[660] = 16'b0000000000100000;
    assign weights2[661] = 16'b0000000000111100;
    assign weights2[662] = 16'b0000000001111011;
    assign weights2[663] = 16'b0000000000101101;
    assign weights2[664] = 16'b1111111101011010;
    assign weights2[665] = 16'b1111111111110000;
    assign weights2[666] = 16'b0000000000000100;
    assign weights2[667] = 16'b0000000010111001;
    assign weights2[668] = 16'b1111111111100111;
    assign weights2[669] = 16'b1111111110110110;
    assign weights2[670] = 16'b1111111111110001;
    assign weights2[671] = 16'b0000000000110110;
    assign weights2[672] = 16'b0000000000000100;
    assign weights2[673] = 16'b1111111111100000;
    assign weights2[674] = 16'b1111111110100000;
    assign weights2[675] = 16'b1111111110101001;
    assign weights2[676] = 16'b0000000000100101;
    assign weights2[677] = 16'b0000000000110001;
    assign weights2[678] = 16'b1111111111100000;
    assign weights2[679] = 16'b1111111111111101;
    assign weights2[680] = 16'b1111111111111001;
    assign weights2[681] = 16'b0000000000011011;
    assign weights2[682] = 16'b1111111111100110;
    assign weights2[683] = 16'b1111111101101111;
    assign weights2[684] = 16'b1111111111111011;
    assign weights2[685] = 16'b1111111111010101;
    assign weights2[686] = 16'b0000000000011100;
    assign weights2[687] = 16'b0000000001110000;
    assign weights2[688] = 16'b1111111111110000;
    assign weights2[689] = 16'b1111111111110010;
    assign weights2[690] = 16'b0000000000100110;
    assign weights2[691] = 16'b1111111111100101;
    assign weights2[692] = 16'b1111111111111101;
    assign weights2[693] = 16'b0000000000010110;
    assign weights2[694] = 16'b0000000000000000;
    assign weights2[695] = 16'b1111111111110110;
    assign weights2[696] = 16'b0000000000110100;
    assign weights2[697] = 16'b1111111110001101;
    assign weights2[698] = 16'b0000000000000010;
    assign weights2[699] = 16'b1111111111101001;
    assign weights2[700] = 16'b0000000001000001;
    assign weights2[701] = 16'b1111111111110000;
    assign weights2[702] = 16'b1111111111110001;
    assign weights2[703] = 16'b1111111111010101;
    assign weights2[704] = 16'b0000000000000100;
    assign weights2[705] = 16'b1111111101111111;
    assign weights2[706] = 16'b1111111111100000;
    assign weights2[707] = 16'b1111111111001001;
    assign weights2[708] = 16'b0000000000010101;
    assign weights2[709] = 16'b1111111111101111;
    assign weights2[710] = 16'b0000000000000000;
    assign weights2[711] = 16'b0000000000010010;
    assign weights2[712] = 16'b0000000000111111;
    assign weights2[713] = 16'b0000000000000100;
    assign weights2[714] = 16'b1111111111001101;
    assign weights2[715] = 16'b1111111111111011;
    assign weights2[716] = 16'b1111111111000011;
    assign weights2[717] = 16'b1111111101011101;
    assign weights2[718] = 16'b1111111110010001;
    assign weights2[719] = 16'b1111111111101010;
    assign weights2[720] = 16'b0000000000100101;
    assign weights2[721] = 16'b1111111111010110;
    assign weights2[722] = 16'b0000000000001000;
    assign weights2[723] = 16'b1111111111011111;
    assign weights2[724] = 16'b1111111100100011;
    assign weights2[725] = 16'b0000000000001011;
    assign weights2[726] = 16'b0000000000011110;
    assign weights2[727] = 16'b0000000000101110;
    assign weights2[728] = 16'b1111111111100000;
    assign weights2[729] = 16'b1111111111001110;
    assign weights2[730] = 16'b0000000000001010;
    assign weights2[731] = 16'b1111111110000111;
    assign weights2[732] = 16'b1111111111000001;
    assign weights2[733] = 16'b1111111110110000;
    assign weights2[734] = 16'b1111111110101011;
    assign weights2[735] = 16'b1111111110010001;
    assign weights2[736] = 16'b1111111111010111;
    assign weights2[737] = 16'b0000000000110100;
    assign weights2[738] = 16'b1111111111000111;
    assign weights2[739] = 16'b0000000000001010;
    assign weights2[740] = 16'b0000000000101100;
    assign weights2[741] = 16'b1111111111000101;
    assign weights2[742] = 16'b1111111111101000;
    assign weights2[743] = 16'b1111111111010111;
    assign weights2[744] = 16'b0000000000001001;
    assign weights2[745] = 16'b1111111111110110;
    assign weights2[746] = 16'b1111111101101100;
    assign weights2[747] = 16'b1111111111100010;
    assign weights2[748] = 16'b1111111111110010;
    assign weights2[749] = 16'b0000000000001100;
    assign weights2[750] = 16'b1111111111111000;
    assign weights2[751] = 16'b1111111111010100;
    assign weights2[752] = 16'b1111111111111010;
    assign weights2[753] = 16'b1111111111000011;
    assign weights2[754] = 16'b1111111111100101;
    assign weights2[755] = 16'b0000000000000000;
    assign weights2[756] = 16'b1111111111110101;
    assign weights2[757] = 16'b1111111111100001;
    assign weights2[758] = 16'b0000000000000000;
    assign weights2[759] = 16'b1111111111001000;
    assign weights2[760] = 16'b1111111110111111;
    assign weights2[761] = 16'b1111111111010111;
    assign weights2[762] = 16'b1111111111111010;
    assign weights2[763] = 16'b1111111111000010;
    assign weights2[764] = 16'b1111111111011101;
    assign weights2[765] = 16'b1111111110111110;
    assign weights2[766] = 16'b0000000000001111;
    assign weights2[767] = 16'b0000000000100011;
    assign weights2[768] = 16'b1111111101111001;
    assign weights2[769] = 16'b0000000000000101;
    assign weights2[770] = 16'b0000000001010011;
    assign weights2[771] = 16'b0000000000111001;
    assign weights2[772] = 16'b1111111111111111;
    assign weights2[773] = 16'b1111111101100000;
    assign weights2[774] = 16'b0000000000000000;
    assign weights2[775] = 16'b0000000000100001;
    assign weights2[776] = 16'b0000000000011000;
    assign weights2[777] = 16'b1111111111100100;
    assign weights2[778] = 16'b1111111111100001;
    assign weights2[779] = 16'b0000000000100001;
    assign weights2[780] = 16'b1111111111101111;
    assign weights2[781] = 16'b0000000000001100;
    assign weights2[782] = 16'b0000000000011011;
    assign weights2[783] = 16'b0000000000000100;
    assign weights2[784] = 16'b1111111111100100;
    assign weights2[785] = 16'b0000000000100111;
    assign weights2[786] = 16'b0000000000001000;
    assign weights2[787] = 16'b0000000000001001;
    assign weights2[788] = 16'b0000000000011111;
    assign weights2[789] = 16'b0000000001101011;
    assign weights2[790] = 16'b1111111111011010;
    assign weights2[791] = 16'b0000000000001010;
    assign weights2[792] = 16'b0000000010111111;
    assign weights2[793] = 16'b0000000000110101;
    assign weights2[794] = 16'b0000000000011110;
    assign weights2[795] = 16'b0000000000101011;
    assign weights2[796] = 16'b0000000000101010;
    assign weights2[797] = 16'b0000000010001110;
    assign weights2[798] = 16'b0000000000000000;
    assign weights2[799] = 16'b0000000000011011;
    assign weights2[800] = 16'b1111111111010100;
    assign weights2[801] = 16'b0000000000000001;
    assign weights2[802] = 16'b0000000001000000;
    assign weights2[803] = 16'b0000000001100101;
    assign weights2[804] = 16'b1111111111110110;
    assign weights2[805] = 16'b0000000000010111;
    assign weights2[806] = 16'b0000000000011011;
    assign weights2[807] = 16'b0000000000001110;
    assign weights2[808] = 16'b1111111111100010;
    assign weights2[809] = 16'b0000000000001001;
    assign weights2[810] = 16'b0000000001001100;
    assign weights2[811] = 16'b0000000010011011;
    assign weights2[812] = 16'b1111111110101011;
    assign weights2[813] = 16'b0000000001001111;
    assign weights2[814] = 16'b0000000000101111;
    assign weights2[815] = 16'b0000000000100101;
    assign weights2[816] = 16'b0000000000100100;
    assign weights2[817] = 16'b0000000001110111;
    assign weights2[818] = 16'b0000000001101101;
    assign weights2[819] = 16'b0000000000011001;
    assign weights2[820] = 16'b0000000000111011;
    assign weights2[821] = 16'b0000000000011000;
    assign weights2[822] = 16'b0000000000000000;
    assign weights2[823] = 16'b0000000000001000;
    assign weights2[824] = 16'b0000000000001100;
    assign weights2[825] = 16'b0000000010010111;
    assign weights2[826] = 16'b1111111111100011;
    assign weights2[827] = 16'b0000000000100000;
    assign weights2[828] = 16'b0000000000100000;
    assign weights2[829] = 16'b0000000001011111;
    assign weights2[830] = 16'b0000000000111001;
    assign weights2[831] = 16'b1111111111101101;
    assign weights2[832] = 16'b1111111111011100;
    assign weights2[833] = 16'b1111111101111111;
    assign weights2[834] = 16'b0000000000000111;
    assign weights2[835] = 16'b0000000000101001;
    assign weights2[836] = 16'b1111111110100011;
    assign weights2[837] = 16'b1111111111111100;
    assign weights2[838] = 16'b0000000000000000;
    assign weights2[839] = 16'b1111111111110110;
    assign weights2[840] = 16'b0000000000010000;
    assign weights2[841] = 16'b1111111110010010;
    assign weights2[842] = 16'b0000000000010111;
    assign weights2[843] = 16'b1111111111001110;
    assign weights2[844] = 16'b1111111110001011;
    assign weights2[845] = 16'b1111111110100100;
    assign weights2[846] = 16'b0000000000000110;
    assign weights2[847] = 16'b1111111111111101;
    assign weights2[848] = 16'b1111111111111110;
    assign weights2[849] = 16'b1111111110110111;
    assign weights2[850] = 16'b1111111111001011;
    assign weights2[851] = 16'b1111111110101101;
    assign weights2[852] = 16'b1111111110100011;
    assign weights2[853] = 16'b1111111110111111;
    assign weights2[854] = 16'b1111111110110111;
    assign weights2[855] = 16'b0000000000001001;
    assign weights2[856] = 16'b1111111111111111;
    assign weights2[857] = 16'b1111111111111110;
    assign weights2[858] = 16'b1111111110011100;
    assign weights2[859] = 16'b1111111110000100;
    assign weights2[860] = 16'b1111111111000101;
    assign weights2[861] = 16'b1111111111110111;
    assign weights2[862] = 16'b1111111111010110;
    assign weights2[863] = 16'b1111111111111111;
    assign weights2[864] = 16'b1111111111101111;
    assign weights2[865] = 16'b1111111111001001;
    assign weights2[866] = 16'b0000000000000111;
    assign weights2[867] = 16'b1111111111001000;
    assign weights2[868] = 16'b0000000000011101;
    assign weights2[869] = 16'b0000000000001100;
    assign weights2[870] = 16'b0000000000010111;
    assign weights2[871] = 16'b1111111111110111;
    assign weights2[872] = 16'b0000000000001011;
    assign weights2[873] = 16'b1111111111111111;
    assign weights2[874] = 16'b1111111111010101;
    assign weights2[875] = 16'b0000000000100110;
    assign weights2[876] = 16'b1111111111110010;
    assign weights2[877] = 16'b0000000000101011;
    assign weights2[878] = 16'b1111111111001010;
    assign weights2[879] = 16'b1111111110111001;
    assign weights2[880] = 16'b1111111111010010;
    assign weights2[881] = 16'b1111111111110100;
    assign weights2[882] = 16'b1111111110101001;
    assign weights2[883] = 16'b0000000000001101;
    assign weights2[884] = 16'b1111111101111011;
    assign weights2[885] = 16'b1111111111101001;
    assign weights2[886] = 16'b0000000000000000;
    assign weights2[887] = 16'b1111111110110101;
    assign weights2[888] = 16'b1111111110011101;
    assign weights2[889] = 16'b0000000000101011;
    assign weights2[890] = 16'b0000000000100110;
    assign weights2[891] = 16'b1111111111000101;
    assign weights2[892] = 16'b1111111110110111;
    assign weights2[893] = 16'b1111111111110101;
    assign weights2[894] = 16'b1111111110101101;
    assign weights2[895] = 16'b1111111111111010;
    assign weights2[896] = 16'b0000000000000111;
    assign weights2[897] = 16'b1111111111101000;
    assign weights2[898] = 16'b1111111110100011;
    assign weights2[899] = 16'b1111111101111000;
    assign weights2[900] = 16'b1111111111010010;
    assign weights2[901] = 16'b1111111110100010;
    assign weights2[902] = 16'b0000000000000000;
    assign weights2[903] = 16'b1111111111111100;
    assign weights2[904] = 16'b1111111110100110;
    assign weights2[905] = 16'b1111111111101100;
    assign weights2[906] = 16'b1111111111000100;
    assign weights2[907] = 16'b1111111110101010;
    assign weights2[908] = 16'b1111111111101010;
    assign weights2[909] = 16'b1111111111100100;
    assign weights2[910] = 16'b0000000000000110;
    assign weights2[911] = 16'b0000000000000010;
    assign weights2[912] = 16'b0000000001001101;
    assign weights2[913] = 16'b1111111110101100;
    assign weights2[914] = 16'b1111111111000011;
    assign weights2[915] = 16'b1111111110110001;
    assign weights2[916] = 16'b0000000001100011;
    assign weights2[917] = 16'b1111111111101100;
    assign weights2[918] = 16'b1111111111101110;
    assign weights2[919] = 16'b1111111111100110;
    assign weights2[920] = 16'b1111111101011011;
    assign weights2[921] = 16'b0000000000100011;
    assign weights2[922] = 16'b1111111110111111;
    assign weights2[923] = 16'b1111111111001110;
    assign weights2[924] = 16'b0000000001001100;
    assign weights2[925] = 16'b1111111110110010;
    assign weights2[926] = 16'b1111111110011101;
    assign weights2[927] = 16'b0000000000000111;
    assign weights2[928] = 16'b0000000000010100;
    assign weights2[929] = 16'b1111111110110011;
    assign weights2[930] = 16'b1111111110000111;
    assign weights2[931] = 16'b1111111110001100;
    assign weights2[932] = 16'b1111111111011001;
    assign weights2[933] = 16'b0000000000000010;
    assign weights2[934] = 16'b1111111111001000;
    assign weights2[935] = 16'b1111111111110011;
    assign weights2[936] = 16'b1111111111110111;
    assign weights2[937] = 16'b0000000000001101;
    assign weights2[938] = 16'b0000000000011111;
    assign weights2[939] = 16'b1111111101101100;
    assign weights2[940] = 16'b0000000000011100;
    assign weights2[941] = 16'b1111111111010010;
    assign weights2[942] = 16'b0000000001010000;
    assign weights2[943] = 16'b1111111111011101;
    assign weights2[944] = 16'b1111111111100011;
    assign weights2[945] = 16'b0000000000101010;
    assign weights2[946] = 16'b0000000000001100;
    assign weights2[947] = 16'b0000000000010110;
    assign weights2[948] = 16'b0000000000011111;
    assign weights2[949] = 16'b0000000000001011;
    assign weights2[950] = 16'b0000000000000000;
    assign weights2[951] = 16'b1111111111101101;
    assign weights2[952] = 16'b0000000000000011;
    assign weights2[953] = 16'b1111111101111110;
    assign weights2[954] = 16'b0000000000000010;
    assign weights2[955] = 16'b0000000001001011;
    assign weights2[956] = 16'b0000000010000010;
    assign weights2[957] = 16'b0000000000010110;
    assign weights2[958] = 16'b1111111111010000;
    assign weights2[959] = 16'b1111111111010110;
    assign weights2[960] = 16'b1111111111000101;
    assign weights2[961] = 16'b1111111101000011;
    assign weights2[962] = 16'b0000000000011101;
    assign weights2[963] = 16'b0000000000011110;
    assign weights2[964] = 16'b0000000000001000;
    assign weights2[965] = 16'b0000000000100000;
    assign weights2[966] = 16'b0000000000000000;
    assign weights2[967] = 16'b1111111111111010;
    assign weights2[968] = 16'b0000000000000011;
    assign weights2[969] = 16'b0000000000000001;
    assign weights2[970] = 16'b0000000000000101;
    assign weights2[971] = 16'b1111111101001010;
    assign weights2[972] = 16'b1111111110111111;
    assign weights2[973] = 16'b1111111101111001;
    assign weights2[974] = 16'b0000000000001001;
    assign weights2[975] = 16'b0000000000010101;
    assign weights2[976] = 16'b1111111101100111;
    assign weights2[977] = 16'b0000000000111001;
    assign weights2[978] = 16'b1111111101000101;
    assign weights2[979] = 16'b1111111110100110;
    assign weights2[980] = 16'b1111111110110111;
    assign weights2[981] = 16'b0000000001100000;
    assign weights2[982] = 16'b1111111101000111;
    assign weights2[983] = 16'b1111111111111111;
    assign weights2[984] = 16'b0000000000111001;
    assign weights2[985] = 16'b1111111111011010;
    assign weights2[986] = 16'b1111111111111010;
    assign weights2[987] = 16'b1111111110001101;
    assign weights2[988] = 16'b0000000000110000;
    assign weights2[989] = 16'b0000000000101111;
    assign weights2[990] = 16'b0000000001011101;
    assign weights2[991] = 16'b0000000000000010;
    assign weights2[992] = 16'b1111111111111100;
    assign weights2[993] = 16'b0000000000001011;
    assign weights2[994] = 16'b0000000000010011;
    assign weights2[995] = 16'b1111111111111001;
    assign weights2[996] = 16'b0000000000000101;
    assign weights2[997] = 16'b0000000000001010;
    assign weights2[998] = 16'b0000000001001010;
    assign weights2[999] = 16'b1111111101111100;
    assign weights2[1000] = 16'b1111111111010111;
    assign weights2[1001] = 16'b1111111101111011;
    assign weights2[1002] = 16'b1111111111110010;
    assign weights2[1003] = 16'b0000000000110101;
    assign weights2[1004] = 16'b1111111111101101;
    assign weights2[1005] = 16'b0000000000101000;
    assign weights2[1006] = 16'b0000000000110011;
    assign weights2[1007] = 16'b1111111100111100;
    assign weights2[1008] = 16'b0000000000010010;
    assign weights2[1009] = 16'b0000000000101010;
    assign weights2[1010] = 16'b0000000000100110;
    assign weights2[1011] = 16'b1111111111010110;
    assign weights2[1012] = 16'b1111111110100000;
    assign weights2[1013] = 16'b1111111101110010;
    assign weights2[1014] = 16'b0000000000000000;
    assign weights2[1015] = 16'b1111111111110110;
    assign weights2[1016] = 16'b1111111110000011;
    assign weights2[1017] = 16'b0000000000110110;
    assign weights2[1018] = 16'b1111111111100010;
    assign weights2[1019] = 16'b1111111101110001;
    assign weights2[1020] = 16'b1111111101000010;
    assign weights2[1021] = 16'b0000000000010111;
    assign weights2[1022] = 16'b1111111111111000;
    assign weights2[1023] = 16'b0000000000100110;
    assign weights2[1024] = 16'b0000000000010010;
    assign weights2[1025] = 16'b0000000001101100;
    assign weights2[1026] = 16'b0000000001010010;
    assign weights2[1027] = 16'b0000000000101111;
    assign weights2[1028] = 16'b1111111101111010;
    assign weights2[1029] = 16'b0000000000110000;
    assign weights2[1030] = 16'b0000000000000000;
    assign weights2[1031] = 16'b0000000000110101;
    assign weights2[1032] = 16'b1111111111011110;
    assign weights2[1033] = 16'b1111111110100000;
    assign weights2[1034] = 16'b0000000000010011;
    assign weights2[1035] = 16'b0000000000100110;
    assign weights2[1036] = 16'b0000000001000110;
    assign weights2[1037] = 16'b0000000010000000;
    assign weights2[1038] = 16'b0000000001011011;
    assign weights2[1039] = 16'b1111111110111011;
    assign weights2[1040] = 16'b1111111111100110;
    assign weights2[1041] = 16'b0000000000100110;
    assign weights2[1042] = 16'b0000000000001111;
    assign weights2[1043] = 16'b0000000000011011;
    assign weights2[1044] = 16'b0000000001010001;
    assign weights2[1045] = 16'b0000000001001010;
    assign weights2[1046] = 16'b0000000000001100;
    assign weights2[1047] = 16'b1111111111010000;
    assign weights2[1048] = 16'b0000000000101011;
    assign weights2[1049] = 16'b0000000000010110;
    assign weights2[1050] = 16'b1111111110101011;
    assign weights2[1051] = 16'b0000000001000101;
    assign weights2[1052] = 16'b0000000001011111;
    assign weights2[1053] = 16'b0000000000111000;
    assign weights2[1054] = 16'b0000000001000111;
    assign weights2[1055] = 16'b0000000001000110;
    assign weights2[1056] = 16'b0000000000000101;
    assign weights2[1057] = 16'b1111111101111101;
    assign weights2[1058] = 16'b0000000000101000;
    assign weights2[1059] = 16'b1111111101100101;
    assign weights2[1060] = 16'b0000000000110111;
    assign weights2[1061] = 16'b0000000001001111;
    assign weights2[1062] = 16'b0000000000101001;
    assign weights2[1063] = 16'b0000000000101001;
    assign weights2[1064] = 16'b1111111110101111;
    assign weights2[1065] = 16'b0000000000001101;
    assign weights2[1066] = 16'b0000000000000100;
    assign weights2[1067] = 16'b0000000000011101;
    assign weights2[1068] = 16'b0000000000000111;
    assign weights2[1069] = 16'b1111111111111111;
    assign weights2[1070] = 16'b0000000000111010;
    assign weights2[1071] = 16'b0000000001011000;
    assign weights2[1072] = 16'b1111111111001101;
    assign weights2[1073] = 16'b0000000000101001;
    assign weights2[1074] = 16'b0000000001010101;
    assign weights2[1075] = 16'b1111111111100001;
    assign weights2[1076] = 16'b1111111111110000;
    assign weights2[1077] = 16'b0000000000101000;
    assign weights2[1078] = 16'b0000000000000000;
    assign weights2[1079] = 16'b1111111110000110;
    assign weights2[1080] = 16'b0000000001111001;
    assign weights2[1081] = 16'b0000000000011011;
    assign weights2[1082] = 16'b0000000000011001;
    assign weights2[1083] = 16'b0000000000001011;
    assign weights2[1084] = 16'b0000000000001101;
    assign weights2[1085] = 16'b0000000000101000;
    assign weights2[1086] = 16'b1111111110101110;
    assign weights2[1087] = 16'b1111111110110011;
    assign weights2[1088] = 16'b1111111110110110;
    assign weights2[1089] = 16'b0000000000000100;
    assign weights2[1090] = 16'b1111111111001011;
    assign weights2[1091] = 16'b1111111111110100;
    assign weights2[1092] = 16'b0000000001101111;
    assign weights2[1093] = 16'b1111111111110100;
    assign weights2[1094] = 16'b0000000000000000;
    assign weights2[1095] = 16'b1111111110110110;
    assign weights2[1096] = 16'b1111111101111100;
    assign weights2[1097] = 16'b0000000000101110;
    assign weights2[1098] = 16'b1111111111111010;
    assign weights2[1099] = 16'b1111111110101110;
    assign weights2[1100] = 16'b1111111111010010;
    assign weights2[1101] = 16'b0000000000011011;
    assign weights2[1102] = 16'b0000000000100000;
    assign weights2[1103] = 16'b1111111100101001;
    assign weights2[1104] = 16'b1111111111100110;
    assign weights2[1105] = 16'b1111111101110110;
    assign weights2[1106] = 16'b1111111101101110;
    assign weights2[1107] = 16'b1111111110010100;
    assign weights2[1108] = 16'b1111111111011001;
    assign weights2[1109] = 16'b1111111101111110;
    assign weights2[1110] = 16'b1111111110011110;
    assign weights2[1111] = 16'b1111111101001111;
    assign weights2[1112] = 16'b0000000000001010;
    assign weights2[1113] = 16'b1111111111011011;
    assign weights2[1114] = 16'b0000000000011110;
    assign weights2[1115] = 16'b1111111110111000;
    assign weights2[1116] = 16'b1111111111100111;
    assign weights2[1117] = 16'b1111111111110111;
    assign weights2[1118] = 16'b1111111110100111;
    assign weights2[1119] = 16'b0000000000100000;
    assign weights2[1120] = 16'b1111111111110011;
    assign weights2[1121] = 16'b0000000000011100;
    assign weights2[1122] = 16'b1111111111111001;
    assign weights2[1123] = 16'b1111111111000000;
    assign weights2[1124] = 16'b1111111111111100;
    assign weights2[1125] = 16'b0000000000110100;
    assign weights2[1126] = 16'b1111111111100001;
    assign weights2[1127] = 16'b0000000000111000;
    assign weights2[1128] = 16'b1111111111011001;
    assign weights2[1129] = 16'b0000000000011000;
    assign weights2[1130] = 16'b1111111110111101;
    assign weights2[1131] = 16'b0000000000000101;
    assign weights2[1132] = 16'b1111111111111100;
    assign weights2[1133] = 16'b1111111111111110;
    assign weights2[1134] = 16'b0000000000000000;
    assign weights2[1135] = 16'b1111111111101101;
    assign weights2[1136] = 16'b1111111101000000;
    assign weights2[1137] = 16'b1111111110111010;
    assign weights2[1138] = 16'b1111111111111010;
    assign weights2[1139] = 16'b0000000000000100;
    assign weights2[1140] = 16'b1111111111010000;
    assign weights2[1141] = 16'b0000000000000111;
    assign weights2[1142] = 16'b0000000000000000;
    assign weights2[1143] = 16'b1111111111111000;
    assign weights2[1144] = 16'b0000000000011000;
    assign weights2[1145] = 16'b1111111111111100;
    assign weights2[1146] = 16'b1111111111110101;
    assign weights2[1147] = 16'b1111111111000101;
    assign weights2[1148] = 16'b1111111111100010;
    assign weights2[1149] = 16'b1111111111010011;
    assign weights2[1150] = 16'b1111111110000000;
    assign weights2[1151] = 16'b0000000000100000;
    assign weights2[1152] = 16'b0000000001110100;
    assign weights2[1153] = 16'b0000000001101101;
    assign weights2[1154] = 16'b1111111111111010;
    assign weights2[1155] = 16'b0000000000000011;
    assign weights2[1156] = 16'b1111111111110110;
    assign weights2[1157] = 16'b0000000000100111;
    assign weights2[1158] = 16'b0000000000000000;
    assign weights2[1159] = 16'b1111111110110001;
    assign weights2[1160] = 16'b0000000000000101;
    assign weights2[1161] = 16'b1111111111111100;
    assign weights2[1162] = 16'b1111111111101100;
    assign weights2[1163] = 16'b0000000000111110;
    assign weights2[1164] = 16'b0000000001101011;
    assign weights2[1165] = 16'b0000000001101110;
    assign weights2[1166] = 16'b1111111111101011;
    assign weights2[1167] = 16'b0000000000001001;
    assign weights2[1168] = 16'b0000000001000101;
    assign weights2[1169] = 16'b0000000000010101;
    assign weights2[1170] = 16'b0000000000111110;
    assign weights2[1171] = 16'b0000000000110001;
    assign weights2[1172] = 16'b0000000000000011;
    assign weights2[1173] = 16'b0000000001000110;
    assign weights2[1174] = 16'b0000000001011101;
    assign weights2[1175] = 16'b1111111111100001;
    assign weights2[1176] = 16'b1111111111011110;
    assign weights2[1177] = 16'b0000000000110000;
    assign weights2[1178] = 16'b0000000000000011;
    assign weights2[1179] = 16'b0000000001011011;
    assign weights2[1180] = 16'b1111111111011010;
    assign weights2[1181] = 16'b1111111111110001;
    assign weights2[1182] = 16'b0000000001000011;
    assign weights2[1183] = 16'b1111111111100110;
    assign weights2[1184] = 16'b0000000001001010;
    assign weights2[1185] = 16'b1111111111111101;
    assign weights2[1186] = 16'b1111111111101110;
    assign weights2[1187] = 16'b0000000000001110;
    assign weights2[1188] = 16'b1111111101111011;
    assign weights2[1189] = 16'b1111111110110111;
    assign weights2[1190] = 16'b1111111111100110;
    assign weights2[1191] = 16'b1111111111010000;
    assign weights2[1192] = 16'b1111111111101001;
    assign weights2[1193] = 16'b0000000000000101;
    assign weights2[1194] = 16'b0000000000101001;
    assign weights2[1195] = 16'b1111111111001011;
    assign weights2[1196] = 16'b0000000001001001;
    assign weights2[1197] = 16'b1111111111111101;
    assign weights2[1198] = 16'b1111111111101101;
    assign weights2[1199] = 16'b0000000010000101;
    assign weights2[1200] = 16'b0000000000101010;
    assign weights2[1201] = 16'b0000000001010110;
    assign weights2[1202] = 16'b1111111111111010;
    assign weights2[1203] = 16'b1111111111110111;
    assign weights2[1204] = 16'b0000000010000011;
    assign weights2[1205] = 16'b0000000000010101;
    assign weights2[1206] = 16'b0000000000000000;
    assign weights2[1207] = 16'b0000000000001111;
    assign weights2[1208] = 16'b0000000001010000;
    assign weights2[1209] = 16'b1111111111011110;
    assign weights2[1210] = 16'b1111111110110111;
    assign weights2[1211] = 16'b0000000000101110;
    assign weights2[1212] = 16'b0000000001111101;
    assign weights2[1213] = 16'b0000000000110001;
    assign weights2[1214] = 16'b0000000000101101;
    assign weights2[1215] = 16'b1111111111110000;
    assign weights2[1216] = 16'b1111111111110011;
    assign weights2[1217] = 16'b0000000000010100;
    assign weights2[1218] = 16'b0000000000101110;
    assign weights2[1219] = 16'b0000000010001001;
    assign weights2[1220] = 16'b0000000000110101;
    assign weights2[1221] = 16'b0000000000010011;
    assign weights2[1222] = 16'b0000000000000000;
    assign weights2[1223] = 16'b1111111111011000;
    assign weights2[1224] = 16'b0000000001101001;
    assign weights2[1225] = 16'b0000000000001001;
    assign weights2[1226] = 16'b0000000000000010;
    assign weights2[1227] = 16'b0000000000010011;
    assign weights2[1228] = 16'b0000000000000011;
    assign weights2[1229] = 16'b0000000000011010;
    assign weights2[1230] = 16'b0000000000001001;
    assign weights2[1231] = 16'b0000000000000010;
    assign weights2[1232] = 16'b1111111111010100;
    assign weights2[1233] = 16'b0000000000010101;
    assign weights2[1234] = 16'b0000000000000010;
    assign weights2[1235] = 16'b1111111111111011;
    assign weights2[1236] = 16'b1111111110101011;
    assign weights2[1237] = 16'b0000000000101110;
    assign weights2[1238] = 16'b0000000000001111;
    assign weights2[1239] = 16'b0000000001001110;
    assign weights2[1240] = 16'b0000000010000101;
    assign weights2[1241] = 16'b1111111110111110;
    assign weights2[1242] = 16'b0000000000111010;
    assign weights2[1243] = 16'b0000000000101001;
    assign weights2[1244] = 16'b1111111101111101;
    assign weights2[1245] = 16'b0000000000110011;
    assign weights2[1246] = 16'b0000000000111010;
    assign weights2[1247] = 16'b0000000000010000;
    assign weights2[1248] = 16'b0000000000001000;
    assign weights2[1249] = 16'b0000000001001000;
    assign weights2[1250] = 16'b0000000001110110;
    assign weights2[1251] = 16'b0000000001011101;
    assign weights2[1252] = 16'b0000000000011010;
    assign weights2[1253] = 16'b0000000000000111;
    assign weights2[1254] = 16'b0000000000100101;
    assign weights2[1255] = 16'b0000000000000100;
    assign weights2[1256] = 16'b1111111111111101;
    assign weights2[1257] = 16'b0000000000000000;
    assign weights2[1258] = 16'b1111111111110000;
    assign weights2[1259] = 16'b0000000010000101;
    assign weights2[1260] = 16'b0000000000001000;
    assign weights2[1261] = 16'b0000000000001111;
    assign weights2[1262] = 16'b1111111101010011;
    assign weights2[1263] = 16'b0000000000110010;
    assign weights2[1264] = 16'b0000000000001100;
    assign weights2[1265] = 16'b1111111111111100;
    assign weights2[1266] = 16'b1111111110100101;
    assign weights2[1267] = 16'b1111111111010011;
    assign weights2[1268] = 16'b0000000000001010;
    assign weights2[1269] = 16'b1111111111110110;
    assign weights2[1270] = 16'b0000000000000000;
    assign weights2[1271] = 16'b0000000000100111;
    assign weights2[1272] = 16'b0000000000100110;
    assign weights2[1273] = 16'b0000000001101101;
    assign weights2[1274] = 16'b1111111111110011;
    assign weights2[1275] = 16'b1111111110101111;
    assign weights2[1276] = 16'b1111111110100110;
    assign weights2[1277] = 16'b1111111111100000;
    assign weights2[1278] = 16'b0000000000110000;
    assign weights2[1279] = 16'b0000000000011011;
    assign weights2[1280] = 16'b1111111111001000;
    assign weights2[1281] = 16'b1111111111101111;
    assign weights2[1282] = 16'b1111111111001011;
    assign weights2[1283] = 16'b1111111101100011;
    assign weights2[1284] = 16'b1111111111101011;
    assign weights2[1285] = 16'b1111111110010111;
    assign weights2[1286] = 16'b0000000000000000;
    assign weights2[1287] = 16'b0000000000110110;
    assign weights2[1288] = 16'b0000000000100110;
    assign weights2[1289] = 16'b1111111111110011;
    assign weights2[1290] = 16'b1111111110010001;
    assign weights2[1291] = 16'b1111111110011110;
    assign weights2[1292] = 16'b1111111111111011;
    assign weights2[1293] = 16'b1111111111110011;
    assign weights2[1294] = 16'b1111111110011001;
    assign weights2[1295] = 16'b0000000000000010;
    assign weights2[1296] = 16'b0000000000000000;
    assign weights2[1297] = 16'b1111111110101110;
    assign weights2[1298] = 16'b1111111110100001;
    assign weights2[1299] = 16'b1111111110111011;
    assign weights2[1300] = 16'b1111111111011110;
    assign weights2[1301] = 16'b1111111110100001;
    assign weights2[1302] = 16'b1111111110100000;
    assign weights2[1303] = 16'b0000000000001111;
    assign weights2[1304] = 16'b1111111111011011;
    assign weights2[1305] = 16'b0000000000100101;
    assign weights2[1306] = 16'b1111111111101100;
    assign weights2[1307] = 16'b1111111111101111;
    assign weights2[1308] = 16'b0000000001010101;
    assign weights2[1309] = 16'b0000000001001011;
    assign weights2[1310] = 16'b1111111110001110;
    assign weights2[1311] = 16'b1111111101110010;
    assign weights2[1312] = 16'b1111111111000000;
    assign weights2[1313] = 16'b1111111111111000;
    assign weights2[1314] = 16'b1111111100001011;
    assign weights2[1315] = 16'b0000000000011010;
    assign weights2[1316] = 16'b0000000001010000;
    assign weights2[1317] = 16'b1111111110111010;
    assign weights2[1318] = 16'b1111111110110010;
    assign weights2[1319] = 16'b1111111111010010;
    assign weights2[1320] = 16'b1111111111111000;
    assign weights2[1321] = 16'b1111111111111111;
    assign weights2[1322] = 16'b0000000000100110;
    assign weights2[1323] = 16'b0000000000010111;
    assign weights2[1324] = 16'b1111111110110100;
    assign weights2[1325] = 16'b0000000001100001;
    assign weights2[1326] = 16'b0000000001111001;
    assign weights2[1327] = 16'b1111111111100110;
    assign weights2[1328] = 16'b0000000000001100;
    assign weights2[1329] = 16'b0000000000111000;
    assign weights2[1330] = 16'b0000000001101111;
    assign weights2[1331] = 16'b0000000000110100;
    assign weights2[1332] = 16'b1111111111110001;
    assign weights2[1333] = 16'b0000000000000011;
    assign weights2[1334] = 16'b0000000000000000;
    assign weights2[1335] = 16'b1111111111110001;
    assign weights2[1336] = 16'b1111111111101011;
    assign weights2[1337] = 16'b0000000000000101;
    assign weights2[1338] = 16'b0000000000000001;
    assign weights2[1339] = 16'b0000000000001010;
    assign weights2[1340] = 16'b0000000000001100;
    assign weights2[1341] = 16'b0000000000111010;
    assign weights2[1342] = 16'b0000000000010001;
    assign weights2[1343] = 16'b0000000000000011;
    assign weights2[1344] = 16'b1111111100110100;
    assign weights2[1345] = 16'b1111111111111011;
    assign weights2[1346] = 16'b1111111110111111;
    assign weights2[1347] = 16'b1111111111101011;
    assign weights2[1348] = 16'b0000000000011100;
    assign weights2[1349] = 16'b1111111110010111;
    assign weights2[1350] = 16'b0000000000000000;
    assign weights2[1351] = 16'b0000000000101011;
    assign weights2[1352] = 16'b0000000000011110;
    assign weights2[1353] = 16'b0000000000001100;
    assign weights2[1354] = 16'b0000000000100111;
    assign weights2[1355] = 16'b1111111110000100;
    assign weights2[1356] = 16'b0000000000000110;
    assign weights2[1357] = 16'b0000000000011100;
    assign weights2[1358] = 16'b0000000000000001;
    assign weights2[1359] = 16'b0000000000000101;
    assign weights2[1360] = 16'b1111111111000100;
    assign weights2[1361] = 16'b1111111111111000;
    assign weights2[1362] = 16'b1111111100111111;
    assign weights2[1363] = 16'b1111111110110011;
    assign weights2[1364] = 16'b1111111110010111;
    assign weights2[1365] = 16'b1111111110110011;
    assign weights2[1366] = 16'b1111111100011111;
    assign weights2[1367] = 16'b0000000000010101;
    assign weights2[1368] = 16'b0000000000100010;
    assign weights2[1369] = 16'b1111111111001110;
    assign weights2[1370] = 16'b0000000000100110;
    assign weights2[1371] = 16'b1111111111101001;
    assign weights2[1372] = 16'b0000000010000111;
    assign weights2[1373] = 16'b0000000000101001;
    assign weights2[1374] = 16'b1111111101111000;
    assign weights2[1375] = 16'b0000000000001101;
    assign weights2[1376] = 16'b1111111110100100;
    assign weights2[1377] = 16'b0000000000100000;
    assign weights2[1378] = 16'b0000000000000001;
    assign weights2[1379] = 16'b1111111111100010;
    assign weights2[1380] = 16'b1111111110011101;
    assign weights2[1381] = 16'b1111111111111010;
    assign weights2[1382] = 16'b1111111111111010;
    assign weights2[1383] = 16'b0000000000101110;
    assign weights2[1384] = 16'b1111111111111010;
    assign weights2[1385] = 16'b0000000000110101;
    assign weights2[1386] = 16'b1111111111011111;
    assign weights2[1387] = 16'b0000000000101110;
    assign weights2[1388] = 16'b1111111110000110;
    assign weights2[1389] = 16'b0000000000101011;
    assign weights2[1390] = 16'b0000000010010001;
    assign weights2[1391] = 16'b1111111111110001;
    assign weights2[1392] = 16'b1111111111111001;
    assign weights2[1393] = 16'b1111111111010100;
    assign weights2[1394] = 16'b0000000001101001;
    assign weights2[1395] = 16'b0000000000001011;
    assign weights2[1396] = 16'b1111111110101100;
    assign weights2[1397] = 16'b0000000000001110;
    assign weights2[1398] = 16'b1111111111111111;
    assign weights2[1399] = 16'b1111111111111101;
    assign weights2[1400] = 16'b0000000000011000;
    assign weights2[1401] = 16'b0000000000101010;
    assign weights2[1402] = 16'b0000000000000101;
    assign weights2[1403] = 16'b1111111110101101;
    assign weights2[1404] = 16'b1111111111101101;
    assign weights2[1405] = 16'b1111111111110100;
    assign weights2[1406] = 16'b1111111111110000;
    assign weights2[1407] = 16'b0000000000010011;
    assign weights2[1408] = 16'b0000000000000100;
    assign weights2[1409] = 16'b1111111110101110;
    assign weights2[1410] = 16'b1111111110011011;
    assign weights2[1411] = 16'b1111111111100000;
    assign weights2[1412] = 16'b1111111110111001;
    assign weights2[1413] = 16'b1111111111100011;
    assign weights2[1414] = 16'b0000000000000000;
    assign weights2[1415] = 16'b0000000000101010;
    assign weights2[1416] = 16'b1111111111100110;
    assign weights2[1417] = 16'b1111111111101010;
    assign weights2[1418] = 16'b0000000000001110;
    assign weights2[1419] = 16'b0000000000000000;
    assign weights2[1420] = 16'b1111111111111011;
    assign weights2[1421] = 16'b0000000000101010;
    assign weights2[1422] = 16'b1111111101010111;
    assign weights2[1423] = 16'b0000000001011101;
    assign weights2[1424] = 16'b1111111111111000;
    assign weights2[1425] = 16'b1111111110000100;
    assign weights2[1426] = 16'b0000000000001010;
    assign weights2[1427] = 16'b1111111111110100;
    assign weights2[1428] = 16'b1111111111011011;
    assign weights2[1429] = 16'b1111111111011011;
    assign weights2[1430] = 16'b1111111111111111;
    assign weights2[1431] = 16'b1111111110101000;
    assign weights2[1432] = 16'b1111111111011011;
    assign weights2[1433] = 16'b1111111111111101;
    assign weights2[1434] = 16'b1111111111011000;
    assign weights2[1435] = 16'b1111111110110100;
    assign weights2[1436] = 16'b0000000001111111;
    assign weights2[1437] = 16'b0000000000001110;
    assign weights2[1438] = 16'b1111111111111000;
    assign weights2[1439] = 16'b1111111110000110;
    assign weights2[1440] = 16'b0000000000000111;
    assign weights2[1441] = 16'b0000000000000100;
    assign weights2[1442] = 16'b1111111111001101;
    assign weights2[1443] = 16'b0000000010110110;
    assign weights2[1444] = 16'b1111111111100001;
    assign weights2[1445] = 16'b1111111101010011;
    assign weights2[1446] = 16'b1111111111000001;
    assign weights2[1447] = 16'b1111111111110010;
    assign weights2[1448] = 16'b0000000000001111;
    assign weights2[1449] = 16'b1111111111101111;
    assign weights2[1450] = 16'b1111111111110011;
    assign weights2[1451] = 16'b1111111111101010;
    assign weights2[1452] = 16'b1111111111111111;
    assign weights2[1453] = 16'b1111111111111100;
    assign weights2[1454] = 16'b0000000000110001;
    assign weights2[1455] = 16'b0000000000011010;
    assign weights2[1456] = 16'b0000000010011110;
    assign weights2[1457] = 16'b1111111111000011;
    assign weights2[1458] = 16'b0000000000100000;
    assign weights2[1459] = 16'b0000000000011000;
    assign weights2[1460] = 16'b1111111111011000;
    assign weights2[1461] = 16'b1111111111000011;
    assign weights2[1462] = 16'b0000000000000000;
    assign weights2[1463] = 16'b1111111111100001;
    assign weights2[1464] = 16'b1111111111010100;
    assign weights2[1465] = 16'b1111111111100110;
    assign weights2[1466] = 16'b1111111111110101;
    assign weights2[1467] = 16'b0000000000000101;
    assign weights2[1468] = 16'b1111111111011111;
    assign weights2[1469] = 16'b1111111111111001;
    assign weights2[1470] = 16'b0000000001111100;
    assign weights2[1471] = 16'b1111111110101111;
    assign weights2[1472] = 16'b0000000000101011;
    assign weights2[1473] = 16'b1111111111111001;
    assign weights2[1474] = 16'b0000000000011010;
    assign weights2[1475] = 16'b1111111110001010;
    assign weights2[1476] = 16'b1111111110001111;
    assign weights2[1477] = 16'b0000000001001100;
    assign weights2[1478] = 16'b0000000000000000;
    assign weights2[1479] = 16'b1111111111101010;
    assign weights2[1480] = 16'b1111111111110101;
    assign weights2[1481] = 16'b1111111111101100;
    assign weights2[1482] = 16'b1111111111100100;
    assign weights2[1483] = 16'b1111111111111011;
    assign weights2[1484] = 16'b1111111111110110;
    assign weights2[1485] = 16'b0000000000000000;
    assign weights2[1486] = 16'b0000000000010100;
    assign weights2[1487] = 16'b0000000000000011;
    assign weights2[1488] = 16'b0000000000101110;
    assign weights2[1489] = 16'b0000000000001100;
    assign weights2[1490] = 16'b1111111111111001;
    assign weights2[1491] = 16'b0000000000100110;
    assign weights2[1492] = 16'b0000000000000111;
    assign weights2[1493] = 16'b1111111111110001;
    assign weights2[1494] = 16'b0000000000010011;
    assign weights2[1495] = 16'b1111111111100010;
    assign weights2[1496] = 16'b1111111110010101;
    assign weights2[1497] = 16'b1111111110111111;
    assign weights2[1498] = 16'b1111111101111011;
    assign weights2[1499] = 16'b1111111111110001;
    assign weights2[1500] = 16'b1111111111001111;
    assign weights2[1501] = 16'b1111111110000011;
    assign weights2[1502] = 16'b0000000001001001;
    assign weights2[1503] = 16'b0000000000000110;
    assign weights2[1504] = 16'b0000000001100111;
    assign weights2[1505] = 16'b1111111101000110;
    assign weights2[1506] = 16'b1111111111001100;
    assign weights2[1507] = 16'b1111111100110101;
    assign weights2[1508] = 16'b1111111111011110;
    assign weights2[1509] = 16'b0000000000001000;
    assign weights2[1510] = 16'b0000000000010100;
    assign weights2[1511] = 16'b1111111111110111;
    assign weights2[1512] = 16'b1111111111101111;
    assign weights2[1513] = 16'b0000000000000010;
    assign weights2[1514] = 16'b1111111111101011;
    assign weights2[1515] = 16'b1111111101101110;
    assign weights2[1516] = 16'b0000000001100110;
    assign weights2[1517] = 16'b1111111110101010;
    assign weights2[1518] = 16'b1111111111000101;
    assign weights2[1519] = 16'b1111111111110001;
    assign weights2[1520] = 16'b1111111111110101;
    assign weights2[1521] = 16'b1111111111010011;
    assign weights2[1522] = 16'b1111111110111001;
    assign weights2[1523] = 16'b1111111111101000;
    assign weights2[1524] = 16'b1111111111101010;
    assign weights2[1525] = 16'b1111111111111111;
    assign weights2[1526] = 16'b0000000000000000;
    assign weights2[1527] = 16'b1111111111010010;
    assign weights2[1528] = 16'b1111111111110111;
    assign weights2[1529] = 16'b1111111110010000;
    assign weights2[1530] = 16'b0000000000000000;
    assign weights2[1531] = 16'b1111111111101101;
    assign weights2[1532] = 16'b0000000000011100;
    assign weights2[1533] = 16'b1111111110100101;
    assign weights2[1534] = 16'b1111111110100110;
    assign weights2[1535] = 16'b1111111111100101;
    assign weights2[1536] = 16'b0000000000010100;
    assign weights2[1537] = 16'b1111111111100111;
    assign weights2[1538] = 16'b0000000001100001;
    assign weights2[1539] = 16'b0000000001111001;
    assign weights2[1540] = 16'b0000000000010001;
    assign weights2[1541] = 16'b0000000000000111;
    assign weights2[1542] = 16'b0000000000000000;
    assign weights2[1543] = 16'b1111111110100001;
    assign weights2[1544] = 16'b0000000000001101;
    assign weights2[1545] = 16'b0000000000001111;
    assign weights2[1546] = 16'b1111111100011011;
    assign weights2[1547] = 16'b1111111111111101;
    assign weights2[1548] = 16'b1111111111111000;
    assign weights2[1549] = 16'b1111111110111001;
    assign weights2[1550] = 16'b0000000000000101;
    assign weights2[1551] = 16'b0000000000010001;
    assign weights2[1552] = 16'b1111111111110111;
    assign weights2[1553] = 16'b0000000000011110;
    assign weights2[1554] = 16'b1111111111110000;
    assign weights2[1555] = 16'b0000000000000100;
    assign weights2[1556] = 16'b1111111111001000;
    assign weights2[1557] = 16'b0000000000110010;
    assign weights2[1558] = 16'b1111111111101110;
    assign weights2[1559] = 16'b0000000000001000;
    assign weights2[1560] = 16'b0000000001101011;
    assign weights2[1561] = 16'b0000000000010110;
    assign weights2[1562] = 16'b0000000000100110;
    assign weights2[1563] = 16'b1111111111111101;
    assign weights2[1564] = 16'b1111111110001101;
    assign weights2[1565] = 16'b0000000000111101;
    assign weights2[1566] = 16'b0000000000011111;
    assign weights2[1567] = 16'b1111111111111000;
    assign weights2[1568] = 16'b0000000000011111;
    assign weights2[1569] = 16'b0000000000010101;
    assign weights2[1570] = 16'b0000000001100110;
    assign weights2[1571] = 16'b0000000001100111;
    assign weights2[1572] = 16'b1111111110110101;
    assign weights2[1573] = 16'b1111111111111000;
    assign weights2[1574] = 16'b0000000000011110;
    assign weights2[1575] = 16'b1111111110011100;
    assign weights2[1576] = 16'b1111111111111011;
    assign weights2[1577] = 16'b1111111111001000;
    assign weights2[1578] = 16'b0000000000100111;
    assign weights2[1579] = 16'b0000000010000001;
    assign weights2[1580] = 16'b0000000000100001;
    assign weights2[1581] = 16'b0000000001010000;
    assign weights2[1582] = 16'b1111111110100000;
    assign weights2[1583] = 16'b1111111111010111;
    assign weights2[1584] = 16'b0000000000110111;
    assign weights2[1585] = 16'b0000000001001100;
    assign weights2[1586] = 16'b1111111111000101;
    assign weights2[1587] = 16'b1111111111111011;
    assign weights2[1588] = 16'b1111111111100110;
    assign weights2[1589] = 16'b0000000000000011;
    assign weights2[1590] = 16'b0000000000000000;
    assign weights2[1591] = 16'b0000000001001001;
    assign weights2[1592] = 16'b0000000000000000;
    assign weights2[1593] = 16'b0000000001111111;
    assign weights2[1594] = 16'b1111111110011110;
    assign weights2[1595] = 16'b0000000000010100;
    assign weights2[1596] = 16'b1111111111001001;
    assign weights2[1597] = 16'b0000000000101101;
    assign weights2[1598] = 16'b0000000001010011;
    assign weights2[1599] = 16'b0000000000011110;
    assign weights2[1600] = 16'b1111111110110000;
    assign weights2[1601] = 16'b1111111111001111;
    assign weights2[1602] = 16'b1111111111111111;
    assign weights2[1603] = 16'b0000000000100110;
    assign weights2[1604] = 16'b0000000000000100;
    assign weights2[1605] = 16'b1111111111101101;
    assign weights2[1606] = 16'b0000000000000000;
    assign weights2[1607] = 16'b1111111111101010;
    assign weights2[1608] = 16'b1111111111111110;
    assign weights2[1609] = 16'b0000000000010010;
    assign weights2[1610] = 16'b1111111111110110;
    assign weights2[1611] = 16'b1111111101111111;
    assign weights2[1612] = 16'b1111111111000011;
    assign weights2[1613] = 16'b1111111111101000;
    assign weights2[1614] = 16'b0000000000111100;
    assign weights2[1615] = 16'b1111111111110101;
    assign weights2[1616] = 16'b0000000000000110;
    assign weights2[1617] = 16'b1111111110110100;
    assign weights2[1618] = 16'b1111111110000010;
    assign weights2[1619] = 16'b1111111110100010;
    assign weights2[1620] = 16'b0000000000000100;
    assign weights2[1621] = 16'b1111111111010010;
    assign weights2[1622] = 16'b1111111101111100;
    assign weights2[1623] = 16'b0000000000011100;
    assign weights2[1624] = 16'b1111111111111111;
    assign weights2[1625] = 16'b1111111110111100;
    assign weights2[1626] = 16'b1111111111110110;
    assign weights2[1627] = 16'b1111111110110001;
    assign weights2[1628] = 16'b1111111110101111;
    assign weights2[1629] = 16'b1111111111110010;
    assign weights2[1630] = 16'b1111111110110101;
    assign weights2[1631] = 16'b0000000000101100;
    assign weights2[1632] = 16'b1111111111111000;
    assign weights2[1633] = 16'b1111111111011011;
    assign weights2[1634] = 16'b0000000000011110;
    assign weights2[1635] = 16'b1111111110010111;
    assign weights2[1636] = 16'b0000000000101000;
    assign weights2[1637] = 16'b0000000000111011;
    assign weights2[1638] = 16'b1111111111101111;
    assign weights2[1639] = 16'b1111111101011110;
    assign weights2[1640] = 16'b1111111111110011;
    assign weights2[1641] = 16'b0000000000111010;
    assign weights2[1642] = 16'b1111111110010111;
    assign weights2[1643] = 16'b1111111111101001;
    assign weights2[1644] = 16'b1111111111111001;
    assign weights2[1645] = 16'b0000000000001011;
    assign weights2[1646] = 16'b1111111110011000;
    assign weights2[1647] = 16'b1111111110101010;
    assign weights2[1648] = 16'b1111111111000110;
    assign weights2[1649] = 16'b1111111111010111;
    assign weights2[1650] = 16'b1111111110101001;
    assign weights2[1651] = 16'b1111111111110010;
    assign weights2[1652] = 16'b1111111110000011;
    assign weights2[1653] = 16'b0000000000100101;
    assign weights2[1654] = 16'b0000000000000000;
    assign weights2[1655] = 16'b1111111111101001;
    assign weights2[1656] = 16'b1111111111111100;
    assign weights2[1657] = 16'b1111111111110011;
    assign weights2[1658] = 16'b0000000000110001;
    assign weights2[1659] = 16'b1111111110100101;
    assign weights2[1660] = 16'b1111111111101001;
    assign weights2[1661] = 16'b1111111110110110;
    assign weights2[1662] = 16'b1111111110101011;
    assign weights2[1663] = 16'b1111111111100010;
    assign weights2[1664] = 16'b1111111111110010;
    assign weights2[1665] = 16'b0000000000111001;
    assign weights2[1666] = 16'b1111111111111111;
    assign weights2[1667] = 16'b0000000001101111;
    assign weights2[1668] = 16'b1111111111100000;
    assign weights2[1669] = 16'b0000000000010011;
    assign weights2[1670] = 16'b0000000000000000;
    assign weights2[1671] = 16'b1111111111111001;
    assign weights2[1672] = 16'b1111111111110111;
    assign weights2[1673] = 16'b1111111111101100;
    assign weights2[1674] = 16'b0000000000111111;
    assign weights2[1675] = 16'b1111111111010001;
    assign weights2[1676] = 16'b0000000000100101;
    assign weights2[1677] = 16'b0000000000111000;
    assign weights2[1678] = 16'b0000000000000111;
    assign weights2[1679] = 16'b0000000000000011;
    assign weights2[1680] = 16'b1111111111111100;
    assign weights2[1681] = 16'b1111111111101000;
    assign weights2[1682] = 16'b1111111111100100;
    assign weights2[1683] = 16'b1111111111011011;
    assign weights2[1684] = 16'b1111111110110101;
    assign weights2[1685] = 16'b1111111111011000;
    assign weights2[1686] = 16'b1111111111101101;
    assign weights2[1687] = 16'b1111111111101001;
    assign weights2[1688] = 16'b0000000001011101;
    assign weights2[1689] = 16'b1111111110000001;
    assign weights2[1690] = 16'b1111111111100011;
    assign weights2[1691] = 16'b0000000000000010;
    assign weights2[1692] = 16'b1111111111000100;
    assign weights2[1693] = 16'b1111111111110100;
    assign weights2[1694] = 16'b0000000000110010;
    assign weights2[1695] = 16'b0000000000010001;
    assign weights2[1696] = 16'b0000000000011110;
    assign weights2[1697] = 16'b1111111111110100;
    assign weights2[1698] = 16'b0000000001101110;
    assign weights2[1699] = 16'b1111111111001001;
    assign weights2[1700] = 16'b1111111111011000;
    assign weights2[1701] = 16'b0000000000000100;
    assign weights2[1702] = 16'b0000000000010111;
    assign weights2[1703] = 16'b0000000000010011;
    assign weights2[1704] = 16'b1111111111110110;
    assign weights2[1705] = 16'b0000000000110011;
    assign weights2[1706] = 16'b1111111110110001;
    assign weights2[1707] = 16'b0000000000110010;
    assign weights2[1708] = 16'b0000000000010111;
    assign weights2[1709] = 16'b1111111111010000;
    assign weights2[1710] = 16'b1111111101001011;
    assign weights2[1711] = 16'b0000000000010111;
    assign weights2[1712] = 16'b0000000000011011;
    assign weights2[1713] = 16'b1111111110101101;
    assign weights2[1714] = 16'b1111111100111110;
    assign weights2[1715] = 16'b1111111111101100;
    assign weights2[1716] = 16'b1111111111000000;
    assign weights2[1717] = 16'b0000000000000000;
    assign weights2[1718] = 16'b0000000000000000;
    assign weights2[1719] = 16'b1111111111101110;
    assign weights2[1720] = 16'b0000000001010100;
    assign weights2[1721] = 16'b0000000000110010;
    assign weights2[1722] = 16'b0000000001001011;
    assign weights2[1723] = 16'b1111111110011001;
    assign weights2[1724] = 16'b1111111111001011;
    assign weights2[1725] = 16'b1111111101000110;
    assign weights2[1726] = 16'b0000000000000101;
    assign weights2[1727] = 16'b1111111111000000;
    assign weights2[1728] = 16'b1111111111100110;
    assign weights2[1729] = 16'b0000000001010010;
    assign weights2[1730] = 16'b1111111111011000;
    assign weights2[1731] = 16'b0000000000010011;
    assign weights2[1732] = 16'b1111111110000001;
    assign weights2[1733] = 16'b1111111111100101;
    assign weights2[1734] = 16'b0000000000000000;
    assign weights2[1735] = 16'b0000000000100111;
    assign weights2[1736] = 16'b1111111111011110;
    assign weights2[1737] = 16'b1111111111111011;
    assign weights2[1738] = 16'b0000000000010011;
    assign weights2[1739] = 16'b0000000001010100;
    assign weights2[1740] = 16'b0000000000010101;
    assign weights2[1741] = 16'b0000000001111001;
    assign weights2[1742] = 16'b0000000000011110;
    assign weights2[1743] = 16'b1111111111100110;
    assign weights2[1744] = 16'b0000000000010001;
    assign weights2[1745] = 16'b1111111111110111;
    assign weights2[1746] = 16'b0000000000101100;
    assign weights2[1747] = 16'b0000000001011101;
    assign weights2[1748] = 16'b0000000001001101;
    assign weights2[1749] = 16'b1111111111101000;
    assign weights2[1750] = 16'b0000000000110010;
    assign weights2[1751] = 16'b1111111110011000;
    assign weights2[1752] = 16'b0000000000000111;
    assign weights2[1753] = 16'b0000000000001010;
    assign weights2[1754] = 16'b0000000000001101;
    assign weights2[1755] = 16'b0000000001011010;
    assign weights2[1756] = 16'b0000000001001111;
    assign weights2[1757] = 16'b0000000000000011;
    assign weights2[1758] = 16'b0000000000110100;
    assign weights2[1759] = 16'b0000000000100011;
    assign weights2[1760] = 16'b1111111111111100;
    assign weights2[1761] = 16'b0000000000000001;
    assign weights2[1762] = 16'b0000000000010011;
    assign weights2[1763] = 16'b1111111101010000;
    assign weights2[1764] = 16'b1111111111111111;
    assign weights2[1765] = 16'b0000000000100100;
    assign weights2[1766] = 16'b1111111111011101;
    assign weights2[1767] = 16'b0000000010000110;
    assign weights2[1768] = 16'b1111111111111110;
    assign weights2[1769] = 16'b0000000000110111;
    assign weights2[1770] = 16'b0000000000001000;
    assign weights2[1771] = 16'b1111111111111101;
    assign weights2[1772] = 16'b1111111111001010;
    assign weights2[1773] = 16'b1111111111101100;
    assign weights2[1774] = 16'b0000000000010111;
    assign weights2[1775] = 16'b0000000010011101;
    assign weights2[1776] = 16'b1111111111010111;
    assign weights2[1777] = 16'b1111111111110110;
    assign weights2[1778] = 16'b1111111111110111;
    assign weights2[1779] = 16'b0000000000001101;
    assign weights2[1780] = 16'b0000000000010101;
    assign weights2[1781] = 16'b0000000001100001;
    assign weights2[1782] = 16'b0000000000000000;
    assign weights2[1783] = 16'b1111111110111100;
    assign weights2[1784] = 16'b0000000010000010;
    assign weights2[1785] = 16'b0000000000000101;
    assign weights2[1786] = 16'b0000000000001010;
    assign weights2[1787] = 16'b0000000000010100;
    assign weights2[1788] = 16'b0000000000101010;
    assign weights2[1789] = 16'b1111111111111010;
    assign weights2[1790] = 16'b1111111110111111;
    assign weights2[1791] = 16'b1111111111000110;
    assign weights2[1792] = 16'b0000000000110101;
    assign weights2[1793] = 16'b1111111111101110;
    assign weights2[1794] = 16'b1111111111100111;
    assign weights2[1795] = 16'b1111111111111011;
    assign weights2[1796] = 16'b1111111111110010;
    assign weights2[1797] = 16'b0000000000100100;
    assign weights2[1798] = 16'b0000000000000000;
    assign weights2[1799] = 16'b0000000000001101;
    assign weights2[1800] = 16'b0000000000110101;
    assign weights2[1801] = 16'b1111111111110110;
    assign weights2[1802] = 16'b0000000000001000;
    assign weights2[1803] = 16'b0000000000111111;
    assign weights2[1804] = 16'b1111111111111011;
    assign weights2[1805] = 16'b1111111111110000;
    assign weights2[1806] = 16'b1111111111100100;
    assign weights2[1807] = 16'b0000000000000101;
    assign weights2[1808] = 16'b0000000000110000;
    assign weights2[1809] = 16'b0000000001000001;
    assign weights2[1810] = 16'b0000000001100111;
    assign weights2[1811] = 16'b0000000010010101;
    assign weights2[1812] = 16'b1111111110011100;
    assign weights2[1813] = 16'b0000000000110111;
    assign weights2[1814] = 16'b0000000010010010;
    assign weights2[1815] = 16'b0000000001001010;
    assign weights2[1816] = 16'b1111111111000111;
    assign weights2[1817] = 16'b1111111101010010;
    assign weights2[1818] = 16'b0000000000000001;
    assign weights2[1819] = 16'b0000000000010001;
    assign weights2[1820] = 16'b1111111111000101;
    assign weights2[1821] = 16'b1111111101001110;
    assign weights2[1822] = 16'b0000000001110101;
    assign weights2[1823] = 16'b1111111111100001;
    assign weights2[1824] = 16'b0000000000010000;
    assign weights2[1825] = 16'b0000000000011101;
    assign weights2[1826] = 16'b0000000000000101;
    assign weights2[1827] = 16'b0000000000000000;
    assign weights2[1828] = 16'b0000000000100111;
    assign weights2[1829] = 16'b1111111111011100;
    assign weights2[1830] = 16'b1111111111111101;
    assign weights2[1831] = 16'b1111111110011110;
    assign weights2[1832] = 16'b0000000000001011;
    assign weights2[1833] = 16'b0000000000001111;
    assign weights2[1834] = 16'b1111111111000011;
    assign weights2[1835] = 16'b1111111111010111;
    assign weights2[1836] = 16'b0000000000010000;
    assign weights2[1837] = 16'b1111111111100010;
    assign weights2[1838] = 16'b1111111110111001;
    assign weights2[1839] = 16'b0000000000000010;
    assign weights2[1840] = 16'b0000000000010000;
    assign weights2[1841] = 16'b1111111110111110;
    assign weights2[1842] = 16'b1111111101100000;
    assign weights2[1843] = 16'b1111111111001101;
    assign weights2[1844] = 16'b0000000000000101;
    assign weights2[1845] = 16'b1111111111100010;
    assign weights2[1846] = 16'b0000000000000000;
    assign weights2[1847] = 16'b1111111111101001;
    assign weights2[1848] = 16'b1111111111111100;
    assign weights2[1849] = 16'b1111111110101000;
    assign weights2[1850] = 16'b1111111111111100;
    assign weights2[1851] = 16'b1111111101000010;
    assign weights2[1852] = 16'b0000000000000111;
    assign weights2[1853] = 16'b1111111110101011;
    assign weights2[1854] = 16'b0000000000000100;
    assign weights2[1855] = 16'b1111111110101011;
    assign weights2[1856] = 16'b0000000001011111;
    assign weights2[1857] = 16'b0000000000011101;
    assign weights2[1858] = 16'b0000000001011000;
    assign weights2[1859] = 16'b0000000000011011;
    assign weights2[1860] = 16'b1111111111111111;
    assign weights2[1861] = 16'b0000000001101101;
    assign weights2[1862] = 16'b0000000000000000;
    assign weights2[1863] = 16'b1111111111110101;
    assign weights2[1864] = 16'b0000000000100011;
    assign weights2[1865] = 16'b1111111111111011;
    assign weights2[1866] = 16'b1111111111110010;
    assign weights2[1867] = 16'b0000000000111010;
    assign weights2[1868] = 16'b0000000000011010;
    assign weights2[1869] = 16'b0000000000000100;
    assign weights2[1870] = 16'b0000000000110110;
    assign weights2[1871] = 16'b0000000000000000;
    assign weights2[1872] = 16'b0000000000111000;
    assign weights2[1873] = 16'b0000000010001110;
    assign weights2[1874] = 16'b0000000000111110;
    assign weights2[1875] = 16'b0000000001110011;
    assign weights2[1876] = 16'b0000000000100100;
    assign weights2[1877] = 16'b0000000010100100;
    assign weights2[1878] = 16'b0000000001101010;
    assign weights2[1879] = 16'b0000000000100100;
    assign weights2[1880] = 16'b1111111111110100;
    assign weights2[1881] = 16'b1111111110101101;
    assign weights2[1882] = 16'b0000000000011010;
    assign weights2[1883] = 16'b0000000001011000;
    assign weights2[1884] = 16'b1111111111101001;
    assign weights2[1885] = 16'b1111111110010000;
    assign weights2[1886] = 16'b0000000010110100;
    assign weights2[1887] = 16'b0000000000110011;
    assign weights2[1888] = 16'b0000000000110010;
    assign weights2[1889] = 16'b0000000000100110;
    assign weights2[1890] = 16'b0000000000100010;
    assign weights2[1891] = 16'b0000000000101010;
    assign weights2[1892] = 16'b1111111111010011;
    assign weights2[1893] = 16'b0000000000101100;
    assign weights2[1894] = 16'b0000000000101110;
    assign weights2[1895] = 16'b1111111111100100;
    assign weights2[1896] = 16'b1111111111011011;
    assign weights2[1897] = 16'b1111111111101111;
    assign weights2[1898] = 16'b1111111111111000;
    assign weights2[1899] = 16'b1111111111010110;
    assign weights2[1900] = 16'b0000000000110111;
    assign weights2[1901] = 16'b1111111101110100;
    assign weights2[1902] = 16'b1111111111011011;
    assign weights2[1903] = 16'b0000000000101101;
    assign weights2[1904] = 16'b0000000000001010;
    assign weights2[1905] = 16'b0000000000101001;
    assign weights2[1906] = 16'b1111111110101111;
    assign weights2[1907] = 16'b1111111111000000;
    assign weights2[1908] = 16'b0000000000110000;
    assign weights2[1909] = 16'b1111111111111111;
    assign weights2[1910] = 16'b0000000000000000;
    assign weights2[1911] = 16'b0000000000000010;
    assign weights2[1912] = 16'b0000000000011010;
    assign weights2[1913] = 16'b1111111111010001;
    assign weights2[1914] = 16'b1111111111100011;
    assign weights2[1915] = 16'b1111111110101111;
    assign weights2[1916] = 16'b0000000000011101;
    assign weights2[1917] = 16'b1111111111011000;
    assign weights2[1918] = 16'b0000000000001010;
    assign weights2[1919] = 16'b0000000000000001;
    assign weights2[1920] = 16'b1111111111111001;
    assign weights2[1921] = 16'b0000000010111100;
    assign weights2[1922] = 16'b0000000001011010;
    assign weights2[1923] = 16'b0000000000001101;
    assign weights2[1924] = 16'b1111111111100011;
    assign weights2[1925] = 16'b0000000000011111;
    assign weights2[1926] = 16'b0000000000000000;
    assign weights2[1927] = 16'b0000000001110001;
    assign weights2[1928] = 16'b0000000000111010;
    assign weights2[1929] = 16'b1111111111101101;
    assign weights2[1930] = 16'b0000000000111011;
    assign weights2[1931] = 16'b0000000000010100;
    assign weights2[1932] = 16'b0000000010101101;
    assign weights2[1933] = 16'b0000000010001001;
    assign weights2[1934] = 16'b1111111111111010;
    assign weights2[1935] = 16'b1111111111111010;
    assign weights2[1936] = 16'b1111111111010001;
    assign weights2[1937] = 16'b0000000001001110;
    assign weights2[1938] = 16'b1111111111110110;
    assign weights2[1939] = 16'b1111111111100011;
    assign weights2[1940] = 16'b1111111110001100;
    assign weights2[1941] = 16'b0000000001010011;
    assign weights2[1942] = 16'b0000000000000001;
    assign weights2[1943] = 16'b0000000000000111;
    assign weights2[1944] = 16'b0000000000010110;
    assign weights2[1945] = 16'b0000000000001011;
    assign weights2[1946] = 16'b1111111111111110;
    assign weights2[1947] = 16'b0000000000110101;
    assign weights2[1948] = 16'b0000000010001001;
    assign weights2[1949] = 16'b0000000001001000;
    assign weights2[1950] = 16'b0000000001000010;
    assign weights2[1951] = 16'b1111111111011110;
    assign weights2[1952] = 16'b1111111111010111;
    assign weights2[1953] = 16'b1111111111111001;
    assign weights2[1954] = 16'b0000000000000010;
    assign weights2[1955] = 16'b0000000001000001;
    assign weights2[1956] = 16'b0000000001100101;
    assign weights2[1957] = 16'b1111111111101101;
    assign weights2[1958] = 16'b0000000000011101;
    assign weights2[1959] = 16'b1111111111010010;
    assign weights2[1960] = 16'b1111111111001001;
    assign weights2[1961] = 16'b1111111111101000;
    assign weights2[1962] = 16'b0000000000000101;
    assign weights2[1963] = 16'b0000000000011001;
    assign weights2[1964] = 16'b1111111111101010;
    assign weights2[1965] = 16'b0000000000011111;
    assign weights2[1966] = 16'b0000000010010010;
    assign weights2[1967] = 16'b0000000001010010;
    assign weights2[1968] = 16'b0000000000100101;
    assign weights2[1969] = 16'b0000000000101011;
    assign weights2[1970] = 16'b0000000010011110;
    assign weights2[1971] = 16'b1111111111011000;
    assign weights2[1972] = 16'b1111111111100100;
    assign weights2[1973] = 16'b1111111111001101;
    assign weights2[1974] = 16'b0000000000000000;
    assign weights2[1975] = 16'b1111111111110000;
    assign weights2[1976] = 16'b1111111111111100;
    assign weights2[1977] = 16'b0000000000011110;
    assign weights2[1978] = 16'b1111111111110001;
    assign weights2[1979] = 16'b1111111111100111;
    assign weights2[1980] = 16'b1111111111101110;
    assign weights2[1981] = 16'b0000000000011010;
    assign weights2[1982] = 16'b0000000001010100;
    assign weights2[1983] = 16'b0000000000000101;
    assign weights2[1984] = 16'b0000000000001001;
    assign weights2[1985] = 16'b1111111101101111;
    assign weights2[1986] = 16'b0000000000100110;
    assign weights2[1987] = 16'b0000000000010011;
    assign weights2[1988] = 16'b1111111110111101;
    assign weights2[1989] = 16'b0000000000101110;
    assign weights2[1990] = 16'b0000000000000000;
    assign weights2[1991] = 16'b1111111111100110;
    assign weights2[1992] = 16'b0000000000100111;
    assign weights2[1993] = 16'b1111111110110100;
    assign weights2[1994] = 16'b0000000000000110;
    assign weights2[1995] = 16'b1111111101001001;
    assign weights2[1996] = 16'b1111111111111111;
    assign weights2[1997] = 16'b1111111110100000;
    assign weights2[1998] = 16'b0000000000011111;
    assign weights2[1999] = 16'b1111111111111001;
    assign weights2[2000] = 16'b1111111110011111;
    assign weights2[2001] = 16'b0000000000100001;
    assign weights2[2002] = 16'b1111111110000101;
    assign weights2[2003] = 16'b1111111111000100;
    assign weights2[2004] = 16'b1111111111011100;
    assign weights2[2005] = 16'b0000000000111101;
    assign weights2[2006] = 16'b1111111110101100;
    assign weights2[2007] = 16'b0000000000011001;
    assign weights2[2008] = 16'b0000000000100100;
    assign weights2[2009] = 16'b0000000000110101;
    assign weights2[2010] = 16'b1111111110100101;
    assign weights2[2011] = 16'b1111111110011010;
    assign weights2[2012] = 16'b0000000000001001;
    assign weights2[2013] = 16'b0000000000111001;
    assign weights2[2014] = 16'b0000000000111100;
    assign weights2[2015] = 16'b0000000000010010;
    assign weights2[2016] = 16'b0000000000011111;
    assign weights2[2017] = 16'b1111111111000101;
    assign weights2[2018] = 16'b0000000000010110;
    assign weights2[2019] = 16'b0000000000110101;
    assign weights2[2020] = 16'b0000000000000100;
    assign weights2[2021] = 16'b0000000000010100;
    assign weights2[2022] = 16'b0000000000101101;
    assign weights2[2023] = 16'b1111111101101100;
    assign weights2[2024] = 16'b1111111101110011;
    assign weights2[2025] = 16'b1111111101001110;
    assign weights2[2026] = 16'b0000000000001001;
    assign weights2[2027] = 16'b0000000000011111;
    assign weights2[2028] = 16'b0000000000101110;
    assign weights2[2029] = 16'b0000000000111001;
    assign weights2[2030] = 16'b1111111111101100;
    assign weights2[2031] = 16'b1111111101010111;
    assign weights2[2032] = 16'b1111111111101110;
    assign weights2[2033] = 16'b0000000000110110;
    assign weights2[2034] = 16'b0000000000100100;
    assign weights2[2035] = 16'b1111111111010001;
    assign weights2[2036] = 16'b1111111111010100;
    assign weights2[2037] = 16'b1111111110000111;
    assign weights2[2038] = 16'b0000000000000000;
    assign weights2[2039] = 16'b1111111110111010;
    assign weights2[2040] = 16'b1111111110011101;
    assign weights2[2041] = 16'b0000000000100101;
    assign weights2[2042] = 16'b0000000000000111;
    assign weights2[2043] = 16'b1111111110101100;
    assign weights2[2044] = 16'b1111111110001000;
    assign weights2[2045] = 16'b0000000000111001;
    assign weights2[2046] = 16'b1111111111100111;
    assign weights2[2047] = 16'b1111111111010000;
    assign biases2[0] = 16'b0000000010000011;
    assign biases2[1] = 16'b0000000001110011;
    assign biases2[2] = 16'b0000000010001011;
    assign biases2[3] = 16'b0000000011010100;
    assign biases2[4] = 16'b0000000010101100;
    assign biases2[5] = 16'b0000000000111101;
    assign biases2[6] = 16'b0000000011111100;
    assign biases2[7] = 16'b0000000011110111;
    assign biases2[8] = 16'b0000000010110001;
    assign biases2[9] = 16'b1111111110001000;
    assign biases2[10] = 16'b0000000000100001;
    assign biases2[11] = 16'b0000000100101101;
    assign biases2[12] = 16'b1111111101101000;
    assign biases2[13] = 16'b0000000110110010;
    assign biases2[14] = 16'b0000000100000101;
    assign biases2[15] = 16'b0000000010011100;
    assign biases2[16] = 16'b0000000000010100;
    assign biases2[17] = 16'b0000000100100011;
    assign biases2[18] = 16'b1111111101111111;
    assign biases2[19] = 16'b1111111110010101;
    assign biases2[20] = 16'b0000000011101001;
    assign biases2[21] = 16'b0000000010101111;
    assign biases2[22] = 16'b0000000011010101;
    assign biases2[23] = 16'b0000000100011011;
    assign biases2[24] = 16'b1111111111010110;
    assign biases2[25] = 16'b0000000101010010;
    assign biases2[26] = 16'b0000000010000000;
    assign biases2[27] = 16'b0000000000000111;
    assign biases2[28] = 16'b0000000001011011;
    assign biases2[29] = 16'b1111111100101010;
    assign biases2[30] = 16'b1111111110011101;
    assign biases2[31] = 16'b0000000001110000;
    assign weights3[0] = 16'b0000000001111011;
    assign weights3[1] = 16'b1111111110001010;
    assign weights3[2] = 16'b0000000000111111;
    assign weights3[3] = 16'b0000000010110101;
    assign weights3[4] = 16'b1111111101101011;
    assign weights3[5] = 16'b0000000000110001;
    assign weights3[6] = 16'b0000000010011111;
    assign weights3[7] = 16'b0000000000000000;
    assign weights3[8] = 16'b1111111101101001;
    assign weights3[9] = 16'b1111111101101000;
    assign weights3[10] = 16'b1111111101111110;
    assign weights3[11] = 16'b1111111111101110;
    assign weights3[12] = 16'b0000000000010110;
    assign weights3[13] = 16'b0000000000100100;
    assign weights3[14] = 16'b0000000001100010;
    assign weights3[15] = 16'b1111111111011101;
    assign weights3[16] = 16'b1111111101001100;
    assign weights3[17] = 16'b1111111110100000;
    assign weights3[18] = 16'b0000000001001101;
    assign weights3[19] = 16'b1111111110101111;
    assign weights3[20] = 16'b0000000001000001;
    assign weights3[21] = 16'b1111111101101101;
    assign weights3[22] = 16'b0000000001000000;
    assign weights3[23] = 16'b0000000000011101;
    assign weights3[24] = 16'b0000000001000100;
    assign weights3[25] = 16'b1111111110010100;
    assign weights3[26] = 16'b1111111110100000;
    assign weights3[27] = 16'b1111111110101011;
    assign weights3[28] = 16'b1111111110101010;
    assign weights3[29] = 16'b1111111110101010;
    assign weights3[30] = 16'b1111111101111001;
    assign weights3[31] = 16'b0000000000011010;
    assign weights3[32] = 16'b1111111110000100;
    assign weights3[33] = 16'b1111111110000010;
    assign weights3[34] = 16'b0000000000100111;
    assign weights3[35] = 16'b1111111110100111;
    assign weights3[36] = 16'b0000000000110110;
    assign weights3[37] = 16'b0000000000000110;
    assign weights3[38] = 16'b1111111100000000;
    assign weights3[39] = 16'b0000000001110000;
    assign weights3[40] = 16'b1111111111100011;
    assign weights3[41] = 16'b0000000000000011;
    assign weights3[42] = 16'b1111111111011101;
    assign weights3[43] = 16'b1111111110101101;
    assign weights3[44] = 16'b0000000001001011;
    assign weights3[45] = 16'b0000000001101011;
    assign weights3[46] = 16'b1111111101101010;
    assign weights3[47] = 16'b0000000010000111;
    assign weights3[48] = 16'b0000000001001011;
    assign weights3[49] = 16'b1111111100100011;
    assign weights3[50] = 16'b0000000000000101;
    assign weights3[51] = 16'b0000000000110001;
    assign weights3[52] = 16'b0000000000011111;
    assign weights3[53] = 16'b1111111101011101;
    assign weights3[54] = 16'b1111111101111001;
    assign weights3[55] = 16'b0000000000010100;
    assign weights3[56] = 16'b0000000000110110;
    assign weights3[57] = 16'b0000000001010010;
    assign weights3[58] = 16'b0000000001000001;
    assign weights3[59] = 16'b1111111101101010;
    assign weights3[60] = 16'b0000000000001001;
    assign weights3[61] = 16'b0000000001001101;
    assign weights3[62] = 16'b0000000001011100;
    assign weights3[63] = 16'b0000000011000111;
    assign weights3[64] = 16'b0000000001001011;
    assign weights3[65] = 16'b1111111110001110;
    assign weights3[66] = 16'b0000000000101000;
    assign weights3[67] = 16'b1111111101101011;
    assign weights3[68] = 16'b1111111110011001;
    assign weights3[69] = 16'b0000000000011101;
    assign weights3[70] = 16'b1111111111011101;
    assign weights3[71] = 16'b1111111111010010;
    assign weights3[72] = 16'b1111111110101100;
    assign weights3[73] = 16'b0000000000110010;
    assign weights3[74] = 16'b0000000000110101;
    assign weights3[75] = 16'b0000000001111000;
    assign weights3[76] = 16'b0000000000001100;
    assign weights3[77] = 16'b1111111101011010;
    assign weights3[78] = 16'b1111111110111110;
    assign weights3[79] = 16'b1111111101111110;
    assign weights3[80] = 16'b1111111110100000;
    assign weights3[81] = 16'b0000000000010111;
    assign weights3[82] = 16'b0000000001000000;
    assign weights3[83] = 16'b0000000000111000;
    assign weights3[84] = 16'b1111111110001110;
    assign weights3[85] = 16'b1111111110110010;
    assign weights3[86] = 16'b1111111111111100;
    assign weights3[87] = 16'b0000000000000001;
    assign weights3[88] = 16'b0000000000110110;
    assign weights3[89] = 16'b1111111101011101;
    assign weights3[90] = 16'b1111111101100110;
    assign weights3[91] = 16'b1111111111111010;
    assign weights3[92] = 16'b0000000001001101;
    assign weights3[93] = 16'b0000000001010110;
    assign weights3[94] = 16'b0000000000000101;
    assign weights3[95] = 16'b1111111110011001;
    assign weights3[96] = 16'b1111111111000010;
    assign weights3[97] = 16'b0000000001000101;
    assign weights3[98] = 16'b0000000000110010;
    assign weights3[99] = 16'b1111111101111100;
    assign weights3[100] = 16'b1111111110110110;
    assign weights3[101] = 16'b1111111110101100;
    assign weights3[102] = 16'b1111111110111011;
    assign weights3[103] = 16'b1111111110111111;
    assign weights3[104] = 16'b0000000000110011;
    assign weights3[105] = 16'b1111111110111101;
    assign weights3[106] = 16'b0000000000110000;
    assign weights3[107] = 16'b1111111111011001;
    assign weights3[108] = 16'b1111111110110100;
    assign weights3[109] = 16'b1111111101101001;
    assign weights3[110] = 16'b1111111111011100;
    assign weights3[111] = 16'b1111111101100011;
    assign weights3[112] = 16'b0000000001000110;
    assign weights3[113] = 16'b1111111110101010;
    assign weights3[114] = 16'b0000000000111111;
    assign weights3[115] = 16'b0000000000010011;
    assign weights3[116] = 16'b1111111101101111;
    assign weights3[117] = 16'b1111111110011111;
    assign weights3[118] = 16'b0000000000110110;
    assign weights3[119] = 16'b0000000001000100;
    assign weights3[120] = 16'b1111111111001011;
    assign weights3[121] = 16'b1111111110101001;
    assign weights3[122] = 16'b0000000000111001;
    assign weights3[123] = 16'b0000000000110011;
    assign weights3[124] = 16'b0000000001001011;
    assign weights3[125] = 16'b0000000001000011;
    assign weights3[126] = 16'b0000000000100111;
    assign weights3[127] = 16'b1111111110011101;
    assign weights3[128] = 16'b1111111111011101;
    assign weights3[129] = 16'b1111111110101010;
    assign weights3[130] = 16'b1111111100011000;
    assign weights3[131] = 16'b1111111111101100;
    assign weights3[132] = 16'b0000000001010011;
    assign weights3[133] = 16'b0000000001000001;
    assign weights3[134] = 16'b0000000001100101;
    assign weights3[135] = 16'b1111111110010100;
    assign weights3[136] = 16'b1111111110000100;
    assign weights3[137] = 16'b0000000000011110;
    assign weights3[138] = 16'b1111111110100101;
    assign weights3[139] = 16'b1111111111010110;
    assign weights3[140] = 16'b0000000001000001;
    assign weights3[141] = 16'b0000000000111000;
    assign weights3[142] = 16'b1111111101111000;
    assign weights3[143] = 16'b1111111111111101;
    assign weights3[144] = 16'b0000000000011001;
    assign weights3[145] = 16'b0000000001101110;
    assign weights3[146] = 16'b1111111101110110;
    assign weights3[147] = 16'b0000000000111010;
    assign weights3[148] = 16'b1111111111010010;
    assign weights3[149] = 16'b0000000001000001;
    assign weights3[150] = 16'b1111111110001111;
    assign weights3[151] = 16'b1111111110001011;
    assign weights3[152] = 16'b0000000000111001;
    assign weights3[153] = 16'b0000000001011011;
    assign weights3[154] = 16'b0000000001001110;
    assign weights3[155] = 16'b0000000000111000;
    assign weights3[156] = 16'b1111111110000110;
    assign weights3[157] = 16'b1111111110100111;
    assign weights3[158] = 16'b1111111101011111;
    assign weights3[159] = 16'b1111111101011101;
    assign weights3[160] = 16'b1111111110111101;
    assign weights3[161] = 16'b0000000001001010;
    assign weights3[162] = 16'b1111111111111110;
    assign weights3[163] = 16'b1111111110000100;
    assign weights3[164] = 16'b1111111110100011;
    assign weights3[165] = 16'b1111111110111010;
    assign weights3[166] = 16'b1111111110110010;
    assign weights3[167] = 16'b1111111111010110;
    assign weights3[168] = 16'b0000000001010100;
    assign weights3[169] = 16'b1111111111110111;
    assign weights3[170] = 16'b0000000000101111;
    assign weights3[171] = 16'b1111111110110110;
    assign weights3[172] = 16'b0000000001000101;
    assign weights3[173] = 16'b1111111101110110;
    assign weights3[174] = 16'b0000000000111111;
    assign weights3[175] = 16'b1111111111000110;
    assign weights3[176] = 16'b0000000000111111;
    assign weights3[177] = 16'b1111111110101111;
    assign weights3[178] = 16'b0000000000101011;
    assign weights3[179] = 16'b1111111111100001;
    assign weights3[180] = 16'b0000000001010010;
    assign weights3[181] = 16'b0000000001001001;
    assign weights3[182] = 16'b0000000000110001;
    assign weights3[183] = 16'b1111111101000100;
    assign weights3[184] = 16'b1111111110101101;
    assign weights3[185] = 16'b1111111110100000;
    assign weights3[186] = 16'b1111111111001011;
    assign weights3[187] = 16'b0000000000101111;
    assign weights3[188] = 16'b1111111110101010;
    assign weights3[189] = 16'b1111111110011000;
    assign weights3[190] = 16'b0000000000110100;
    assign weights3[191] = 16'b1111111110110111;
    assign weights3[192] = 16'b0000000001011101;
    assign weights3[193] = 16'b1111111111110000;
    assign weights3[194] = 16'b1111111110011011;
    assign weights3[195] = 16'b0000000001110011;
    assign weights3[196] = 16'b1111111110001110;
    assign weights3[197] = 16'b1111111100110001;
    assign weights3[198] = 16'b0000000010000001;
    assign weights3[199] = 16'b1111111110001011;
    assign weights3[200] = 16'b0000000001001001;
    assign weights3[201] = 16'b0000000000101100;
    assign weights3[202] = 16'b1111111100100100;
    assign weights3[203] = 16'b0000000001001001;
    assign weights3[204] = 16'b0000000001000001;
    assign weights3[205] = 16'b1111111111011100;
    assign weights3[206] = 16'b1111111110111110;
    assign weights3[207] = 16'b0000000010101000;
    assign weights3[208] = 16'b1111111101111100;
    assign weights3[209] = 16'b0000000000111101;
    assign weights3[210] = 16'b1111111101001111;
    assign weights3[211] = 16'b0000000000101110;
    assign weights3[212] = 16'b0000000001100010;
    assign weights3[213] = 16'b0000000001011111;
    assign weights3[214] = 16'b0000000000101001;
    assign weights3[215] = 16'b1111111100011010;
    assign weights3[216] = 16'b0000000000110000;
    assign weights3[217] = 16'b1111111110000110;
    assign weights3[218] = 16'b1111111111101001;
    assign weights3[219] = 16'b1111111101010101;
    assign weights3[220] = 16'b1111111110001001;
    assign weights3[221] = 16'b1111111111001101;
    assign weights3[222] = 16'b0000000000101111;
    assign weights3[223] = 16'b0000000000010001;
    assign weights3[224] = 16'b1111111101110011;
    assign weights3[225] = 16'b1111111101100001;
    assign weights3[226] = 16'b0000000000110011;
    assign weights3[227] = 16'b1111111110101111;
    assign weights3[228] = 16'b0000000001100100;
    assign weights3[229] = 16'b0000000001001111;
    assign weights3[230] = 16'b1111111110000001;
    assign weights3[231] = 16'b0000000010000010;
    assign weights3[232] = 16'b1111111101111111;
    assign weights3[233] = 16'b0000000000101100;
    assign weights3[234] = 16'b0000000000101111;
    assign weights3[235] = 16'b1111111111011100;
    assign weights3[236] = 16'b0000000001000000;
    assign weights3[237] = 16'b1111111110101011;
    assign weights3[238] = 16'b0000000001010000;
    assign weights3[239] = 16'b1111111100111100;
    assign weights3[240] = 16'b0000000001010101;
    assign weights3[241] = 16'b1111111111010111;
    assign weights3[242] = 16'b0000000000111000;
    assign weights3[243] = 16'b1111111110101111;
    assign weights3[244] = 16'b1111111110001100;
    assign weights3[245] = 16'b1111111111010000;
    assign weights3[246] = 16'b1111111100111111;
    assign weights3[247] = 16'b0000000001000110;
    assign weights3[248] = 16'b1111111110101000;
    assign weights3[249] = 16'b1111111111001000;
    assign weights3[250] = 16'b1111111110001110;
    assign weights3[251] = 16'b0000000001000010;
    assign weights3[252] = 16'b0000000000110010;
    assign weights3[253] = 16'b0000000001001111;
    assign weights3[254] = 16'b1111111110001111;
    assign weights3[255] = 16'b1111111110111111;
    assign weights3[256] = 16'b1111111111101110;
    assign weights3[257] = 16'b0000000000100110;
    assign weights3[258] = 16'b0000000000101110;
    assign weights3[259] = 16'b1111111101100001;
    assign weights3[260] = 16'b1111111110011111;
    assign weights3[261] = 16'b1111111110100000;
    assign weights3[262] = 16'b1111111101111011;
    assign weights3[263] = 16'b0000000010010011;
    assign weights3[264] = 16'b0000000001000011;
    assign weights3[265] = 16'b1111111110101001;
    assign weights3[266] = 16'b1111111111111100;
    assign weights3[267] = 16'b0000000001101101;
    assign weights3[268] = 16'b1111111111010001;
    assign weights3[269] = 16'b0000000001100000;
    assign weights3[270] = 16'b0000000000111011;
    assign weights3[271] = 16'b1111111111001011;
    assign weights3[272] = 16'b1111111110111110;
    assign weights3[273] = 16'b1111111101110000;
    assign weights3[274] = 16'b1111111111000101;
    assign weights3[275] = 16'b1111111111100011;
    assign weights3[276] = 16'b0000000000111010;
    assign weights3[277] = 16'b0000000000011101;
    assign weights3[278] = 16'b0000000000010110;
    assign weights3[279] = 16'b0000000000100110;
    assign weights3[280] = 16'b1111111111001010;
    assign weights3[281] = 16'b0000000001101000;
    assign weights3[282] = 16'b0000000000010010;
    assign weights3[283] = 16'b1111111111001110;
    assign weights3[284] = 16'b0000000000110011;
    assign weights3[285] = 16'b1111111111001011;
    assign weights3[286] = 16'b1111111111001111;
    assign weights3[287] = 16'b0000000000010110;
    assign weights3[288] = 16'b1111111111101101;
    assign weights3[289] = 16'b0000000000111111;
    assign weights3[290] = 16'b1111111110010010;
    assign weights3[291] = 16'b0000000000001110;
    assign weights3[292] = 16'b0000000001010011;
    assign weights3[293] = 16'b0000000001000001;
    assign weights3[294] = 16'b0000000001101111;
    assign weights3[295] = 16'b1111111111001111;
    assign weights3[296] = 16'b1111111111001010;
    assign weights3[297] = 16'b1111111111001000;
    assign weights3[298] = 16'b0000000000100000;
    assign weights3[299] = 16'b1111111111000110;
    assign weights3[300] = 16'b1111111101110110;
    assign weights3[301] = 16'b0000000000010011;
    assign weights3[302] = 16'b0000000001001001;
    assign weights3[303] = 16'b1111111110001010;
    assign weights3[304] = 16'b0000000000111101;
    assign weights3[305] = 16'b0000000001110010;
    assign weights3[306] = 16'b0000000000000110;
    assign weights3[307] = 16'b1111111101100110;
    assign weights3[308] = 16'b1111111110111001;
    assign weights3[309] = 16'b0000000000001010;
    assign weights3[310] = 16'b1111111110000010;
    assign weights3[311] = 16'b0000000001100010;
    assign weights3[312] = 16'b1111111101110010;
    assign weights3[313] = 16'b0000000001000110;
    assign weights3[314] = 16'b0000000000011011;
    assign weights3[315] = 16'b0000000000101011;
    assign weights3[316] = 16'b1111111101011110;
    assign weights3[317] = 16'b1111111111011111;
    assign weights3[318] = 16'b1111111111011101;
    assign weights3[319] = 16'b1111111101111110;
    assign biases3[0] = 16'b0000000000000100;
    assign biases3[1] = 16'b1111111011110110;
    assign biases3[2] = 16'b0000000000011001;
    assign biases3[3] = 16'b1111111111110100;
    assign biases3[4] = 16'b0000000001000000;
    assign biases3[5] = 16'b0000000000110111;
    assign biases3[6] = 16'b1111111110001101;
    assign biases3[7] = 16'b1111111101100110;
    assign biases3[8] = 16'b0000000011001010;
    assign biases3[9] = 16'b0000000010001111;

endmodule
