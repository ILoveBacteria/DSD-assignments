//////////////////////////////////////////////////////////////////////////////////
// AXI4 Lite Slave Example
// By:
//        Ali Jahanian
// 
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps

module axi4_lite_slave #(
    parameter ADDRESS = 32,
    parameter DATA_WIDTH = 32
    )
    (
        // Global Signals
        input                           ACLK, // # of used = 1
        input                           ARESETN, // # of used = 1

        // Read Address Channel INPUTS
        input           [ADDRESS-1:0]   S_ARADDR, // # of used = 4
        input                           S_ARVALID, // # of used = 2

        // Read Data Channel INPUTS
        input                           S_RREADY, // # of used = 1

        // Write Address Channel INPUTS
        /* verilator lint_off UNUSED */
        input           [ADDRESS-1:0]   S_AWADDR, // # of used = 4
        input                           S_AWVALID, // # of used = 2

        // Write Data  Channel INPUTS
        input          [DATA_WIDTH-1:0] S_WDATA, // # of used = 2
        input          [3:0]            S_WSTRB, // # of used = 0
        input                           S_WVALID, // # of used = 1

        // Write Response Channel INPUTS
        input                           S_BREADY, // # of used = 1

        // Read Address Channel OUTPUTS
        output                     S_ARREADY, // # of used = 2

        // Read Data Channel OUTPUTS
        output [DATA_WIDTH-1:0]    S_RDATA, // # of used = 1
        output          [1:0]      S_RRESP, // # of used = 1
        output                     S_RVALID, // # of used = 2

        // Write Address Channel OUTPUTS
        output                     S_AWREADY, // # of used = 2
        output                     S_WREADY, // # of used = 2
        
        // Write Response Channel OUTPUTS
        output          [1:0]      S_BRESP, // # of used = 1
        output                     S_BVALID // # of used = 2
    );

    localparam REG_NUM       = 32;
    localparam IDLE          = 0;
    localparam WRITE_CHANNEL = 1;
    localparam WRESP_CHANNEL = 2;
    localparam RADDR_CHANNEL = 3;
    localparam RDATA_CHANNEL = 4;
    localparam MY_STATE      = 5;

    reg start;
    wire clk;
    reg rst;
    reg [783:0] in_features;
    reg [783:0] not_reversed_in_features;
    wire [3:0] prediction;
    wire done;

    NeuralNetwork my_NeuralNetwork (clk, rst, start, in_features, prediction, done);

    assign clk = ACLK;
   
    reg  [2:0] state, next_state;
    reg  [ADDRESS-1:0] read_addr;
    wire [ADDRESS-1:0] S_ARADDR_T;
    wire [ADDRESS-1:0] S_AWADDR_T;
    reg  [DATA_WIDTH-1:0] register [0:REG_NUM-1]; // 32 ta register 32bits
    
    // Address Read
    assign S_ARREADY = (state == RADDR_CHANNEL) ? 1 : 0;
    
    // Read
    assign S_RVALID = (state == RDATA_CHANNEL) ? 1 : 0;
    assign S_RDATA  = (state == RDATA_CHANNEL) ? register[read_addr] : 0;
    assign S_RRESP  = (state == RDATA_CHANNEL) ? 2'b00 : 0;

    // Address Write
    assign S_AWREADY = (state == WRITE_CHANNEL) ? 1 : 0;

    // Write
    assign S_WREADY = (state == WRITE_CHANNEL) ? 1 : 0;

    // Response
    assign S_BVALID = (state == WRESP_CHANNEL) ? 1 : 0;
    assign S_BRESP  = (state == WRESP_CHANNEL )? 0:0;

    assign S_ARADDR_T = S_ARADDR[ADDRESS-1:2]; // Read address 
    assign S_AWADDR_T = S_AWADDR[ADDRESS-1:2]; // Write address 
    
    always @(posedge ACLK) begin
        // Reset the register array
        if (~ARESETN) begin
            state <= IDLE;
        end
        else begin
            state <= next_state;
            if (state == WRITE_CHANNEL) begin
                register[S_AWADDR_T] <= S_WDATA;
            end
            else if (state == RADDR_CHANNEL) begin
                read_addr <= S_ARADDR_T;
            end
            else if (state == IDLE) begin
                start <= 0;
                rst <= 1;
            end
            else if (state == MY_STATE) begin
                start <= 1;
                rst <= 0;
                in_features = {register[23], register[22], register[21], register[20], register[19], register[18], register[17], register[16], register[15], register[14], register[13], register[12], register[11], register[10], register[9], register[8], register[7], register[6], register[5], register[4], register[3], register[2], register[1], register[0]};
                // in_features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000011111100000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000000000000000000101111111000000000000000000010100000111000000000000000001110000000110000000000000000110000000001000000000000000011000000000100000000000000000100000000010000000000000000010000000001000000000000000000110000001000000000000000000001111111000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                register[24] <= {28'h0000000, prediction};
            end
        end
    end

    // State machine
    always @(*) begin
        next_state = state;
        case (state)
            IDLE: begin
                if (S_AWVALID) begin
                    next_state = WRITE_CHANNEL;
                end 
                else if (S_ARVALID) begin
                    next_state = RADDR_CHANNEL;
                end 
                else begin
                    next_state = IDLE;
                end
            end

            RADDR_CHANNEL: begin
                if (S_ARVALID && S_ARREADY && S_ARADDR_T == 24)
                    next_state = MY_STATE;
                else if (S_ARVALID && S_ARREADY)
                    next_state = RDATA_CHANNEL;
            end

            MY_STATE: begin
                if (done)
                    next_state = RDATA_CHANNEL;
            end

            RDATA_CHANNEL: begin
                if (S_RVALID && S_RREADY)
                    next_state = IDLE;
            end

            WRITE_CHANNEL: begin
                if (S_AWVALID && S_AWREADY && S_WREADY && S_WVALID)
                    next_state = WRESP_CHANNEL;
            end

            WRESP_CHANNEL: begin
                if (S_BVALID && S_BREADY) 
                    next_state = IDLE;
            end

            default: begin
                next_state = IDLE;
            end 
        endcase
    end
endmodule

module NeuralNetwork (
    input clk,
    input rst,
    input start,
    input [783:0] in_features, // 784 input features
    output reg [3:0] prediction, // 10 output classes (ArgMax index)
    output reg done
);

    // register to hold the input features
    reg [783:0] features;

    // state machine
    localparam IDLE = 0, COMPUTE = 1;
    reg state;
    reg [2:0] count_clocks; 

    // Define the parameters for layer sizes
    parameter INPUT_SIZE = 784;
    parameter HIDDEN1_SIZE = 64;
    parameter HIDDEN2_SIZE = 32;
    parameter OUTPUT_SIZE = 10;
    
    // Define memory for weights and biases (assumed preloaded)
    (* ram_style = "block" *) reg signed [15:0] weights1 [0:50175];
    (* ram_style = "block" *) reg signed [15:0] biases1 [0:63];
    
    (* ram_style = "block" *) reg signed [15:0] weights2 [0:2047];
    (* ram_style = "block" *) reg signed [15:0] biases2 [0:31];
    
    (* ram_style = "block" *) reg signed [15:0] weights3 [0:319];
    (* ram_style = "block" *) reg signed [15:0] biases3 [0:9];

    // Layer Outputs
    reg signed [15:0] hidden1 [0:HIDDEN1_SIZE-1];
    reg signed [15:0] hidden2 [0:HIDDEN2_SIZE-1];
    reg signed [15:0] output_layer [0:OUTPUT_SIZE-1];
    
    // ReLU activation function
    function signed [15:0] relu;
        input signed [15:0] x;
        begin
            relu = (x > 0) ? x : 0;
        end
    endfunction

    integer i, j;

    // ============================================
    // combinational Computation of the neurons
    // ============================================

    // layer 1
    reg signed [15:0] new_hidden1 [0:HIDDEN1_SIZE-1];
    always @(*) begin
        for (i = 0; i < HIDDEN1_SIZE; i = i + 1) begin
            new_hidden1[i] = biases1[i];
            for (j = 0; j < INPUT_SIZE; j = j + 1) begin
                new_hidden1[i] = new_hidden1[i] + (features[j] == 1 ? weights1[i*INPUT_SIZE+j] : 0); 
            end
            new_hidden1[i] = relu(new_hidden1[i]); 
        end
    end

    // layer 2
    reg signed [15:0] new_hidden2 [0:HIDDEN2_SIZE-1];
    reg signed [31:0] multiplier_out2 [0:HIDDEN2_SIZE-1][0:HIDDEN1_SIZE-1];
    reg signed [15:0] shift_out2 [0:HIDDEN2_SIZE-1][0:HIDDEN1_SIZE-1];
    always @(*) begin
        for (i = 0; i < HIDDEN2_SIZE; i = i + 1) begin
            new_hidden2[i] = biases2[i];
            for (j = 0; j < HIDDEN1_SIZE; j = j + 1) begin
                multiplier_out2[i][j] = hidden1[j] * weights2[i*HIDDEN1_SIZE+j];
                shift_out2[i][j] = multiplier_out2[i][j] >> 8;
                new_hidden2[i] = new_hidden2[i] + shift_out2[i][j];
            end
            new_hidden2[i] = relu(new_hidden2[i]);
        end
    end

    // Output Layer computation
    reg signed [15:0] new_output_layer [0:OUTPUT_SIZE-1];
    reg signed [31:0] multiplier_out3 [0:OUTPUT_SIZE-1][0:HIDDEN2_SIZE-1];
    reg signed [15:0] shift_out3 [0:OUTPUT_SIZE-1][0:HIDDEN2_SIZE-1];
    always @(*) begin
        for (i = 0; i < OUTPUT_SIZE; i = i + 1) begin
            new_output_layer[i] = biases3[i];
            for (j = 0; j < HIDDEN2_SIZE; j = j + 1) begin
                multiplier_out3[i][j] = hidden2[j] * weights3[i*HIDDEN2_SIZE+j];
                shift_out3[i][j] = multiplier_out3[i][j] >> 8;
                new_output_layer[i] = new_output_layer[i] + shift_out3[i][j];
            end
        end
    end

    // ArgMax operation
    reg [3:0] new_prediction;
    always @(*) begin
        new_prediction = 0;
        for (i = 1; i < OUTPUT_SIZE; i = i + 1) begin
            if (output_layer[i] > output_layer[new_prediction]) begin
                new_prediction = i;
            end
        end
    end
    

    // ============================================
    // Sequential update of the neurons
    // ============================================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            done <= 0;
            count_clocks <= 0;
            prediction <= 0;
            for (i = 0; i < INPUT_SIZE; i = i + 1) begin
                features[i] <= 0;
            end
        end 
        else if (state == IDLE) begin
            if (start) begin
                // Load the input features
                for (i = 0; i < INPUT_SIZE; i = i + 1) begin
                    features[i] <= in_features[i];
                end
                state <= COMPUTE;
                done <= 0;
                count_clocks <= 0;
            end
        end 
        else begin
            // Layer 1 computation
            for (i = 0; i < HIDDEN1_SIZE; i = i + 1) begin
                hidden1[i] <= new_hidden1[i];
            end

            // Layer 2 computation
            for (i = 0; i < HIDDEN2_SIZE; i = i + 1) begin
                hidden2[i] <= new_hidden2[i];
            end

            // Output Layer computation
            for (i = 0; i < OUTPUT_SIZE; i = i + 1) begin
                output_layer[i] <= new_output_layer[i];
            end

            // ArgMax operation
            prediction <= new_prediction;

            // Update state or increment the clock counter
            if (count_clocks >= 3) begin
                state <= IDLE;
                done <= 1;
            end
            else begin
                count_clocks <= count_clocks + 1;
            end
        end
    end

    
    always @(posedge clk) begin
        weights1[0] <= 16'b0000000000000000;
        weights1[1] <= 16'b0000000000000000;
        weights1[2] <= 16'b0000000000000000;
        weights1[3] <= 16'b0000000000000000;
        weights1[4] <= 16'b0000000000001100;
        weights1[5] <= 16'b0000000000011010;
        weights1[6] <= 16'b0000000000100111;
        weights1[7] <= 16'b0000000000101010;
        weights1[8] <= 16'b0000000000111110;
        weights1[9] <= 16'b0000000001001001;
        weights1[10] <= 16'b0000000000111111;
        weights1[11] <= 16'b0000000001000001;
        weights1[12] <= 16'b0000000000110011;
        weights1[13] <= 16'b0000000000100101;
        weights1[14] <= 16'b0000000000100000;
        weights1[15] <= 16'b0000000000011110;
        weights1[16] <= 16'b0000000000000110;
        weights1[17] <= 16'b0000000000000101;
        weights1[18] <= 16'b0000000000011001;
        weights1[19] <= 16'b1111111111110101;
        weights1[20] <= 16'b0000000000000011;
        weights1[21] <= 16'b0000000000000011;
        weights1[22] <= 16'b0000000000001111;
        weights1[23] <= 16'b1111111111110101;
        weights1[24] <= 16'b1111111111101011;
        weights1[25] <= 16'b1111111111101100;
        weights1[26] <= 16'b1111111111110100;
        weights1[27] <= 16'b1111111111111010;
        weights1[28] <= 16'b0000000000000000;
        weights1[29] <= 16'b0000000000000000;
        weights1[30] <= 16'b0000000000000000;
        weights1[31] <= 16'b0000000000001010;
        weights1[32] <= 16'b0000000000010101;
        weights1[33] <= 16'b0000000000100100;
        weights1[34] <= 16'b0000000000101010;
        weights1[35] <= 16'b0000000001000010;
        weights1[36] <= 16'b0000000001010011;
        weights1[37] <= 16'b0000000001000111;
        weights1[38] <= 16'b0000000001010010;
        weights1[39] <= 16'b0000000001011010;
        weights1[40] <= 16'b0000000001001000;
        weights1[41] <= 16'b0000000000101000;
        weights1[42] <= 16'b0000000000100111;
        weights1[43] <= 16'b0000000000011010;
        weights1[44] <= 16'b0000000000011110;
        weights1[45] <= 16'b0000000000011100;
        weights1[46] <= 16'b0000000000000010;
        weights1[47] <= 16'b0000000000000110;
        weights1[48] <= 16'b1111111111110111;
        weights1[49] <= 16'b0000000000010000;
        weights1[50] <= 16'b0000000000001010;
        weights1[51] <= 16'b0000000000000110;
        weights1[52] <= 16'b1111111111111001;
        weights1[53] <= 16'b1111111111111010;
        weights1[54] <= 16'b1111111111110000;
        weights1[55] <= 16'b1111111111101110;
        weights1[56] <= 16'b0000000000000000;
        weights1[57] <= 16'b0000000000000000;
        weights1[58] <= 16'b0000000000000111;
        weights1[59] <= 16'b0000000000001110;
        weights1[60] <= 16'b0000000000011000;
        weights1[61] <= 16'b0000000000011101;
        weights1[62] <= 16'b0000000000100100;
        weights1[63] <= 16'b0000000000110001;
        weights1[64] <= 16'b0000000000111101;
        weights1[65] <= 16'b0000000001000101;
        weights1[66] <= 16'b0000000001001001;
        weights1[67] <= 16'b0000000001000110;
        weights1[68] <= 16'b0000000001001101;
        weights1[69] <= 16'b0000000001000010;
        weights1[70] <= 16'b0000000000101111;
        weights1[71] <= 16'b0000000000011111;
        weights1[72] <= 16'b0000000000101100;
        weights1[73] <= 16'b0000000000100100;
        weights1[74] <= 16'b0000000000001111;
        weights1[75] <= 16'b0000000000001000;
        weights1[76] <= 16'b0000000000010000;
        weights1[77] <= 16'b0000000000011110;
        weights1[78] <= 16'b0000000000000100;
        weights1[79] <= 16'b0000000000000110;
        weights1[80] <= 16'b0000000000001111;
        weights1[81] <= 16'b1111111111110010;
        weights1[82] <= 16'b1111111111110110;
        weights1[83] <= 16'b1111111111110010;
        weights1[84] <= 16'b0000000000000000;
        weights1[85] <= 16'b0000000000000011;
        weights1[86] <= 16'b0000000000001001;
        weights1[87] <= 16'b0000000000010000;
        weights1[88] <= 16'b0000000000011000;
        weights1[89] <= 16'b0000000000010111;
        weights1[90] <= 16'b0000000000010111;
        weights1[91] <= 16'b0000000000101100;
        weights1[92] <= 16'b0000000000110001;
        weights1[93] <= 16'b0000000000111101;
        weights1[94] <= 16'b0000000000111111;
        weights1[95] <= 16'b0000000001000101;
        weights1[96] <= 16'b0000000001010111;
        weights1[97] <= 16'b0000000001010101;
        weights1[98] <= 16'b0000000001001001;
        weights1[99] <= 16'b0000000000110110;
        weights1[100] <= 16'b0000000000010010;
        weights1[101] <= 16'b0000000000101000;
        weights1[102] <= 16'b0000000000011111;
        weights1[103] <= 16'b0000000000011110;
        weights1[104] <= 16'b0000000000010100;
        weights1[105] <= 16'b0000000000010000;
        weights1[106] <= 16'b0000000000011001;
        weights1[107] <= 16'b0000000000001001;
        weights1[108] <= 16'b0000000000000110;
        weights1[109] <= 16'b0000000000000100;
        weights1[110] <= 16'b1111111111111000;
        weights1[111] <= 16'b1111111111101010;
        weights1[112] <= 16'b0000000000000011;
        weights1[113] <= 16'b0000000000000101;
        weights1[114] <= 16'b1111111111111101;
        weights1[115] <= 16'b1111111111110111;
        weights1[116] <= 16'b1111111111110100;
        weights1[117] <= 16'b1111111111110100;
        weights1[118] <= 16'b1111111111111101;
        weights1[119] <= 16'b0000000000000111;
        weights1[120] <= 16'b0000000000100010;
        weights1[121] <= 16'b0000000000011101;
        weights1[122] <= 16'b0000000000101010;
        weights1[123] <= 16'b0000000001000011;
        weights1[124] <= 16'b0000000000110111;
        weights1[125] <= 16'b0000000001100100;
        weights1[126] <= 16'b0000000001100000;
        weights1[127] <= 16'b0000000001001000;
        weights1[128] <= 16'b0000000000110101;
        weights1[129] <= 16'b0000000000100110;
        weights1[130] <= 16'b0000000000011101;
        weights1[131] <= 16'b0000000000010110;
        weights1[132] <= 16'b0000000000010101;
        weights1[133] <= 16'b0000000000001110;
        weights1[134] <= 16'b0000000000010001;
        weights1[135] <= 16'b0000000000010001;
        weights1[136] <= 16'b0000000000001001;
        weights1[137] <= 16'b0000000000000100;
        weights1[138] <= 16'b0000000000001011;
        weights1[139] <= 16'b1111111111110111;
        weights1[140] <= 16'b1111111111111110;
        weights1[141] <= 16'b1111111111110011;
        weights1[142] <= 16'b1111111111101111;
        weights1[143] <= 16'b1111111111100000;
        weights1[144] <= 16'b1111111111010010;
        weights1[145] <= 16'b1111111111001110;
        weights1[146] <= 16'b1111111111010011;
        weights1[147] <= 16'b1111111111100001;
        weights1[148] <= 16'b1111111111010101;
        weights1[149] <= 16'b1111111111001011;
        weights1[150] <= 16'b1111111111101000;
        weights1[151] <= 16'b1111111111101011;
        weights1[152] <= 16'b0000000000010001;
        weights1[153] <= 16'b0000000000110111;
        weights1[154] <= 16'b0000000001000111;
        weights1[155] <= 16'b0000000001010110;
        weights1[156] <= 16'b0000000001010001;
        weights1[157] <= 16'b0000000001000100;
        weights1[158] <= 16'b0000000000100011;
        weights1[159] <= 16'b0000000000010011;
        weights1[160] <= 16'b0000000000101100;
        weights1[161] <= 16'b0000000000100010;
        weights1[162] <= 16'b0000000000011100;
        weights1[163] <= 16'b0000000000011011;
        weights1[164] <= 16'b0000000000010010;
        weights1[165] <= 16'b0000000000010001;
        weights1[166] <= 16'b0000000000010010;
        weights1[167] <= 16'b1111111111111101;
        weights1[168] <= 16'b1111111111111000;
        weights1[169] <= 16'b1111111111100110;
        weights1[170] <= 16'b1111111111001101;
        weights1[171] <= 16'b1111111110111011;
        weights1[172] <= 16'b1111111110100110;
        weights1[173] <= 16'b1111111110011111;
        weights1[174] <= 16'b1111111110100100;
        weights1[175] <= 16'b1111111110101001;
        weights1[176] <= 16'b1111111110011100;
        weights1[177] <= 16'b1111111110011100;
        weights1[178] <= 16'b1111111110011011;
        weights1[179] <= 16'b1111111110111111;
        weights1[180] <= 16'b1111111110100111;
        weights1[181] <= 16'b1111111111000111;
        weights1[182] <= 16'b1111111111101011;
        weights1[183] <= 16'b0000000000100111;
        weights1[184] <= 16'b0000000000111101;
        weights1[185] <= 16'b0000000001000101;
        weights1[186] <= 16'b0000000000101111;
        weights1[187] <= 16'b0000000000101010;
        weights1[188] <= 16'b0000000000011100;
        weights1[189] <= 16'b0000000000010110;
        weights1[190] <= 16'b0000000000100100;
        weights1[191] <= 16'b0000000000001001;
        weights1[192] <= 16'b0000000000010110;
        weights1[193] <= 16'b0000000000011101;
        weights1[194] <= 16'b0000000000001011;
        weights1[195] <= 16'b0000000000001110;
        weights1[196] <= 16'b1111111111110110;
        weights1[197] <= 16'b1111111111001110;
        weights1[198] <= 16'b1111111110110101;
        weights1[199] <= 16'b1111111110011010;
        weights1[200] <= 16'b1111111101110101;
        weights1[201] <= 16'b1111111101110010;
        weights1[202] <= 16'b1111111110000001;
        weights1[203] <= 16'b1111111110000011;
        weights1[204] <= 16'b1111111101101011;
        weights1[205] <= 16'b1111111101110101;
        weights1[206] <= 16'b1111111101101110;
        weights1[207] <= 16'b1111111110010001;
        weights1[208] <= 16'b1111111110001010;
        weights1[209] <= 16'b1111111110001111;
        weights1[210] <= 16'b1111111110100011;
        weights1[211] <= 16'b1111111111001001;
        weights1[212] <= 16'b1111111111111110;
        weights1[213] <= 16'b0000000000101100;
        weights1[214] <= 16'b0000000000101111;
        weights1[215] <= 16'b0000000000101100;
        weights1[216] <= 16'b0000000000101010;
        weights1[217] <= 16'b0000000000101110;
        weights1[218] <= 16'b0000000000100000;
        weights1[219] <= 16'b0000000000100111;
        weights1[220] <= 16'b0000000000101011;
        weights1[221] <= 16'b0000000000010110;
        weights1[222] <= 16'b0000000000001001;
        weights1[223] <= 16'b0000000000010101;
        weights1[224] <= 16'b1111111111101001;
        weights1[225] <= 16'b1111111111000010;
        weights1[226] <= 16'b1111111110100101;
        weights1[227] <= 16'b1111111110010100;
        weights1[228] <= 16'b1111111101111001;
        weights1[229] <= 16'b1111111101110111;
        weights1[230] <= 16'b1111111101111100;
        weights1[231] <= 16'b1111111110001101;
        weights1[232] <= 16'b1111111101111111;
        weights1[233] <= 16'b1111111110000110;
        weights1[234] <= 16'b1111111110110010;
        weights1[235] <= 16'b1111111110101101;
        weights1[236] <= 16'b1111111111001010;
        weights1[237] <= 16'b1111111110111001;
        weights1[238] <= 16'b1111111111001001;
        weights1[239] <= 16'b1111111110111011;
        weights1[240] <= 16'b1111111111001101;
        weights1[241] <= 16'b1111111111111110;
        weights1[242] <= 16'b0000000000011001;
        weights1[243] <= 16'b0000000000101111;
        weights1[244] <= 16'b0000000000000011;
        weights1[245] <= 16'b0000000000110010;
        weights1[246] <= 16'b0000000000010110;
        weights1[247] <= 16'b0000000000011010;
        weights1[248] <= 16'b0000000000010100;
        weights1[249] <= 16'b0000000000000011;
        weights1[250] <= 16'b0000000000100000;
        weights1[251] <= 16'b0000000000001111;
        weights1[252] <= 16'b1111111111101000;
        weights1[253] <= 16'b1111111111000111;
        weights1[254] <= 16'b1111111110101101;
        weights1[255] <= 16'b1111111110011111;
        weights1[256] <= 16'b1111111110100010;
        weights1[257] <= 16'b1111111110100000;
        weights1[258] <= 16'b1111111110110010;
        weights1[259] <= 16'b1111111110110011;
        weights1[260] <= 16'b1111111110100101;
        weights1[261] <= 16'b1111111111100101;
        weights1[262] <= 16'b1111111111011010;
        weights1[263] <= 16'b1111111111101110;
        weights1[264] <= 16'b1111111111101000;
        weights1[265] <= 16'b1111111111100011;
        weights1[266] <= 16'b1111111111001011;
        weights1[267] <= 16'b1111111111001000;
        weights1[268] <= 16'b1111111111001101;
        weights1[269] <= 16'b1111111111100100;
        weights1[270] <= 16'b1111111111101010;
        weights1[271] <= 16'b0000000000000010;
        weights1[272] <= 16'b0000000000000001;
        weights1[273] <= 16'b0000000000011001;
        weights1[274] <= 16'b0000000000100100;
        weights1[275] <= 16'b0000000000011101;
        weights1[276] <= 16'b0000000000010000;
        weights1[277] <= 16'b0000000000010001;
        weights1[278] <= 16'b0000000000010100;
        weights1[279] <= 16'b0000000000010010;
        weights1[280] <= 16'b1111111111111100;
        weights1[281] <= 16'b1111111111101010;
        weights1[282] <= 16'b1111111111011001;
        weights1[283] <= 16'b1111111111100010;
        weights1[284] <= 16'b1111111111110000;
        weights1[285] <= 16'b0000000000000010;
        weights1[286] <= 16'b0000000000000101;
        weights1[287] <= 16'b0000000000000000;
        weights1[288] <= 16'b0000000000010010;
        weights1[289] <= 16'b0000000000011001;
        weights1[290] <= 16'b1111111111111101;
        weights1[291] <= 16'b1111111111101111;
        weights1[292] <= 16'b1111111111110011;
        weights1[293] <= 16'b1111111111101111;
        weights1[294] <= 16'b1111111111100110;
        weights1[295] <= 16'b1111111111110001;
        weights1[296] <= 16'b1111111111011010;
        weights1[297] <= 16'b1111111111011101;
        weights1[298] <= 16'b1111111111011101;
        weights1[299] <= 16'b1111111111100111;
        weights1[300] <= 16'b1111111111101100;
        weights1[301] <= 16'b0000000000000101;
        weights1[302] <= 16'b0000000000011001;
        weights1[303] <= 16'b0000000000011100;
        weights1[304] <= 16'b0000000000011001;
        weights1[305] <= 16'b0000000000011000;
        weights1[306] <= 16'b0000000000011010;
        weights1[307] <= 16'b0000000000011100;
        weights1[308] <= 16'b0000000000001000;
        weights1[309] <= 16'b0000000000010011;
        weights1[310] <= 16'b0000000000100010;
        weights1[311] <= 16'b0000000000101011;
        weights1[312] <= 16'b0000000000110011;
        weights1[313] <= 16'b0000000000111001;
        weights1[314] <= 16'b0000000001000100;
        weights1[315] <= 16'b0000000000101111;
        weights1[316] <= 16'b0000000000011111;
        weights1[317] <= 16'b0000000000010101;
        weights1[318] <= 16'b0000000000001010;
        weights1[319] <= 16'b1111111111111011;
        weights1[320] <= 16'b1111111111101111;
        weights1[321] <= 16'b1111111111111000;
        weights1[322] <= 16'b1111111111100000;
        weights1[323] <= 16'b1111111111100101;
        weights1[324] <= 16'b1111111111111010;
        weights1[325] <= 16'b1111111111110011;
        weights1[326] <= 16'b1111111111100001;
        weights1[327] <= 16'b1111111111110000;
        weights1[328] <= 16'b1111111111101010;
        weights1[329] <= 16'b0000000000000001;
        weights1[330] <= 16'b0000000000010000;
        weights1[331] <= 16'b0000000000001001;
        weights1[332] <= 16'b0000000000001101;
        weights1[333] <= 16'b0000000000011100;
        weights1[334] <= 16'b0000000000011101;
        weights1[335] <= 16'b0000000000001100;
        weights1[336] <= 16'b0000000000011011;
        weights1[337] <= 16'b0000000000101001;
        weights1[338] <= 16'b0000000000110111;
        weights1[339] <= 16'b0000000000111101;
        weights1[340] <= 16'b0000000000111010;
        weights1[341] <= 16'b0000000000100001;
        weights1[342] <= 16'b0000000000010100;
        weights1[343] <= 16'b1111111111101110;
        weights1[344] <= 16'b0000000000001110;
        weights1[345] <= 16'b0000000000000000;
        weights1[346] <= 16'b1111111111110000;
        weights1[347] <= 16'b0000000000000001;
        weights1[348] <= 16'b1111111111110111;
        weights1[349] <= 16'b1111111111110000;
        weights1[350] <= 16'b1111111111101011;
        weights1[351] <= 16'b1111111111110111;
        weights1[352] <= 16'b1111111111101010;
        weights1[353] <= 16'b1111111111110101;
        weights1[354] <= 16'b1111111111101011;
        weights1[355] <= 16'b1111111111101100;
        weights1[356] <= 16'b1111111111111000;
        weights1[357] <= 16'b1111111111110010;
        weights1[358] <= 16'b0000000000000010;
        weights1[359] <= 16'b0000000000001100;
        weights1[360] <= 16'b0000000000010100;
        weights1[361] <= 16'b0000000000000111;
        weights1[362] <= 16'b0000000000010100;
        weights1[363] <= 16'b0000000000010011;
        weights1[364] <= 16'b0000000000101101;
        weights1[365] <= 16'b0000000000101011;
        weights1[366] <= 16'b0000000000110110;
        weights1[367] <= 16'b0000000000111000;
        weights1[368] <= 16'b0000000000101100;
        weights1[369] <= 16'b0000000000001110;
        weights1[370] <= 16'b0000000000000111;
        weights1[371] <= 16'b0000000000000001;
        weights1[372] <= 16'b0000000000001011;
        weights1[373] <= 16'b1111111111110111;
        weights1[374] <= 16'b0000000000011010;
        weights1[375] <= 16'b1111111111111010;
        weights1[376] <= 16'b1111111111110010;
        weights1[377] <= 16'b1111111111101110;
        weights1[378] <= 16'b1111111111011000;
        weights1[379] <= 16'b1111111111110101;
        weights1[380] <= 16'b1111111111101000;
        weights1[381] <= 16'b1111111111110000;
        weights1[382] <= 16'b1111111111100110;
        weights1[383] <= 16'b1111111111111111;
        weights1[384] <= 16'b1111111111110000;
        weights1[385] <= 16'b1111111111101111;
        weights1[386] <= 16'b0000000000001010;
        weights1[387] <= 16'b1111111111110111;
        weights1[388] <= 16'b1111111111111101;
        weights1[389] <= 16'b0000000000001110;
        weights1[390] <= 16'b0000000000000101;
        weights1[391] <= 16'b0000000000010011;
        weights1[392] <= 16'b0000000000110010;
        weights1[393] <= 16'b0000000000010010;
        weights1[394] <= 16'b0000000000011110;
        weights1[395] <= 16'b0000000000010011;
        weights1[396] <= 16'b0000000000001000;
        weights1[397] <= 16'b0000000000010000;
        weights1[398] <= 16'b0000000000000011;
        weights1[399] <= 16'b0000000000010010;
        weights1[400] <= 16'b1111111111111000;
        weights1[401] <= 16'b0000000000000111;
        weights1[402] <= 16'b0000000000000010;
        weights1[403] <= 16'b0000000000001111;
        weights1[404] <= 16'b0000000000000101;
        weights1[405] <= 16'b1111111111111111;
        weights1[406] <= 16'b0000000000000011;
        weights1[407] <= 16'b1111111111100110;
        weights1[408] <= 16'b1111111111111011;
        weights1[409] <= 16'b1111111111111100;
        weights1[410] <= 16'b1111111111100100;
        weights1[411] <= 16'b1111111111111000;
        weights1[412] <= 16'b1111111111101011;
        weights1[413] <= 16'b1111111111110110;
        weights1[414] <= 16'b0000000000000001;
        weights1[415] <= 16'b0000000000010000;
        weights1[416] <= 16'b1111111111111110;
        weights1[417] <= 16'b1111111111101000;
        weights1[418] <= 16'b1111111111111101;
        weights1[419] <= 16'b0000000000011011;
        weights1[420] <= 16'b0000000000010001;
        weights1[421] <= 16'b0000000000010101;
        weights1[422] <= 16'b1111111111111111;
        weights1[423] <= 16'b0000000000010100;
        weights1[424] <= 16'b1111111111110110;
        weights1[425] <= 16'b0000000000000001;
        weights1[426] <= 16'b0000000000001101;
        weights1[427] <= 16'b1111111111110011;
        weights1[428] <= 16'b0000000000010011;
        weights1[429] <= 16'b1111111111111100;
        weights1[430] <= 16'b0000000000001000;
        weights1[431] <= 16'b0000000000000111;
        weights1[432] <= 16'b0000000000000001;
        weights1[433] <= 16'b0000000000000000;
        weights1[434] <= 16'b1111111111110001;
        weights1[435] <= 16'b1111111111101110;
        weights1[436] <= 16'b1111111111111100;
        weights1[437] <= 16'b1111111111101101;
        weights1[438] <= 16'b1111111111101111;
        weights1[439] <= 16'b1111111111110010;
        weights1[440] <= 16'b1111111111111100;
        weights1[441] <= 16'b0000000000001001;
        weights1[442] <= 16'b1111111111111111;
        weights1[443] <= 16'b1111111111111010;
        weights1[444] <= 16'b0000000000001111;
        weights1[445] <= 16'b0000000000001001;
        weights1[446] <= 16'b0000000000000110;
        weights1[447] <= 16'b0000000000100111;
        weights1[448] <= 16'b0000000000010001;
        weights1[449] <= 16'b0000000000001100;
        weights1[450] <= 16'b1111111111110001;
        weights1[451] <= 16'b0000000000000001;
        weights1[452] <= 16'b1111111111111011;
        weights1[453] <= 16'b0000000000010110;
        weights1[454] <= 16'b1111111111111100;
        weights1[455] <= 16'b0000000000010000;
        weights1[456] <= 16'b0000000000000101;
        weights1[457] <= 16'b0000000000001110;
        weights1[458] <= 16'b0000000000000001;
        weights1[459] <= 16'b0000000000001001;
        weights1[460] <= 16'b0000000000000011;
        weights1[461] <= 16'b0000000000000101;
        weights1[462] <= 16'b1111111111111111;
        weights1[463] <= 16'b0000000000001101;
        weights1[464] <= 16'b1111111111100100;
        weights1[465] <= 16'b0000000000000100;
        weights1[466] <= 16'b1111111111101101;
        weights1[467] <= 16'b1111111111101111;
        weights1[468] <= 16'b1111111111110001;
        weights1[469] <= 16'b1111111111110110;
        weights1[470] <= 16'b1111111111111001;
        weights1[471] <= 16'b1111111111110010;
        weights1[472] <= 16'b1111111111101000;
        weights1[473] <= 16'b0000000000000100;
        weights1[474] <= 16'b0000000000000110;
        weights1[475] <= 16'b0000000000100101;
        weights1[476] <= 16'b0000000000000101;
        weights1[477] <= 16'b0000000000010001;
        weights1[478] <= 16'b0000000000001110;
        weights1[479] <= 16'b1111111111110000;
        weights1[480] <= 16'b0000000000001000;
        weights1[481] <= 16'b0000000000000011;
        weights1[482] <= 16'b0000000000010000;
        weights1[483] <= 16'b0000000000001001;
        weights1[484] <= 16'b0000000000011001;
        weights1[485] <= 16'b0000000000000000;
        weights1[486] <= 16'b0000000000000111;
        weights1[487] <= 16'b0000000000001101;
        weights1[488] <= 16'b1111111111110110;
        weights1[489] <= 16'b0000000000000111;
        weights1[490] <= 16'b1111111111111100;
        weights1[491] <= 16'b1111111111110110;
        weights1[492] <= 16'b1111111111111001;
        weights1[493] <= 16'b1111111111101101;
        weights1[494] <= 16'b1111111111111011;
        weights1[495] <= 16'b1111111111111001;
        weights1[496] <= 16'b1111111111101100;
        weights1[497] <= 16'b1111111111110010;
        weights1[498] <= 16'b1111111111101101;
        weights1[499] <= 16'b1111111111110001;
        weights1[500] <= 16'b1111111111111010;
        weights1[501] <= 16'b0000000000001100;
        weights1[502] <= 16'b0000000000010110;
        weights1[503] <= 16'b0000000000011110;
        weights1[504] <= 16'b0000000000001100;
        weights1[505] <= 16'b0000000000010001;
        weights1[506] <= 16'b0000000000000001;
        weights1[507] <= 16'b1111111111111111;
        weights1[508] <= 16'b1111111111111010;
        weights1[509] <= 16'b0000000000010101;
        weights1[510] <= 16'b0000000000000101;
        weights1[511] <= 16'b1111111111101001;
        weights1[512] <= 16'b0000000000011100;
        weights1[513] <= 16'b0000000000000001;
        weights1[514] <= 16'b1111111111111001;
        weights1[515] <= 16'b0000000000001001;
        weights1[516] <= 16'b0000000000001111;
        weights1[517] <= 16'b1111111111110101;
        weights1[518] <= 16'b1111111111110010;
        weights1[519] <= 16'b1111111111100100;
        weights1[520] <= 16'b1111111111110110;
        weights1[521] <= 16'b1111111111110111;
        weights1[522] <= 16'b1111111111110011;
        weights1[523] <= 16'b1111111111111000;
        weights1[524] <= 16'b1111111111100110;
        weights1[525] <= 16'b0000000000000101;
        weights1[526] <= 16'b1111111111111101;
        weights1[527] <= 16'b0000000000011100;
        weights1[528] <= 16'b0000000000010101;
        weights1[529] <= 16'b1111111111111100;
        weights1[530] <= 16'b0000000000000001;
        weights1[531] <= 16'b0000000000010011;
        weights1[532] <= 16'b0000000000010001;
        weights1[533] <= 16'b0000000000010001;
        weights1[534] <= 16'b0000000000001100;
        weights1[535] <= 16'b1111111111110101;
        weights1[536] <= 16'b0000000000000001;
        weights1[537] <= 16'b0000000000010101;
        weights1[538] <= 16'b0000000000001011;
        weights1[539] <= 16'b0000000000000100;
        weights1[540] <= 16'b0000000000001110;
        weights1[541] <= 16'b0000000000000100;
        weights1[542] <= 16'b0000000000000001;
        weights1[543] <= 16'b0000000000000100;
        weights1[544] <= 16'b0000000000001010;
        weights1[545] <= 16'b0000000000001011;
        weights1[546] <= 16'b1111111111101110;
        weights1[547] <= 16'b0000000000000100;
        weights1[548] <= 16'b1111111111110101;
        weights1[549] <= 16'b1111111111110010;
        weights1[550] <= 16'b1111111111111111;
        weights1[551] <= 16'b0000000000000100;
        weights1[552] <= 16'b1111111111111110;
        weights1[553] <= 16'b1111111111101101;
        weights1[554] <= 16'b0000000000000000;
        weights1[555] <= 16'b1111111111100111;
        weights1[556] <= 16'b0000000000000000;
        weights1[557] <= 16'b1111111111110001;
        weights1[558] <= 16'b0000000000001000;
        weights1[559] <= 16'b0000000000001110;
        weights1[560] <= 16'b0000000000000101;
        weights1[561] <= 16'b0000000000001100;
        weights1[562] <= 16'b0000000000001010;
        weights1[563] <= 16'b0000000000001100;
        weights1[564] <= 16'b0000000000000011;
        weights1[565] <= 16'b0000000000001000;
        weights1[566] <= 16'b0000000000001011;
        weights1[567] <= 16'b0000000000001100;
        weights1[568] <= 16'b1111111111111110;
        weights1[569] <= 16'b0000000000001101;
        weights1[570] <= 16'b1111111111111011;
        weights1[571] <= 16'b0000000000000001;
        weights1[572] <= 16'b1111111111111110;
        weights1[573] <= 16'b0000000000000100;
        weights1[574] <= 16'b1111111111110000;
        weights1[575] <= 16'b0000000000000010;
        weights1[576] <= 16'b1111111111111101;
        weights1[577] <= 16'b1111111111101101;
        weights1[578] <= 16'b1111111111111110;
        weights1[579] <= 16'b1111111111111100;
        weights1[580] <= 16'b1111111111101110;
        weights1[581] <= 16'b0000000000001100;
        weights1[582] <= 16'b1111111111100010;
        weights1[583] <= 16'b1111111111101000;
        weights1[584] <= 16'b1111111111110000;
        weights1[585] <= 16'b1111111111101111;
        weights1[586] <= 16'b1111111111111011;
        weights1[587] <= 16'b0000000000000011;
        weights1[588] <= 16'b0000000000000010;
        weights1[589] <= 16'b0000000000001010;
        weights1[590] <= 16'b0000000000000100;
        weights1[591] <= 16'b0000000000001011;
        weights1[592] <= 16'b1111111111111010;
        weights1[593] <= 16'b1111111111111000;
        weights1[594] <= 16'b0000000000000010;
        weights1[595] <= 16'b1111111111110100;
        weights1[596] <= 16'b1111111111111110;
        weights1[597] <= 16'b0000000000001001;
        weights1[598] <= 16'b0000000000000011;
        weights1[599] <= 16'b1111111111101110;
        weights1[600] <= 16'b1111111111110011;
        weights1[601] <= 16'b1111111111111100;
        weights1[602] <= 16'b0000000000000011;
        weights1[603] <= 16'b1111111111110101;
        weights1[604] <= 16'b1111111111111111;
        weights1[605] <= 16'b1111111111111001;
        weights1[606] <= 16'b1111111111110111;
        weights1[607] <= 16'b0000000000000100;
        weights1[608] <= 16'b1111111111111110;
        weights1[609] <= 16'b0000000000010001;
        weights1[610] <= 16'b1111111111111110;
        weights1[611] <= 16'b1111111111111100;
        weights1[612] <= 16'b1111111111110011;
        weights1[613] <= 16'b1111111111110011;
        weights1[614] <= 16'b1111111111111000;
        weights1[615] <= 16'b0000000000000001;
        weights1[616] <= 16'b1111111111111110;
        weights1[617] <= 16'b0000000000000100;
        weights1[618] <= 16'b0000000000000101;
        weights1[619] <= 16'b0000000000000111;
        weights1[620] <= 16'b0000000000001000;
        weights1[621] <= 16'b1111111111111100;
        weights1[622] <= 16'b0000000000000101;
        weights1[623] <= 16'b0000000000100001;
        weights1[624] <= 16'b1111111111110001;
        weights1[625] <= 16'b0000000000000011;
        weights1[626] <= 16'b1111111111110001;
        weights1[627] <= 16'b1111111111111101;
        weights1[628] <= 16'b1111111111111100;
        weights1[629] <= 16'b1111111111101111;
        weights1[630] <= 16'b0000000000000010;
        weights1[631] <= 16'b1111111111100010;
        weights1[632] <= 16'b0000000000000110;
        weights1[633] <= 16'b0000000000001011;
        weights1[634] <= 16'b0000000000001000;
        weights1[635] <= 16'b1111111111111011;
        weights1[636] <= 16'b1111111111111110;
        weights1[637] <= 16'b0000000000001000;
        weights1[638] <= 16'b0000000000000000;
        weights1[639] <= 16'b0000000000000000;
        weights1[640] <= 16'b1111111111110100;
        weights1[641] <= 16'b1111111111111100;
        weights1[642] <= 16'b1111111111111100;
        weights1[643] <= 16'b1111111111110110;
        weights1[644] <= 16'b0000000000000010;
        weights1[645] <= 16'b0000000000000001;
        weights1[646] <= 16'b1111111111111101;
        weights1[647] <= 16'b1111111111110110;
        weights1[648] <= 16'b1111111111111001;
        weights1[649] <= 16'b0000000000000001;
        weights1[650] <= 16'b1111111111111010;
        weights1[651] <= 16'b1111111111110101;
        weights1[652] <= 16'b1111111111111100;
        weights1[653] <= 16'b1111111111110001;
        weights1[654] <= 16'b0000000000000101;
        weights1[655] <= 16'b1111111111111000;
        weights1[656] <= 16'b0000000000000101;
        weights1[657] <= 16'b1111111111100010;
        weights1[658] <= 16'b1111111111011100;
        weights1[659] <= 16'b0000000000000101;
        weights1[660] <= 16'b1111111111111011;
        weights1[661] <= 16'b1111111111110110;
        weights1[662] <= 16'b1111111111111111;
        weights1[663] <= 16'b0000000000010101;
        weights1[664] <= 16'b1111111111110001;
        weights1[665] <= 16'b0000000000000010;
        weights1[666] <= 16'b0000000000000101;
        weights1[667] <= 16'b1111111111111101;
        weights1[668] <= 16'b1111111111110010;
        weights1[669] <= 16'b1111111111110101;
        weights1[670] <= 16'b1111111111110100;
        weights1[671] <= 16'b1111111111111001;
        weights1[672] <= 16'b1111111111111011;
        weights1[673] <= 16'b1111111111111101;
        weights1[674] <= 16'b1111111111111011;
        weights1[675] <= 16'b1111111111111010;
        weights1[676] <= 16'b1111111111110001;
        weights1[677] <= 16'b1111111111110110;
        weights1[678] <= 16'b1111111111101000;
        weights1[679] <= 16'b1111111111011100;
        weights1[680] <= 16'b0000000000001110;
        weights1[681] <= 16'b1111111111011001;
        weights1[682] <= 16'b1111111111111101;
        weights1[683] <= 16'b1111111111111010;
        weights1[684] <= 16'b0000000000000011;
        weights1[685] <= 16'b0000000000010000;
        weights1[686] <= 16'b1111111111111101;
        weights1[687] <= 16'b1111111111111111;
        weights1[688] <= 16'b1111111111111111;
        weights1[689] <= 16'b1111111111110011;
        weights1[690] <= 16'b0000000000000111;
        weights1[691] <= 16'b0000000000000100;
        weights1[692] <= 16'b1111111111111010;
        weights1[693] <= 16'b0000000000000011;
        weights1[694] <= 16'b0000000000000110;
        weights1[695] <= 16'b0000000000000011;
        weights1[696] <= 16'b1111111111110110;
        weights1[697] <= 16'b1111111111111001;
        weights1[698] <= 16'b1111111111111101;
        weights1[699] <= 16'b0000000000000000;
        weights1[700] <= 16'b1111111111111110;
        weights1[701] <= 16'b0000000000000000;
        weights1[702] <= 16'b0000000000000100;
        weights1[703] <= 16'b1111111111111101;
        weights1[704] <= 16'b1111111111111010;
        weights1[705] <= 16'b1111111111101101;
        weights1[706] <= 16'b1111111111101111;
        weights1[707] <= 16'b1111111111110101;
        weights1[708] <= 16'b1111111111110111;
        weights1[709] <= 16'b0000000000000000;
        weights1[710] <= 16'b0000000000000001;
        weights1[711] <= 16'b0000000000010000;
        weights1[712] <= 16'b0000000000000101;
        weights1[713] <= 16'b1111111111111001;
        weights1[714] <= 16'b0000000000001010;
        weights1[715] <= 16'b1111111111111001;
        weights1[716] <= 16'b1111111111110100;
        weights1[717] <= 16'b1111111111011010;
        weights1[718] <= 16'b1111111111110011;
        weights1[719] <= 16'b0000000000000001;
        weights1[720] <= 16'b1111111111111111;
        weights1[721] <= 16'b1111111111110111;
        weights1[722] <= 16'b1111111111111110;
        weights1[723] <= 16'b0000000000000000;
        weights1[724] <= 16'b0000000000000100;
        weights1[725] <= 16'b1111111111111111;
        weights1[726] <= 16'b1111111111111111;
        weights1[727] <= 16'b0000000000000100;
        weights1[728] <= 16'b0000000000000000;
        weights1[729] <= 16'b0000000000000010;
        weights1[730] <= 16'b0000000000000001;
        weights1[731] <= 16'b1111111111111100;
        weights1[732] <= 16'b1111111111111010;
        weights1[733] <= 16'b1111111111110110;
        weights1[734] <= 16'b0000000000000110;
        weights1[735] <= 16'b1111111111111001;
        weights1[736] <= 16'b0000000000000011;
        weights1[737] <= 16'b0000000000000001;
        weights1[738] <= 16'b0000000000000110;
        weights1[739] <= 16'b1111111111110100;
        weights1[740] <= 16'b0000000000000011;
        weights1[741] <= 16'b0000000000000001;
        weights1[742] <= 16'b0000000000000100;
        weights1[743] <= 16'b1111111111111010;
        weights1[744] <= 16'b1111111111110111;
        weights1[745] <= 16'b1111111111110000;
        weights1[746] <= 16'b1111111111101011;
        weights1[747] <= 16'b1111111111110010;
        weights1[748] <= 16'b1111111111111110;
        weights1[749] <= 16'b1111111111111001;
        weights1[750] <= 16'b1111111111110001;
        weights1[751] <= 16'b1111111111110111;
        weights1[752] <= 16'b1111111111111011;
        weights1[753] <= 16'b1111111111111010;
        weights1[754] <= 16'b1111111111111100;
        weights1[755] <= 16'b0000000000000001;
        weights1[756] <= 16'b0000000000000000;
        weights1[757] <= 16'b0000000000000000;
        weights1[758] <= 16'b1111111111111101;
        weights1[759] <= 16'b1111111111111111;
        weights1[760] <= 16'b1111111111111010;
        weights1[761] <= 16'b1111111111111000;
        weights1[762] <= 16'b1111111111111111;
        weights1[763] <= 16'b1111111111111110;
        weights1[764] <= 16'b0000000000001001;
        weights1[765] <= 16'b1111111111110111;
        weights1[766] <= 16'b1111111111111110;
        weights1[767] <= 16'b0000000000000111;
        weights1[768] <= 16'b0000000000000100;
        weights1[769] <= 16'b1111111111110100;
        weights1[770] <= 16'b0000000000000011;
        weights1[771] <= 16'b1111111111111101;
        weights1[772] <= 16'b1111111111111001;
        weights1[773] <= 16'b1111111111111000;
        weights1[774] <= 16'b1111111111101001;
        weights1[775] <= 16'b1111111111110101;
        weights1[776] <= 16'b1111111111101110;
        weights1[777] <= 16'b1111111111111001;
        weights1[778] <= 16'b1111111111111011;
        weights1[779] <= 16'b1111111111111100;
        weights1[780] <= 16'b1111111111111011;
        weights1[781] <= 16'b1111111111111110;
        weights1[782] <= 16'b1111111111111111;
        weights1[783] <= 16'b0000000000000000;
        weights1[784] <= 16'b0000000000000000;
        weights1[785] <= 16'b0000000000000000;
        weights1[786] <= 16'b1111111111111110;
        weights1[787] <= 16'b1111111111111111;
        weights1[788] <= 16'b0000000000000000;
        weights1[789] <= 16'b1111111111111110;
        weights1[790] <= 16'b0000000000000001;
        weights1[791] <= 16'b1111111111111000;
        weights1[792] <= 16'b0000000000000000;
        weights1[793] <= 16'b1111111111110110;
        weights1[794] <= 16'b1111111111110001;
        weights1[795] <= 16'b1111111111101100;
        weights1[796] <= 16'b1111111111101010;
        weights1[797] <= 16'b1111111111101101;
        weights1[798] <= 16'b1111111111111010;
        weights1[799] <= 16'b1111111111110101;
        weights1[800] <= 16'b1111111111110000;
        weights1[801] <= 16'b1111111111101100;
        weights1[802] <= 16'b1111111111110101;
        weights1[803] <= 16'b1111111111111001;
        weights1[804] <= 16'b0000000000000011;
        weights1[805] <= 16'b0000000000000010;
        weights1[806] <= 16'b0000000000000011;
        weights1[807] <= 16'b0000000000000011;
        weights1[808] <= 16'b1111111111111111;
        weights1[809] <= 16'b0000000000000000;
        weights1[810] <= 16'b1111111111111110;
        weights1[811] <= 16'b0000000000000000;
        weights1[812] <= 16'b0000000000000000;
        weights1[813] <= 16'b0000000000000000;
        weights1[814] <= 16'b0000000000000010;
        weights1[815] <= 16'b0000000000000001;
        weights1[816] <= 16'b0000000000000100;
        weights1[817] <= 16'b0000000000000110;
        weights1[818] <= 16'b0000000000000110;
        weights1[819] <= 16'b1111111111111110;
        weights1[820] <= 16'b0000000000001011;
        weights1[821] <= 16'b1111111111111011;
        weights1[822] <= 16'b1111111111111000;
        weights1[823] <= 16'b0000000000000001;
        weights1[824] <= 16'b1111111111111000;
        weights1[825] <= 16'b1111111111111011;
        weights1[826] <= 16'b1111111111111100;
        weights1[827] <= 16'b0000000000000100;
        weights1[828] <= 16'b1111111111101100;
        weights1[829] <= 16'b1111111111111000;
        weights1[830] <= 16'b1111111111101111;
        weights1[831] <= 16'b0000000000000011;
        weights1[832] <= 16'b1111111111111101;
        weights1[833] <= 16'b1111111111111110;
        weights1[834] <= 16'b0000000000001101;
        weights1[835] <= 16'b0000000000001001;
        weights1[836] <= 16'b1111111111111111;
        weights1[837] <= 16'b1111111111110011;
        weights1[838] <= 16'b1111111111111100;
        weights1[839] <= 16'b0000000000000000;
        weights1[840] <= 16'b0000000000000000;
        weights1[841] <= 16'b1111111111111111;
        weights1[842] <= 16'b0000000000000011;
        weights1[843] <= 16'b1111111111111011;
        weights1[844] <= 16'b0000000000000111;
        weights1[845] <= 16'b0000000000000011;
        weights1[846] <= 16'b1111111111111011;
        weights1[847] <= 16'b0000000000001000;
        weights1[848] <= 16'b1111111111110110;
        weights1[849] <= 16'b1111111111111100;
        weights1[850] <= 16'b1111111111111111;
        weights1[851] <= 16'b1111111111111111;
        weights1[852] <= 16'b0000000000010111;
        weights1[853] <= 16'b0000000000001011;
        weights1[854] <= 16'b0000000000000010;
        weights1[855] <= 16'b0000000000000001;
        weights1[856] <= 16'b0000000000001000;
        weights1[857] <= 16'b1111111111101010;
        weights1[858] <= 16'b0000000000001010;
        weights1[859] <= 16'b1111111111111101;
        weights1[860] <= 16'b0000000000001010;
        weights1[861] <= 16'b0000000000000000;
        weights1[862] <= 16'b0000000000000000;
        weights1[863] <= 16'b0000000000000010;
        weights1[864] <= 16'b0000000000000011;
        weights1[865] <= 16'b1111111111111010;
        weights1[866] <= 16'b1111111111111001;
        weights1[867] <= 16'b0000000000000000;
        weights1[868] <= 16'b0000000000000000;
        weights1[869] <= 16'b0000000000000001;
        weights1[870] <= 16'b1111111111111010;
        weights1[871] <= 16'b1111111111111011;
        weights1[872] <= 16'b1111111111111110;
        weights1[873] <= 16'b0000000000000100;
        weights1[874] <= 16'b0000000000000000;
        weights1[875] <= 16'b0000000000000111;
        weights1[876] <= 16'b1111111111111001;
        weights1[877] <= 16'b0000000000000011;
        weights1[878] <= 16'b1111111111111011;
        weights1[879] <= 16'b1111111111111110;
        weights1[880] <= 16'b1111111111110111;
        weights1[881] <= 16'b0000000000001011;
        weights1[882] <= 16'b0000000000000110;
        weights1[883] <= 16'b1111111111111001;
        weights1[884] <= 16'b0000000000000010;
        weights1[885] <= 16'b0000000000010010;
        weights1[886] <= 16'b1111111111111111;
        weights1[887] <= 16'b1111111111111011;
        weights1[888] <= 16'b1111111111111011;
        weights1[889] <= 16'b1111111111110111;
        weights1[890] <= 16'b0000000000000110;
        weights1[891] <= 16'b1111111111110111;
        weights1[892] <= 16'b1111111111110101;
        weights1[893] <= 16'b0000000000000001;
        weights1[894] <= 16'b0000000000001011;
        weights1[895] <= 16'b0000000000000111;
        weights1[896] <= 16'b1111111111111110;
        weights1[897] <= 16'b1111111111110111;
        weights1[898] <= 16'b1111111111111001;
        weights1[899] <= 16'b1111111111110101;
        weights1[900] <= 16'b1111111111111101;
        weights1[901] <= 16'b1111111111111000;
        weights1[902] <= 16'b0000000000000100;
        weights1[903] <= 16'b0000000000010101;
        weights1[904] <= 16'b0000000000000101;
        weights1[905] <= 16'b0000000000010000;
        weights1[906] <= 16'b0000000000001100;
        weights1[907] <= 16'b0000000000000011;
        weights1[908] <= 16'b0000000000010110;
        weights1[909] <= 16'b1111111111110011;
        weights1[910] <= 16'b1111111111111100;
        weights1[911] <= 16'b0000000000001100;
        weights1[912] <= 16'b1111111111110101;
        weights1[913] <= 16'b0000000000001010;
        weights1[914] <= 16'b1111111111101100;
        weights1[915] <= 16'b1111111111111110;
        weights1[916] <= 16'b0000000000010000;
        weights1[917] <= 16'b1111111111110000;
        weights1[918] <= 16'b1111111111110010;
        weights1[919] <= 16'b1111111111110101;
        weights1[920] <= 16'b1111111111111010;
        weights1[921] <= 16'b0000000000000101;
        weights1[922] <= 16'b0000000000001000;
        weights1[923] <= 16'b0000000000000100;
        weights1[924] <= 16'b1111111111111100;
        weights1[925] <= 16'b1111111111111101;
        weights1[926] <= 16'b1111111111111010;
        weights1[927] <= 16'b1111111111111010;
        weights1[928] <= 16'b1111111111111010;
        weights1[929] <= 16'b1111111111111100;
        weights1[930] <= 16'b0000000000011010;
        weights1[931] <= 16'b0000000000010000;
        weights1[932] <= 16'b0000000000000101;
        weights1[933] <= 16'b0000000000001011;
        weights1[934] <= 16'b1111111111111000;
        weights1[935] <= 16'b0000000000001001;
        weights1[936] <= 16'b1111111111111111;
        weights1[937] <= 16'b0000000000000111;
        weights1[938] <= 16'b0000000000001101;
        weights1[939] <= 16'b1111111111110101;
        weights1[940] <= 16'b1111111111111111;
        weights1[941] <= 16'b0000000000000110;
        weights1[942] <= 16'b0000000000001000;
        weights1[943] <= 16'b0000000000001000;
        weights1[944] <= 16'b0000000000001011;
        weights1[945] <= 16'b0000000000000110;
        weights1[946] <= 16'b1111111111111111;
        weights1[947] <= 16'b0000000000000000;
        weights1[948] <= 16'b0000000000001111;
        weights1[949] <= 16'b1111111111111101;
        weights1[950] <= 16'b0000000000010111;
        weights1[951] <= 16'b0000000000001001;
        weights1[952] <= 16'b0000000000000001;
        weights1[953] <= 16'b0000000000001101;
        weights1[954] <= 16'b0000000000010111;
        weights1[955] <= 16'b0000000000001001;
        weights1[956] <= 16'b0000000000000011;
        weights1[957] <= 16'b1111111111111001;
        weights1[958] <= 16'b1111111111110101;
        weights1[959] <= 16'b0000000000000001;
        weights1[960] <= 16'b0000000000001101;
        weights1[961] <= 16'b0000000000000010;
        weights1[962] <= 16'b0000000000001001;
        weights1[963] <= 16'b0000000000001000;
        weights1[964] <= 16'b0000000000000100;
        weights1[965] <= 16'b1111111111111010;
        weights1[966] <= 16'b0000000000000111;
        weights1[967] <= 16'b0000000000000101;
        weights1[968] <= 16'b0000000000010000;
        weights1[969] <= 16'b1111111111111000;
        weights1[970] <= 16'b0000000000001011;
        weights1[971] <= 16'b1111111111100101;
        weights1[972] <= 16'b0000000000010000;
        weights1[973] <= 16'b1111111111101101;
        weights1[974] <= 16'b0000000000011010;
        weights1[975] <= 16'b0000000000001110;
        weights1[976] <= 16'b0000000000001100;
        weights1[977] <= 16'b0000000000000001;
        weights1[978] <= 16'b1111111111111001;
        weights1[979] <= 16'b0000000000001001;
        weights1[980] <= 16'b0000000000001000;
        weights1[981] <= 16'b1111111111111101;
        weights1[982] <= 16'b1111111111111001;
        weights1[983] <= 16'b1111111111111011;
        weights1[984] <= 16'b0000000000000011;
        weights1[985] <= 16'b1111111111111111;
        weights1[986] <= 16'b0000000000010100;
        weights1[987] <= 16'b0000000000000101;
        weights1[988] <= 16'b0000000000010001;
        weights1[989] <= 16'b1111111111111101;
        weights1[990] <= 16'b0000000000000000;
        weights1[991] <= 16'b1111111111111111;
        weights1[992] <= 16'b0000000000000100;
        weights1[993] <= 16'b0000000000010101;
        weights1[994] <= 16'b0000000000001110;
        weights1[995] <= 16'b1111111111111011;
        weights1[996] <= 16'b0000000000000101;
        weights1[997] <= 16'b1111111111111110;
        weights1[998] <= 16'b1111111111111110;
        weights1[999] <= 16'b0000000000000011;
        weights1[1000] <= 16'b0000000000001011;
        weights1[1001] <= 16'b0000000000001110;
        weights1[1002] <= 16'b0000000000000110;
        weights1[1003] <= 16'b1111111111111011;
        weights1[1004] <= 16'b1111111111110100;
        weights1[1005] <= 16'b0000000000000000;
        weights1[1006] <= 16'b0000000000000011;
        weights1[1007] <= 16'b0000000000000011;
        weights1[1008] <= 16'b0000000000000100;
        weights1[1009] <= 16'b0000000000000110;
        weights1[1010] <= 16'b1111111111111101;
        weights1[1011] <= 16'b0000000000000000;
        weights1[1012] <= 16'b1111111111111110;
        weights1[1013] <= 16'b0000000000001000;
        weights1[1014] <= 16'b1111111111110100;
        weights1[1015] <= 16'b0000000000000000;
        weights1[1016] <= 16'b0000000000000100;
        weights1[1017] <= 16'b0000000000001000;
        weights1[1018] <= 16'b1111111111111101;
        weights1[1019] <= 16'b0000000000001111;
        weights1[1020] <= 16'b1111111111111100;
        weights1[1021] <= 16'b0000000000000011;
        weights1[1022] <= 16'b0000000000000001;
        weights1[1023] <= 16'b1111111111111011;
        weights1[1024] <= 16'b0000000000001101;
        weights1[1025] <= 16'b0000000000010000;
        weights1[1026] <= 16'b0000000000010111;
        weights1[1027] <= 16'b0000000000000110;
        weights1[1028] <= 16'b1111111111100110;
        weights1[1029] <= 16'b0000000000000100;
        weights1[1030] <= 16'b1111111111111001;
        weights1[1031] <= 16'b1111111111110011;
        weights1[1032] <= 16'b0000000000000100;
        weights1[1033] <= 16'b0000000000000011;
        weights1[1034] <= 16'b1111111111110110;
        weights1[1035] <= 16'b0000000000001110;
        weights1[1036] <= 16'b0000000000000001;
        weights1[1037] <= 16'b1111111111111111;
        weights1[1038] <= 16'b1111111111111010;
        weights1[1039] <= 16'b0000000000001100;
        weights1[1040] <= 16'b0000000000010110;
        weights1[1041] <= 16'b0000000000000010;
        weights1[1042] <= 16'b0000000000000100;
        weights1[1043] <= 16'b0000000000010001;
        weights1[1044] <= 16'b1111111111101001;
        weights1[1045] <= 16'b1111111111111000;
        weights1[1046] <= 16'b0000000000000111;
        weights1[1047] <= 16'b0000000000001111;
        weights1[1048] <= 16'b0000000000010000;
        weights1[1049] <= 16'b0000000000010011;
        weights1[1050] <= 16'b0000000000000110;
        weights1[1051] <= 16'b0000000000001101;
        weights1[1052] <= 16'b1111111111110101;
        weights1[1053] <= 16'b1111111111111110;
        weights1[1054] <= 16'b0000000000000111;
        weights1[1055] <= 16'b0000000000001011;
        weights1[1056] <= 16'b0000000000000000;
        weights1[1057] <= 16'b1111111111110100;
        weights1[1058] <= 16'b1111111111111110;
        weights1[1059] <= 16'b1111111111111101;
        weights1[1060] <= 16'b1111111111101011;
        weights1[1061] <= 16'b1111111111111101;
        weights1[1062] <= 16'b0000000000000100;
        weights1[1063] <= 16'b1111111111110111;
        weights1[1064] <= 16'b0000000000001000;
        weights1[1065] <= 16'b0000000000011101;
        weights1[1066] <= 16'b0000000000001001;
        weights1[1067] <= 16'b0000000000011000;
        weights1[1068] <= 16'b1111111111111100;
        weights1[1069] <= 16'b1111111111111111;
        weights1[1070] <= 16'b0000000000000001;
        weights1[1071] <= 16'b0000000000000100;
        weights1[1072] <= 16'b0000000000001010;
        weights1[1073] <= 16'b1111111111110111;
        weights1[1074] <= 16'b1111111111111111;
        weights1[1075] <= 16'b0000000000000001;
        weights1[1076] <= 16'b0000000000001110;
        weights1[1077] <= 16'b1111111111110000;
        weights1[1078] <= 16'b0000000000000000;
        weights1[1079] <= 16'b0000000000000000;
        weights1[1080] <= 16'b1111111111111001;
        weights1[1081] <= 16'b1111111111111011;
        weights1[1082] <= 16'b1111111111111100;
        weights1[1083] <= 16'b1111111111110011;
        weights1[1084] <= 16'b0000000000010010;
        weights1[1085] <= 16'b1111111111111111;
        weights1[1086] <= 16'b1111111111110100;
        weights1[1087] <= 16'b1111111111111101;
        weights1[1088] <= 16'b0000000000000001;
        weights1[1089] <= 16'b0000000000000100;
        weights1[1090] <= 16'b0000000000000010;
        weights1[1091] <= 16'b0000000000001010;
        weights1[1092] <= 16'b1111111111111011;
        weights1[1093] <= 16'b0000000000001000;
        weights1[1094] <= 16'b1111111111110111;
        weights1[1095] <= 16'b1111111111111111;
        weights1[1096] <= 16'b0000000000010010;
        weights1[1097] <= 16'b1111111111111010;
        weights1[1098] <= 16'b1111111111111001;
        weights1[1099] <= 16'b1111111111111001;
        weights1[1100] <= 16'b1111111111111000;
        weights1[1101] <= 16'b0000000000000001;
        weights1[1102] <= 16'b0000000000010001;
        weights1[1103] <= 16'b1111111111101100;
        weights1[1104] <= 16'b1111111111111110;
        weights1[1105] <= 16'b0000000000000011;
        weights1[1106] <= 16'b1111111111110111;
        weights1[1107] <= 16'b1111111111111010;
        weights1[1108] <= 16'b1111111111110100;
        weights1[1109] <= 16'b1111111111111000;
        weights1[1110] <= 16'b0000000000001001;
        weights1[1111] <= 16'b0000000000000111;
        weights1[1112] <= 16'b1111111111111000;
        weights1[1113] <= 16'b1111111111111100;
        weights1[1114] <= 16'b0000000000010011;
        weights1[1115] <= 16'b1111111111111011;
        weights1[1116] <= 16'b1111111111110000;
        weights1[1117] <= 16'b1111111111111100;
        weights1[1118] <= 16'b0000000000000001;
        weights1[1119] <= 16'b0000000000000110;
        weights1[1120] <= 16'b1111111111110000;
        weights1[1121] <= 16'b1111111111111010;
        weights1[1122] <= 16'b1111111111111101;
        weights1[1123] <= 16'b0000000000000000;
        weights1[1124] <= 16'b0000000000000100;
        weights1[1125] <= 16'b1111111111111011;
        weights1[1126] <= 16'b1111111111111110;
        weights1[1127] <= 16'b1111111111101111;
        weights1[1128] <= 16'b1111111111110001;
        weights1[1129] <= 16'b1111111111111000;
        weights1[1130] <= 16'b1111111111101110;
        weights1[1131] <= 16'b1111111111111101;
        weights1[1132] <= 16'b1111111111110110;
        weights1[1133] <= 16'b0000000000000011;
        weights1[1134] <= 16'b1111111111111110;
        weights1[1135] <= 16'b1111111111111110;
        weights1[1136] <= 16'b1111111111111100;
        weights1[1137] <= 16'b0000000000000000;
        weights1[1138] <= 16'b1111111111110100;
        weights1[1139] <= 16'b1111111111100101;
        weights1[1140] <= 16'b1111111111111001;
        weights1[1141] <= 16'b1111111111111101;
        weights1[1142] <= 16'b0000000000000010;
        weights1[1143] <= 16'b1111111111111110;
        weights1[1144] <= 16'b0000000000000010;
        weights1[1145] <= 16'b1111111111110000;
        weights1[1146] <= 16'b1111111111111100;
        weights1[1147] <= 16'b1111111111111011;
        weights1[1148] <= 16'b1111111111100100;
        weights1[1149] <= 16'b1111111111100110;
        weights1[1150] <= 16'b1111111111101110;
        weights1[1151] <= 16'b1111111111111111;
        weights1[1152] <= 16'b0000000000001011;
        weights1[1153] <= 16'b0000000000001110;
        weights1[1154] <= 16'b1111111111111101;
        weights1[1155] <= 16'b1111111111110001;
        weights1[1156] <= 16'b1111111111110110;
        weights1[1157] <= 16'b0000000000010110;
        weights1[1158] <= 16'b1111111111110001;
        weights1[1159] <= 16'b0000000000001010;
        weights1[1160] <= 16'b0000000000011110;
        weights1[1161] <= 16'b0000000000011000;
        weights1[1162] <= 16'b0000000000010110;
        weights1[1163] <= 16'b0000000000001100;
        weights1[1164] <= 16'b0000000000001001;
        weights1[1165] <= 16'b0000000000001001;
        weights1[1166] <= 16'b1111111111111101;
        weights1[1167] <= 16'b1111111111111101;
        weights1[1168] <= 16'b1111111111111001;
        weights1[1169] <= 16'b1111111111100010;
        weights1[1170] <= 16'b1111111111111100;
        weights1[1171] <= 16'b1111111111110011;
        weights1[1172] <= 16'b0000000000000111;
        weights1[1173] <= 16'b0000000000000111;
        weights1[1174] <= 16'b1111111111110110;
        weights1[1175] <= 16'b1111111111111010;
        weights1[1176] <= 16'b1111111111011001;
        weights1[1177] <= 16'b1111111110111111;
        weights1[1178] <= 16'b1111111111010001;
        weights1[1179] <= 16'b1111111111100000;
        weights1[1180] <= 16'b0000000000000111;
        weights1[1181] <= 16'b0000000000010001;
        weights1[1182] <= 16'b0000000000011101;
        weights1[1183] <= 16'b0000000000010110;
        weights1[1184] <= 16'b0000000000100010;
        weights1[1185] <= 16'b0000000000010000;
        weights1[1186] <= 16'b0000000000000000;
        weights1[1187] <= 16'b0000000000001011;
        weights1[1188] <= 16'b0000000000011001;
        weights1[1189] <= 16'b0000000000010101;
        weights1[1190] <= 16'b0000000000001011;
        weights1[1191] <= 16'b0000000000010010;
        weights1[1192] <= 16'b0000000000000001;
        weights1[1193] <= 16'b1111111111101001;
        weights1[1194] <= 16'b0000000000000101;
        weights1[1195] <= 16'b0000000000000010;
        weights1[1196] <= 16'b1111111111111101;
        weights1[1197] <= 16'b0000000000001011;
        weights1[1198] <= 16'b1111111111100111;
        weights1[1199] <= 16'b1111111111110010;
        weights1[1200] <= 16'b0000000000001110;
        weights1[1201] <= 16'b1111111111111010;
        weights1[1202] <= 16'b1111111111110100;
        weights1[1203] <= 16'b0000000000001000;
        weights1[1204] <= 16'b1111111111001000;
        weights1[1205] <= 16'b1111111110100110;
        weights1[1206] <= 16'b1111111110101010;
        weights1[1207] <= 16'b1111111110110001;
        weights1[1208] <= 16'b1111111111001010;
        weights1[1209] <= 16'b1111111111110010;
        weights1[1210] <= 16'b0000000000101101;
        weights1[1211] <= 16'b0000000000100010;
        weights1[1212] <= 16'b0000000000001001;
        weights1[1213] <= 16'b0000000000001111;
        weights1[1214] <= 16'b0000000000011101;
        weights1[1215] <= 16'b0000000000011001;
        weights1[1216] <= 16'b0000000000001110;
        weights1[1217] <= 16'b0000000000000000;
        weights1[1218] <= 16'b1111111111110111;
        weights1[1219] <= 16'b0000000000000111;
        weights1[1220] <= 16'b1111111111110110;
        weights1[1221] <= 16'b0000000000001001;
        weights1[1222] <= 16'b0000000000001011;
        weights1[1223] <= 16'b1111111111101001;
        weights1[1224] <= 16'b1111111111111101;
        weights1[1225] <= 16'b1111111111111000;
        weights1[1226] <= 16'b1111111111011100;
        weights1[1227] <= 16'b0000000000001011;
        weights1[1228] <= 16'b0000000000000000;
        weights1[1229] <= 16'b1111111111111011;
        weights1[1230] <= 16'b0000000000010000;
        weights1[1231] <= 16'b0000000000000001;
        weights1[1232] <= 16'b1111111111001010;
        weights1[1233] <= 16'b1111111110111000;
        weights1[1234] <= 16'b1111111110100110;
        weights1[1235] <= 16'b1111111101111101;
        weights1[1236] <= 16'b1111111101001001;
        weights1[1237] <= 16'b1111111101110000;
        weights1[1238] <= 16'b1111111110110001;
        weights1[1239] <= 16'b1111111111010100;
        weights1[1240] <= 16'b0000000000000100;
        weights1[1241] <= 16'b0000000000010010;
        weights1[1242] <= 16'b0000000000000100;
        weights1[1243] <= 16'b0000000001000000;
        weights1[1244] <= 16'b0000000000100110;
        weights1[1245] <= 16'b0000000000100010;
        weights1[1246] <= 16'b0000000000001001;
        weights1[1247] <= 16'b1111111111111111;
        weights1[1248] <= 16'b0000000000000010;
        weights1[1249] <= 16'b0000000000000001;
        weights1[1250] <= 16'b1111111111101100;
        weights1[1251] <= 16'b0000000000000010;
        weights1[1252] <= 16'b1111111111110010;
        weights1[1253] <= 16'b1111111111110100;
        weights1[1254] <= 16'b1111111111111101;
        weights1[1255] <= 16'b1111111111110000;
        weights1[1256] <= 16'b1111111111111011;
        weights1[1257] <= 16'b0000000000001101;
        weights1[1258] <= 16'b0000000000010011;
        weights1[1259] <= 16'b0000000000000101;
        weights1[1260] <= 16'b1111111111010001;
        weights1[1261] <= 16'b1111111110110100;
        weights1[1262] <= 16'b1111111110110111;
        weights1[1263] <= 16'b1111111110000010;
        weights1[1264] <= 16'b1111111101011001;
        weights1[1265] <= 16'b1111111100101010;
        weights1[1266] <= 16'b1111111011101011;
        weights1[1267] <= 16'b1111111100011111;
        weights1[1268] <= 16'b1111111101101101;
        weights1[1269] <= 16'b1111111110111100;
        weights1[1270] <= 16'b1111111111100010;
        weights1[1271] <= 16'b0000000000000100;
        weights1[1272] <= 16'b0000000000010100;
        weights1[1273] <= 16'b0000000000001101;
        weights1[1274] <= 16'b0000000000000101;
        weights1[1275] <= 16'b1111111111110011;
        weights1[1276] <= 16'b1111111111101100;
        weights1[1277] <= 16'b1111111111100000;
        weights1[1278] <= 16'b1111111111111000;
        weights1[1279] <= 16'b1111111111101100;
        weights1[1280] <= 16'b1111111111111000;
        weights1[1281] <= 16'b1111111111110010;
        weights1[1282] <= 16'b1111111111110100;
        weights1[1283] <= 16'b0000000000001001;
        weights1[1284] <= 16'b1111111111111011;
        weights1[1285] <= 16'b0000000000000101;
        weights1[1286] <= 16'b0000000000000010;
        weights1[1287] <= 16'b0000000000001010;
        weights1[1288] <= 16'b1111111111011010;
        weights1[1289] <= 16'b1111111111001011;
        weights1[1290] <= 16'b1111111111001010;
        weights1[1291] <= 16'b1111111110111001;
        weights1[1292] <= 16'b1111111110011011;
        weights1[1293] <= 16'b1111111101101101;
        weights1[1294] <= 16'b1111111101000001;
        weights1[1295] <= 16'b1111111100000110;
        weights1[1296] <= 16'b1111111010111000;
        weights1[1297] <= 16'b1111111010101000;
        weights1[1298] <= 16'b1111111010110000;
        weights1[1299] <= 16'b1111111011101101;
        weights1[1300] <= 16'b1111111101000000;
        weights1[1301] <= 16'b1111111101111010;
        weights1[1302] <= 16'b1111111110010111;
        weights1[1303] <= 16'b1111111111001100;
        weights1[1304] <= 16'b1111111111001011;
        weights1[1305] <= 16'b1111111111100101;
        weights1[1306] <= 16'b1111111111110110;
        weights1[1307] <= 16'b1111111111111001;
        weights1[1308] <= 16'b1111111111111000;
        weights1[1309] <= 16'b1111111111111010;
        weights1[1310] <= 16'b0000000000000010;
        weights1[1311] <= 16'b0000000000010010;
        weights1[1312] <= 16'b1111111111111011;
        weights1[1313] <= 16'b0000000000001011;
        weights1[1314] <= 16'b0000000000000011;
        weights1[1315] <= 16'b0000000000001010;
        weights1[1316] <= 16'b1111111111110110;
        weights1[1317] <= 16'b1111111111101111;
        weights1[1318] <= 16'b1111111111110000;
        weights1[1319] <= 16'b1111111111101111;
        weights1[1320] <= 16'b1111111111011010;
        weights1[1321] <= 16'b1111111111100101;
        weights1[1322] <= 16'b1111111111010101;
        weights1[1323] <= 16'b1111111110101110;
        weights1[1324] <= 16'b1111111101010110;
        weights1[1325] <= 16'b1111111100100110;
        weights1[1326] <= 16'b1111111100011100;
        weights1[1327] <= 16'b1111111101000011;
        weights1[1328] <= 16'b1111111101100010;
        weights1[1329] <= 16'b1111111110101010;
        weights1[1330] <= 16'b1111111110110110;
        weights1[1331] <= 16'b1111111110111010;
        weights1[1332] <= 16'b1111111111110010;
        weights1[1333] <= 16'b1111111111110100;
        weights1[1334] <= 16'b1111111111110111;
        weights1[1335] <= 16'b1111111111111100;
        weights1[1336] <= 16'b0000000000011000;
        weights1[1337] <= 16'b1111111111111000;
        weights1[1338] <= 16'b0000000000001010;
        weights1[1339] <= 16'b1111111111111010;
        weights1[1340] <= 16'b0000000000010110;
        weights1[1341] <= 16'b0000000000001000;
        weights1[1342] <= 16'b0000000000010010;
        weights1[1343] <= 16'b0000000000000110;
        weights1[1344] <= 16'b0000000000000010;
        weights1[1345] <= 16'b0000000000000110;
        weights1[1346] <= 16'b0000000000010000;
        weights1[1347] <= 16'b0000000000001110;
        weights1[1348] <= 16'b0000000000010100;
        weights1[1349] <= 16'b0000000000001110;
        weights1[1350] <= 16'b0000000000011000;
        weights1[1351] <= 16'b0000000000010011;
        weights1[1352] <= 16'b0000000000111110;
        weights1[1353] <= 16'b0000000000111010;
        weights1[1354] <= 16'b0000000000101000;
        weights1[1355] <= 16'b0000000000101001;
        weights1[1356] <= 16'b1111111111111001;
        weights1[1357] <= 16'b1111111111110010;
        weights1[1358] <= 16'b0000000000000101;
        weights1[1359] <= 16'b1111111111111011;
        weights1[1360] <= 16'b1111111111111100;
        weights1[1361] <= 16'b0000000000000101;
        weights1[1362] <= 16'b0000000000001011;
        weights1[1363] <= 16'b0000000000001111;
        weights1[1364] <= 16'b0000000000000011;
        weights1[1365] <= 16'b0000000000001001;
        weights1[1366] <= 16'b0000000000010011;
        weights1[1367] <= 16'b0000000000000001;
        weights1[1368] <= 16'b1111111111111110;
        weights1[1369] <= 16'b0000000000001001;
        weights1[1370] <= 16'b0000000000001111;
        weights1[1371] <= 16'b0000000000001011;
        weights1[1372] <= 16'b0000000000010101;
        weights1[1373] <= 16'b0000000000010011;
        weights1[1374] <= 16'b0000000000011100;
        weights1[1375] <= 16'b0000000000011111;
        weights1[1376] <= 16'b0000000000110010;
        weights1[1377] <= 16'b0000000001000101;
        weights1[1378] <= 16'b0000000001011010;
        weights1[1379] <= 16'b0000000001001111;
        weights1[1380] <= 16'b0000000001101100;
        weights1[1381] <= 16'b0000000001011101;
        weights1[1382] <= 16'b0000000001000011;
        weights1[1383] <= 16'b0000000000111111;
        weights1[1384] <= 16'b0000000000101000;
        weights1[1385] <= 16'b0000000000100101;
        weights1[1386] <= 16'b0000000000000111;
        weights1[1387] <= 16'b0000000000001000;
        weights1[1388] <= 16'b0000000000011010;
        weights1[1389] <= 16'b1111111111110111;
        weights1[1390] <= 16'b1111111111110110;
        weights1[1391] <= 16'b0000000000001101;
        weights1[1392] <= 16'b1111111111111000;
        weights1[1393] <= 16'b0000000000000010;
        weights1[1394] <= 16'b1111111111111000;
        weights1[1395] <= 16'b0000000000001010;
        weights1[1396] <= 16'b0000000000000111;
        weights1[1397] <= 16'b0000000000000011;
        weights1[1398] <= 16'b0000000000000101;
        weights1[1399] <= 16'b1111111111111100;
        weights1[1400] <= 16'b0000000000000111;
        weights1[1401] <= 16'b0000000000000111;
        weights1[1402] <= 16'b0000000000100001;
        weights1[1403] <= 16'b0000000000100001;
        weights1[1404] <= 16'b0000000000101011;
        weights1[1405] <= 16'b0000000000101010;
        weights1[1406] <= 16'b0000000000011010;
        weights1[1407] <= 16'b0000000001000101;
        weights1[1408] <= 16'b0000000000111011;
        weights1[1409] <= 16'b0000000000111000;
        weights1[1410] <= 16'b0000000000100110;
        weights1[1411] <= 16'b0000000000111100;
        weights1[1412] <= 16'b0000000000011011;
        weights1[1413] <= 16'b0000000000001110;
        weights1[1414] <= 16'b0000000000101100;
        weights1[1415] <= 16'b0000000000000101;
        weights1[1416] <= 16'b0000000000000101;
        weights1[1417] <= 16'b1111111111111000;
        weights1[1418] <= 16'b0000000000000110;
        weights1[1419] <= 16'b1111111111111101;
        weights1[1420] <= 16'b1111111111111011;
        weights1[1421] <= 16'b0000000000000000;
        weights1[1422] <= 16'b0000000000001101;
        weights1[1423] <= 16'b1111111111110110;
        weights1[1424] <= 16'b0000000000000100;
        weights1[1425] <= 16'b1111111111110101;
        weights1[1426] <= 16'b0000000000000100;
        weights1[1427] <= 16'b0000000000000010;
        weights1[1428] <= 16'b0000000000001001;
        weights1[1429] <= 16'b0000000000000101;
        weights1[1430] <= 16'b0000000000010001;
        weights1[1431] <= 16'b0000000000100001;
        weights1[1432] <= 16'b0000000000100011;
        weights1[1433] <= 16'b0000000001000001;
        weights1[1434] <= 16'b0000000000101111;
        weights1[1435] <= 16'b0000000000000100;
        weights1[1436] <= 16'b1111111111110111;
        weights1[1437] <= 16'b0000000000100000;
        weights1[1438] <= 16'b0000000000011011;
        weights1[1439] <= 16'b0000000000001000;
        weights1[1440] <= 16'b0000000000001100;
        weights1[1441] <= 16'b0000000000100011;
        weights1[1442] <= 16'b1111111111111011;
        weights1[1443] <= 16'b0000000000010011;
        weights1[1444] <= 16'b0000000000000101;
        weights1[1445] <= 16'b0000000000001011;
        weights1[1446] <= 16'b0000000000000111;
        weights1[1447] <= 16'b0000000000000011;
        weights1[1448] <= 16'b0000000000010010;
        weights1[1449] <= 16'b1111111111111010;
        weights1[1450] <= 16'b0000000000001000;
        weights1[1451] <= 16'b0000000000001110;
        weights1[1452] <= 16'b0000000000001011;
        weights1[1453] <= 16'b1111111111110110;
        weights1[1454] <= 16'b1111111111111011;
        weights1[1455] <= 16'b1111111111111110;
        weights1[1456] <= 16'b0000000000000000;
        weights1[1457] <= 16'b1111111111111100;
        weights1[1458] <= 16'b1111111111110010;
        weights1[1459] <= 16'b0000000000010111;
        weights1[1460] <= 16'b0000000000001011;
        weights1[1461] <= 16'b0000000000010010;
        weights1[1462] <= 16'b0000000000101000;
        weights1[1463] <= 16'b0000000000110110;
        weights1[1464] <= 16'b0000000000010100;
        weights1[1465] <= 16'b0000000000100000;
        weights1[1466] <= 16'b0000000000001100;
        weights1[1467] <= 16'b0000000000100010;
        weights1[1468] <= 16'b0000000000000001;
        weights1[1469] <= 16'b0000000000000011;
        weights1[1470] <= 16'b0000000000011011;
        weights1[1471] <= 16'b1111111111111110;
        weights1[1472] <= 16'b0000000000000000;
        weights1[1473] <= 16'b0000000000001110;
        weights1[1474] <= 16'b1111111111111110;
        weights1[1475] <= 16'b1111111111110110;
        weights1[1476] <= 16'b0000000000000101;
        weights1[1477] <= 16'b1111111111111001;
        weights1[1478] <= 16'b0000000000000001;
        weights1[1479] <= 16'b1111111111110110;
        weights1[1480] <= 16'b1111111111101110;
        weights1[1481] <= 16'b1111111111110111;
        weights1[1482] <= 16'b1111111111111110;
        weights1[1483] <= 16'b1111111111111100;
        weights1[1484] <= 16'b1111111111111100;
        weights1[1485] <= 16'b1111111111111110;
        weights1[1486] <= 16'b1111111111110110;
        weights1[1487] <= 16'b1111111111110001;
        weights1[1488] <= 16'b1111111111111010;
        weights1[1489] <= 16'b1111111111111010;
        weights1[1490] <= 16'b1111111111110010;
        weights1[1491] <= 16'b0000000000010010;
        weights1[1492] <= 16'b0000000000000010;
        weights1[1493] <= 16'b0000000000001111;
        weights1[1494] <= 16'b0000000000000111;
        weights1[1495] <= 16'b0000000000001011;
        weights1[1496] <= 16'b0000000000011000;
        weights1[1497] <= 16'b0000000000010010;
        weights1[1498] <= 16'b1111111111111100;
        weights1[1499] <= 16'b0000000000010100;
        weights1[1500] <= 16'b0000000000000001;
        weights1[1501] <= 16'b0000000000000101;
        weights1[1502] <= 16'b0000000000000011;
        weights1[1503] <= 16'b0000000000001001;
        weights1[1504] <= 16'b1111111111111111;
        weights1[1505] <= 16'b0000000000000001;
        weights1[1506] <= 16'b1111111111111110;
        weights1[1507] <= 16'b0000000000000000;
        weights1[1508] <= 16'b1111111111111100;
        weights1[1509] <= 16'b1111111111110011;
        weights1[1510] <= 16'b1111111111111111;
        weights1[1511] <= 16'b1111111111111100;
        weights1[1512] <= 16'b1111111111111101;
        weights1[1513] <= 16'b1111111111111101;
        weights1[1514] <= 16'b1111111111111100;
        weights1[1515] <= 16'b1111111111101111;
        weights1[1516] <= 16'b1111111111011110;
        weights1[1517] <= 16'b1111111111011101;
        weights1[1518] <= 16'b1111111111010111;
        weights1[1519] <= 16'b1111111111001111;
        weights1[1520] <= 16'b1111111111100000;
        weights1[1521] <= 16'b1111111111110101;
        weights1[1522] <= 16'b1111111111111011;
        weights1[1523] <= 16'b1111111111101001;
        weights1[1524] <= 16'b1111111111100111;
        weights1[1525] <= 16'b0000000000000011;
        weights1[1526] <= 16'b0000000000001011;
        weights1[1527] <= 16'b1111111111101111;
        weights1[1528] <= 16'b0000000000011010;
        weights1[1529] <= 16'b1111111111110100;
        weights1[1530] <= 16'b1111111111111010;
        weights1[1531] <= 16'b0000000000000110;
        weights1[1532] <= 16'b0000000000000111;
        weights1[1533] <= 16'b0000000000000000;
        weights1[1534] <= 16'b1111111111101110;
        weights1[1535] <= 16'b1111111111111011;
        weights1[1536] <= 16'b1111111111111010;
        weights1[1537] <= 16'b1111111111111110;
        weights1[1538] <= 16'b1111111111111100;
        weights1[1539] <= 16'b0000000000000000;
        weights1[1540] <= 16'b0000000000000000;
        weights1[1541] <= 16'b1111111111111111;
        weights1[1542] <= 16'b1111111111111001;
        weights1[1543] <= 16'b1111111111101110;
        weights1[1544] <= 16'b1111111111100101;
        weights1[1545] <= 16'b1111111111100001;
        weights1[1546] <= 16'b1111111111100110;
        weights1[1547] <= 16'b1111111111010010;
        weights1[1548] <= 16'b1111111111010000;
        weights1[1549] <= 16'b1111111111011011;
        weights1[1550] <= 16'b1111111111101111;
        weights1[1551] <= 16'b1111111111101010;
        weights1[1552] <= 16'b1111111111111100;
        weights1[1553] <= 16'b1111111111111000;
        weights1[1554] <= 16'b1111111111100001;
        weights1[1555] <= 16'b1111111111100110;
        weights1[1556] <= 16'b1111111111011111;
        weights1[1557] <= 16'b1111111111100101;
        weights1[1558] <= 16'b1111111111110000;
        weights1[1559] <= 16'b1111111111100010;
        weights1[1560] <= 16'b1111111111110001;
        weights1[1561] <= 16'b1111111111101101;
        weights1[1562] <= 16'b1111111111111000;
        weights1[1563] <= 16'b0000000000000011;
        weights1[1564] <= 16'b1111111111111111;
        weights1[1565] <= 16'b0000000000000001;
        weights1[1566] <= 16'b1111111111111101;
        weights1[1567] <= 16'b0000000000000000;
        weights1[1568] <= 16'b0000000000000000;
        weights1[1569] <= 16'b0000000000000000;
        weights1[1570] <= 16'b0000000000000000;
        weights1[1571] <= 16'b0000000000000000;
        weights1[1572] <= 16'b1111111111111110;
        weights1[1573] <= 16'b1111111111111111;
        weights1[1574] <= 16'b1111111111111000;
        weights1[1575] <= 16'b1111111111110101;
        weights1[1576] <= 16'b1111111111111001;
        weights1[1577] <= 16'b0000000000000110;
        weights1[1578] <= 16'b0000000000000100;
        weights1[1579] <= 16'b0000000000001101;
        weights1[1580] <= 16'b0000000000010000;
        weights1[1581] <= 16'b1111111111110101;
        weights1[1582] <= 16'b1111111111111111;
        weights1[1583] <= 16'b0000000000001100;
        weights1[1584] <= 16'b0000000000000010;
        weights1[1585] <= 16'b0000000000000010;
        weights1[1586] <= 16'b0000000000000010;
        weights1[1587] <= 16'b0000000000001000;
        weights1[1588] <= 16'b0000000000000001;
        weights1[1589] <= 16'b1111111111111101;
        weights1[1590] <= 16'b1111111111111100;
        weights1[1591] <= 16'b1111111111111111;
        weights1[1592] <= 16'b0000000000000000;
        weights1[1593] <= 16'b0000000000000001;
        weights1[1594] <= 16'b0000000000000000;
        weights1[1595] <= 16'b0000000000000000;
        weights1[1596] <= 16'b0000000000000000;
        weights1[1597] <= 16'b0000000000000000;
        weights1[1598] <= 16'b0000000000000000;
        weights1[1599] <= 16'b1111111111111111;
        weights1[1600] <= 16'b1111111111111001;
        weights1[1601] <= 16'b1111111111110101;
        weights1[1602] <= 16'b1111111111110101;
        weights1[1603] <= 16'b1111111111110000;
        weights1[1604] <= 16'b1111111111110110;
        weights1[1605] <= 16'b0000000000000101;
        weights1[1606] <= 16'b0000000000010000;
        weights1[1607] <= 16'b0000000000000111;
        weights1[1608] <= 16'b0000000000000010;
        weights1[1609] <= 16'b1111111111101100;
        weights1[1610] <= 16'b1111111111111001;
        weights1[1611] <= 16'b0000000000001101;
        weights1[1612] <= 16'b0000000000000010;
        weights1[1613] <= 16'b1111111111111101;
        weights1[1614] <= 16'b0000000000000101;
        weights1[1615] <= 16'b0000000000000011;
        weights1[1616] <= 16'b0000000000000011;
        weights1[1617] <= 16'b1111111111111000;
        weights1[1618] <= 16'b1111111111111001;
        weights1[1619] <= 16'b1111111111110111;
        weights1[1620] <= 16'b1111111111111011;
        weights1[1621] <= 16'b1111111111111101;
        weights1[1622] <= 16'b1111111111111110;
        weights1[1623] <= 16'b1111111111111111;
        weights1[1624] <= 16'b0000000000000000;
        weights1[1625] <= 16'b0000000000000000;
        weights1[1626] <= 16'b1111111111111111;
        weights1[1627] <= 16'b1111111111111010;
        weights1[1628] <= 16'b1111111111110100;
        weights1[1629] <= 16'b1111111111101101;
        weights1[1630] <= 16'b1111111111101001;
        weights1[1631] <= 16'b1111111111101010;
        weights1[1632] <= 16'b1111111111110110;
        weights1[1633] <= 16'b0000000000000100;
        weights1[1634] <= 16'b0000000000010111;
        weights1[1635] <= 16'b0000000000010000;
        weights1[1636] <= 16'b1111111111110100;
        weights1[1637] <= 16'b0000000000001100;
        weights1[1638] <= 16'b1111111111101111;
        weights1[1639] <= 16'b0000000000000010;
        weights1[1640] <= 16'b0000000000000011;
        weights1[1641] <= 16'b1111111111111011;
        weights1[1642] <= 16'b0000000000000010;
        weights1[1643] <= 16'b0000000000011101;
        weights1[1644] <= 16'b1111111111111100;
        weights1[1645] <= 16'b1111111111111001;
        weights1[1646] <= 16'b1111111111110111;
        weights1[1647] <= 16'b1111111111110101;
        weights1[1648] <= 16'b1111111111110100;
        weights1[1649] <= 16'b1111111111111101;
        weights1[1650] <= 16'b1111111111111111;
        weights1[1651] <= 16'b0000000000000000;
        weights1[1652] <= 16'b0000000000000000;
        weights1[1653] <= 16'b0000000000000000;
        weights1[1654] <= 16'b1111111111111001;
        weights1[1655] <= 16'b1111111111110100;
        weights1[1656] <= 16'b1111111111110010;
        weights1[1657] <= 16'b1111111111100110;
        weights1[1658] <= 16'b1111111111011100;
        weights1[1659] <= 16'b1111111111011100;
        weights1[1660] <= 16'b1111111111101001;
        weights1[1661] <= 16'b0000000000001010;
        weights1[1662] <= 16'b0000000000001100;
        weights1[1663] <= 16'b0000000000000101;
        weights1[1664] <= 16'b1111111111111011;
        weights1[1665] <= 16'b1111111111101101;
        weights1[1666] <= 16'b1111111111111110;
        weights1[1667] <= 16'b1111111111111100;
        weights1[1668] <= 16'b1111111111111010;
        weights1[1669] <= 16'b0000000000000100;
        weights1[1670] <= 16'b0000000000001110;
        weights1[1671] <= 16'b0000000000000000;
        weights1[1672] <= 16'b0000000000000101;
        weights1[1673] <= 16'b1111111111110011;
        weights1[1674] <= 16'b1111111111110010;
        weights1[1675] <= 16'b1111111111110100;
        weights1[1676] <= 16'b1111111111110101;
        weights1[1677] <= 16'b1111111111111101;
        weights1[1678] <= 16'b1111111111111111;
        weights1[1679] <= 16'b0000000000000000;
        weights1[1680] <= 16'b1111111111111110;
        weights1[1681] <= 16'b1111111111111100;
        weights1[1682] <= 16'b0000000000000000;
        weights1[1683] <= 16'b1111111111110001;
        weights1[1684] <= 16'b1111111111101100;
        weights1[1685] <= 16'b1111111111101000;
        weights1[1686] <= 16'b1111111111011001;
        weights1[1687] <= 16'b1111111111011001;
        weights1[1688] <= 16'b1111111111100101;
        weights1[1689] <= 16'b0000000000000101;
        weights1[1690] <= 16'b0000000000001001;
        weights1[1691] <= 16'b0000000000100111;
        weights1[1692] <= 16'b1111111111110101;
        weights1[1693] <= 16'b0000000000001001;
        weights1[1694] <= 16'b1111111111111100;
        weights1[1695] <= 16'b0000000000001000;
        weights1[1696] <= 16'b1111111111110011;
        weights1[1697] <= 16'b0000000000001010;
        weights1[1698] <= 16'b0000000000001000;
        weights1[1699] <= 16'b1111111111101000;
        weights1[1700] <= 16'b1111111111111101;
        weights1[1701] <= 16'b1111111111101111;
        weights1[1702] <= 16'b1111111111010111;
        weights1[1703] <= 16'b1111111111101111;
        weights1[1704] <= 16'b1111111111110101;
        weights1[1705] <= 16'b1111111111111011;
        weights1[1706] <= 16'b1111111111111111;
        weights1[1707] <= 16'b1111111111111111;
        weights1[1708] <= 16'b0000000000000000;
        weights1[1709] <= 16'b1111111111111100;
        weights1[1710] <= 16'b1111111111111100;
        weights1[1711] <= 16'b1111111111111110;
        weights1[1712] <= 16'b1111111111111101;
        weights1[1713] <= 16'b1111111111110111;
        weights1[1714] <= 16'b1111111111011101;
        weights1[1715] <= 16'b1111111111110010;
        weights1[1716] <= 16'b1111111111100000;
        weights1[1717] <= 16'b1111111111111110;
        weights1[1718] <= 16'b0000000000000101;
        weights1[1719] <= 16'b0000000000000111;
        weights1[1720] <= 16'b1111111111101001;
        weights1[1721] <= 16'b1111111111111101;
        weights1[1722] <= 16'b1111111111011100;
        weights1[1723] <= 16'b1111111111110100;
        weights1[1724] <= 16'b1111111111111001;
        weights1[1725] <= 16'b1111111111010000;
        weights1[1726] <= 16'b1111111111100111;
        weights1[1727] <= 16'b1111111111101011;
        weights1[1728] <= 16'b1111111111101110;
        weights1[1729] <= 16'b1111111111011001;
        weights1[1730] <= 16'b1111111111010000;
        weights1[1731] <= 16'b1111111111011100;
        weights1[1732] <= 16'b1111111111110100;
        weights1[1733] <= 16'b1111111111111011;
        weights1[1734] <= 16'b0000000000000100;
        weights1[1735] <= 16'b0000000000000010;
        weights1[1736] <= 16'b0000000000000011;
        weights1[1737] <= 16'b1111111111111110;
        weights1[1738] <= 16'b1111111111111110;
        weights1[1739] <= 16'b1111111111111100;
        weights1[1740] <= 16'b1111111111110010;
        weights1[1741] <= 16'b1111111111101111;
        weights1[1742] <= 16'b1111111111101000;
        weights1[1743] <= 16'b1111111111101000;
        weights1[1744] <= 16'b1111111111011111;
        weights1[1745] <= 16'b1111111111010001;
        weights1[1746] <= 16'b1111111111110010;
        weights1[1747] <= 16'b0000000000010001;
        weights1[1748] <= 16'b0000000000000101;
        weights1[1749] <= 16'b1111111111111110;
        weights1[1750] <= 16'b1111111111101001;
        weights1[1751] <= 16'b1111111111110010;
        weights1[1752] <= 16'b1111111111111000;
        weights1[1753] <= 16'b1111111111110001;
        weights1[1754] <= 16'b1111111111110000;
        weights1[1755] <= 16'b1111111111001100;
        weights1[1756] <= 16'b1111111111011111;
        weights1[1757] <= 16'b1111111111000111;
        weights1[1758] <= 16'b1111111111011100;
        weights1[1759] <= 16'b1111111111101011;
        weights1[1760] <= 16'b1111111111110001;
        weights1[1761] <= 16'b1111111111110001;
        weights1[1762] <= 16'b0000000000000001;
        weights1[1763] <= 16'b0000000000000001;
        weights1[1764] <= 16'b0000000000000100;
        weights1[1765] <= 16'b0000000000001001;
        weights1[1766] <= 16'b0000000000000101;
        weights1[1767] <= 16'b0000000000001000;
        weights1[1768] <= 16'b0000000000000001;
        weights1[1769] <= 16'b0000000000000000;
        weights1[1770] <= 16'b0000000000000000;
        weights1[1771] <= 16'b1111111111101000;
        weights1[1772] <= 16'b1111111111101010;
        weights1[1773] <= 16'b1111111111010110;
        weights1[1774] <= 16'b1111111111101000;
        weights1[1775] <= 16'b0000000000010010;
        weights1[1776] <= 16'b0000000000010011;
        weights1[1777] <= 16'b1111111111111110;
        weights1[1778] <= 16'b1111111111111110;
        weights1[1779] <= 16'b1111111111101011;
        weights1[1780] <= 16'b1111111111110101;
        weights1[1781] <= 16'b0000000000001100;
        weights1[1782] <= 16'b1111111111010110;
        weights1[1783] <= 16'b1111111111101011;
        weights1[1784] <= 16'b1111111111001011;
        weights1[1785] <= 16'b1111111111000110;
        weights1[1786] <= 16'b1111111111100110;
        weights1[1787] <= 16'b1111111111101110;
        weights1[1788] <= 16'b1111111111101000;
        weights1[1789] <= 16'b1111111111110010;
        weights1[1790] <= 16'b0000000000000001;
        weights1[1791] <= 16'b0000000000000010;
        weights1[1792] <= 16'b0000000000001011;
        weights1[1793] <= 16'b0000000000001001;
        weights1[1794] <= 16'b0000000000001000;
        weights1[1795] <= 16'b0000000000001101;
        weights1[1796] <= 16'b0000000000001000;
        weights1[1797] <= 16'b0000000000000101;
        weights1[1798] <= 16'b0000000000010001;
        weights1[1799] <= 16'b1111111111111010;
        weights1[1800] <= 16'b1111111111011110;
        weights1[1801] <= 16'b1111111111101001;
        weights1[1802] <= 16'b1111111111100111;
        weights1[1803] <= 16'b1111111111110110;
        weights1[1804] <= 16'b1111111111110111;
        weights1[1805] <= 16'b0000000000010000;
        weights1[1806] <= 16'b0000000000011010;
        weights1[1807] <= 16'b0000000000001101;
        weights1[1808] <= 16'b1111111111110110;
        weights1[1809] <= 16'b1111111111101001;
        weights1[1810] <= 16'b1111111110111000;
        weights1[1811] <= 16'b1111111111011111;
        weights1[1812] <= 16'b1111111110111011;
        weights1[1813] <= 16'b1111111110111010;
        weights1[1814] <= 16'b1111111111011111;
        weights1[1815] <= 16'b1111111111100010;
        weights1[1816] <= 16'b1111111111100111;
        weights1[1817] <= 16'b1111111111101101;
        weights1[1818] <= 16'b0000000000000001;
        weights1[1819] <= 16'b0000000000000101;
        weights1[1820] <= 16'b0000000000001001;
        weights1[1821] <= 16'b0000000000010000;
        weights1[1822] <= 16'b0000000000001101;
        weights1[1823] <= 16'b0000000000000111;
        weights1[1824] <= 16'b1111111111101110;
        weights1[1825] <= 16'b1111111111111111;
        weights1[1826] <= 16'b0000000000001010;
        weights1[1827] <= 16'b0000000000000100;
        weights1[1828] <= 16'b1111111111110001;
        weights1[1829] <= 16'b1111111111010101;
        weights1[1830] <= 16'b1111111111101001;
        weights1[1831] <= 16'b1111111111110100;
        weights1[1832] <= 16'b1111111111110000;
        weights1[1833] <= 16'b0000000000000001;
        weights1[1834] <= 16'b0000000000101100;
        weights1[1835] <= 16'b0000000000010111;
        weights1[1836] <= 16'b1111111111111110;
        weights1[1837] <= 16'b1111111111100100;
        weights1[1838] <= 16'b1111111111011010;
        weights1[1839] <= 16'b1111111111000011;
        weights1[1840] <= 16'b1111111110101110;
        weights1[1841] <= 16'b1111111111001100;
        weights1[1842] <= 16'b1111111111011001;
        weights1[1843] <= 16'b1111111111100011;
        weights1[1844] <= 16'b1111111111101000;
        weights1[1845] <= 16'b1111111111110011;
        weights1[1846] <= 16'b1111111111111101;
        weights1[1847] <= 16'b1111111111111111;
        weights1[1848] <= 16'b0000000000000111;
        weights1[1849] <= 16'b0000000000000111;
        weights1[1850] <= 16'b0000000000001001;
        weights1[1851] <= 16'b0000000000000100;
        weights1[1852] <= 16'b1111111111111101;
        weights1[1853] <= 16'b1111111111110010;
        weights1[1854] <= 16'b1111111111110010;
        weights1[1855] <= 16'b1111111111110111;
        weights1[1856] <= 16'b0000000000001001;
        weights1[1857] <= 16'b1111111111010110;
        weights1[1858] <= 16'b1111111111100000;
        weights1[1859] <= 16'b1111111111100101;
        weights1[1860] <= 16'b0000000000000000;
        weights1[1861] <= 16'b0000000000010101;
        weights1[1862] <= 16'b0000000000100101;
        weights1[1863] <= 16'b0000000001010010;
        weights1[1864] <= 16'b0000000000000111;
        weights1[1865] <= 16'b1111111111101111;
        weights1[1866] <= 16'b1111111111001001;
        weights1[1867] <= 16'b1111111110010110;
        weights1[1868] <= 16'b1111111110111011;
        weights1[1869] <= 16'b1111111111010001;
        weights1[1870] <= 16'b1111111111100100;
        weights1[1871] <= 16'b1111111111100001;
        weights1[1872] <= 16'b1111111111110100;
        weights1[1873] <= 16'b1111111111110110;
        weights1[1874] <= 16'b1111111111111000;
        weights1[1875] <= 16'b1111111111111111;
        weights1[1876] <= 16'b0000000000001100;
        weights1[1877] <= 16'b0000000000000010;
        weights1[1878] <= 16'b0000000000001001;
        weights1[1879] <= 16'b1111111111110110;
        weights1[1880] <= 16'b0000000000000011;
        weights1[1881] <= 16'b0000000000001111;
        weights1[1882] <= 16'b1111111111110011;
        weights1[1883] <= 16'b1111111111101111;
        weights1[1884] <= 16'b0000000000010010;
        weights1[1885] <= 16'b1111111111100000;
        weights1[1886] <= 16'b1111111111001111;
        weights1[1887] <= 16'b1111111111010000;
        weights1[1888] <= 16'b1111111111100110;
        weights1[1889] <= 16'b0000000000010011;
        weights1[1890] <= 16'b0000000000111010;
        weights1[1891] <= 16'b0000000000011010;
        weights1[1892] <= 16'b0000000000010010;
        weights1[1893] <= 16'b0000000000000101;
        weights1[1894] <= 16'b1111111110011001;
        weights1[1895] <= 16'b1111111110101111;
        weights1[1896] <= 16'b1111111110111110;
        weights1[1897] <= 16'b1111111111010100;
        weights1[1898] <= 16'b1111111111011011;
        weights1[1899] <= 16'b1111111111101010;
        weights1[1900] <= 16'b1111111111101101;
        weights1[1901] <= 16'b1111111111110001;
        weights1[1902] <= 16'b1111111111110101;
        weights1[1903] <= 16'b1111111111111100;
        weights1[1904] <= 16'b0000000000001001;
        weights1[1905] <= 16'b0000000000000110;
        weights1[1906] <= 16'b0000000000000110;
        weights1[1907] <= 16'b0000000000001010;
        weights1[1908] <= 16'b0000000000001101;
        weights1[1909] <= 16'b0000000000011000;
        weights1[1910] <= 16'b1111111111111110;
        weights1[1911] <= 16'b1111111111100010;
        weights1[1912] <= 16'b1111111111101110;
        weights1[1913] <= 16'b1111111111110110;
        weights1[1914] <= 16'b1111111111001010;
        weights1[1915] <= 16'b1111111111010110;
        weights1[1916] <= 16'b0000000000011000;
        weights1[1917] <= 16'b0000000000011010;
        weights1[1918] <= 16'b0000000000101110;
        weights1[1919] <= 16'b0000000000010000;
        weights1[1920] <= 16'b0000000000011000;
        weights1[1921] <= 16'b0000000000000001;
        weights1[1922] <= 16'b1111111110111110;
        weights1[1923] <= 16'b1111111110011001;
        weights1[1924] <= 16'b1111111110110111;
        weights1[1925] <= 16'b1111111111011010;
        weights1[1926] <= 16'b1111111111011101;
        weights1[1927] <= 16'b1111111111110001;
        weights1[1928] <= 16'b1111111111100100;
        weights1[1929] <= 16'b1111111111101111;
        weights1[1930] <= 16'b0000000000000000;
        weights1[1931] <= 16'b1111111111111111;
        weights1[1932] <= 16'b1111111111111111;
        weights1[1933] <= 16'b0000000000000100;
        weights1[1934] <= 16'b0000000000000100;
        weights1[1935] <= 16'b1111111111110110;
        weights1[1936] <= 16'b0000000000000000;
        weights1[1937] <= 16'b1111111111111110;
        weights1[1938] <= 16'b1111111111101110;
        weights1[1939] <= 16'b1111111111100101;
        weights1[1940] <= 16'b1111111111011111;
        weights1[1941] <= 16'b1111111111000000;
        weights1[1942] <= 16'b1111111110101010;
        weights1[1943] <= 16'b1111111111001110;
        weights1[1944] <= 16'b0000000000100011;
        weights1[1945] <= 16'b1111111111111000;
        weights1[1946] <= 16'b0000000000101010;
        weights1[1947] <= 16'b0000000000011010;
        weights1[1948] <= 16'b0000000000001101;
        weights1[1949] <= 16'b1111111111110000;
        weights1[1950] <= 16'b1111111110111001;
        weights1[1951] <= 16'b1111111110110100;
        weights1[1952] <= 16'b1111111110111111;
        weights1[1953] <= 16'b1111111111001111;
        weights1[1954] <= 16'b1111111111011110;
        weights1[1955] <= 16'b1111111111101011;
        weights1[1956] <= 16'b1111111111101011;
        weights1[1957] <= 16'b1111111111110011;
        weights1[1958] <= 16'b1111111111111110;
        weights1[1959] <= 16'b0000000000000001;
        weights1[1960] <= 16'b1111111111111010;
        weights1[1961] <= 16'b1111111111111000;
        weights1[1962] <= 16'b1111111111111101;
        weights1[1963] <= 16'b1111111111111010;
        weights1[1964] <= 16'b0000000000000101;
        weights1[1965] <= 16'b1111111111110110;
        weights1[1966] <= 16'b1111111111110010;
        weights1[1967] <= 16'b1111111111010100;
        weights1[1968] <= 16'b1111111110110110;
        weights1[1969] <= 16'b1111111110101111;
        weights1[1970] <= 16'b1111111111001101;
        weights1[1971] <= 16'b1111111111011000;
        weights1[1972] <= 16'b1111111111110101;
        weights1[1973] <= 16'b1111111111111111;
        weights1[1974] <= 16'b0000000000011110;
        weights1[1975] <= 16'b0000000000010100;
        weights1[1976] <= 16'b0000000000010110;
        weights1[1977] <= 16'b1111111111100110;
        weights1[1978] <= 16'b1111111111001111;
        weights1[1979] <= 16'b1111111110111101;
        weights1[1980] <= 16'b1111111110111001;
        weights1[1981] <= 16'b1111111111001010;
        weights1[1982] <= 16'b1111111111011011;
        weights1[1983] <= 16'b1111111111011011;
        weights1[1984] <= 16'b1111111111101101;
        weights1[1985] <= 16'b1111111111110111;
        weights1[1986] <= 16'b0000000000000110;
        weights1[1987] <= 16'b1111111111110111;
        weights1[1988] <= 16'b1111111111111101;
        weights1[1989] <= 16'b0000000000000001;
        weights1[1990] <= 16'b1111111111111100;
        weights1[1991] <= 16'b1111111111110110;
        weights1[1992] <= 16'b1111111111110111;
        weights1[1993] <= 16'b1111111111101101;
        weights1[1994] <= 16'b1111111111011100;
        weights1[1995] <= 16'b1111111111000110;
        weights1[1996] <= 16'b1111111110101111;
        weights1[1997] <= 16'b1111111111001000;
        weights1[1998] <= 16'b1111111110101100;
        weights1[1999] <= 16'b1111111111101100;
        weights1[2000] <= 16'b1111111111110101;
        weights1[2001] <= 16'b0000000000100010;
        weights1[2002] <= 16'b0000000000001101;
        weights1[2003] <= 16'b0000000000001001;
        weights1[2004] <= 16'b1111111111101001;
        weights1[2005] <= 16'b1111111111010110;
        weights1[2006] <= 16'b1111111111001011;
        weights1[2007] <= 16'b1111111110010100;
        weights1[2008] <= 16'b1111111110100101;
        weights1[2009] <= 16'b1111111111001011;
        weights1[2010] <= 16'b1111111111100010;
        weights1[2011] <= 16'b1111111111100011;
        weights1[2012] <= 16'b1111111111110011;
        weights1[2013] <= 16'b0000000000000010;
        weights1[2014] <= 16'b1111111111111001;
        weights1[2015] <= 16'b1111111111111000;
        weights1[2016] <= 16'b1111111111111010;
        weights1[2017] <= 16'b1111111111111000;
        weights1[2018] <= 16'b1111111111111001;
        weights1[2019] <= 16'b1111111111110001;
        weights1[2020] <= 16'b1111111111100000;
        weights1[2021] <= 16'b1111111111010100;
        weights1[2022] <= 16'b1111111111000010;
        weights1[2023] <= 16'b1111111111000101;
        weights1[2024] <= 16'b1111111111000100;
        weights1[2025] <= 16'b1111111111101100;
        weights1[2026] <= 16'b1111111111011011;
        weights1[2027] <= 16'b1111111111110100;
        weights1[2028] <= 16'b0000000000000110;
        weights1[2029] <= 16'b1111111111111000;
        weights1[2030] <= 16'b0000000000010011;
        weights1[2031] <= 16'b1111111111110001;
        weights1[2032] <= 16'b1111111111110011;
        weights1[2033] <= 16'b1111111111001001;
        weights1[2034] <= 16'b1111111111101100;
        weights1[2035] <= 16'b1111111110110011;
        weights1[2036] <= 16'b1111111110110010;
        weights1[2037] <= 16'b1111111111011001;
        weights1[2038] <= 16'b1111111111100000;
        weights1[2039] <= 16'b1111111111101110;
        weights1[2040] <= 16'b1111111111110100;
        weights1[2041] <= 16'b1111111111111001;
        weights1[2042] <= 16'b1111111111111111;
        weights1[2043] <= 16'b0000000000000001;
        weights1[2044] <= 16'b1111111111111101;
        weights1[2045] <= 16'b1111111111111011;
        weights1[2046] <= 16'b1111111111101111;
        weights1[2047] <= 16'b1111111111011001;
        weights1[2048] <= 16'b1111111111010101;
        weights1[2049] <= 16'b1111111111000111;
        weights1[2050] <= 16'b1111111111100010;
        weights1[2051] <= 16'b1111111111011100;
        weights1[2052] <= 16'b1111111111110011;
        weights1[2053] <= 16'b1111111111101100;
        weights1[2054] <= 16'b1111111111110110;
        weights1[2055] <= 16'b0000000000000101;
        weights1[2056] <= 16'b1111111111111000;
        weights1[2057] <= 16'b0000000000011101;
        weights1[2058] <= 16'b0000000000011001;
        weights1[2059] <= 16'b1111111111101011;
        weights1[2060] <= 16'b1111111111110110;
        weights1[2061] <= 16'b1111111111011010;
        weights1[2062] <= 16'b1111111110111111;
        weights1[2063] <= 16'b1111111110110011;
        weights1[2064] <= 16'b1111111111100011;
        weights1[2065] <= 16'b1111111111011111;
        weights1[2066] <= 16'b1111111111101101;
        weights1[2067] <= 16'b0000000000000001;
        weights1[2068] <= 16'b0000000000000001;
        weights1[2069] <= 16'b1111111111110000;
        weights1[2070] <= 16'b1111111111111101;
        weights1[2071] <= 16'b1111111111111011;
        weights1[2072] <= 16'b0000000000000001;
        weights1[2073] <= 16'b1111111111110010;
        weights1[2074] <= 16'b1111111111101001;
        weights1[2075] <= 16'b1111111111010010;
        weights1[2076] <= 16'b1111111111011010;
        weights1[2077] <= 16'b1111111111011111;
        weights1[2078] <= 16'b1111111111011111;
        weights1[2079] <= 16'b0000000000000010;
        weights1[2080] <= 16'b1111111111111010;
        weights1[2081] <= 16'b0000000000001111;
        weights1[2082] <= 16'b1111111111110000;
        weights1[2083] <= 16'b1111111111101100;
        weights1[2084] <= 16'b1111111111100110;
        weights1[2085] <= 16'b0000000000010100;
        weights1[2086] <= 16'b0000000000010100;
        weights1[2087] <= 16'b0000000000010010;
        weights1[2088] <= 16'b1111111111100000;
        weights1[2089] <= 16'b0000000000000010;
        weights1[2090] <= 16'b0000000000000011;
        weights1[2091] <= 16'b0000000000000001;
        weights1[2092] <= 16'b0000000000100100;
        weights1[2093] <= 16'b1111111111111010;
        weights1[2094] <= 16'b0000000000000101;
        weights1[2095] <= 16'b0000000000100011;
        weights1[2096] <= 16'b0000000000010110;
        weights1[2097] <= 16'b0000000000000001;
        weights1[2098] <= 16'b0000000000000001;
        weights1[2099] <= 16'b0000000000000110;
        weights1[2100] <= 16'b1111111111111100;
        weights1[2101] <= 16'b1111111111110100;
        weights1[2102] <= 16'b1111111111110000;
        weights1[2103] <= 16'b1111111111011000;
        weights1[2104] <= 16'b1111111111100100;
        weights1[2105] <= 16'b1111111111101011;
        weights1[2106] <= 16'b1111111111111101;
        weights1[2107] <= 16'b1111111111110111;
        weights1[2108] <= 16'b1111111111111100;
        weights1[2109] <= 16'b0000000000011100;
        weights1[2110] <= 16'b0000000000001110;
        weights1[2111] <= 16'b1111111111111101;
        weights1[2112] <= 16'b0000000000010000;
        weights1[2113] <= 16'b0000000000011101;
        weights1[2114] <= 16'b0000000000011101;
        weights1[2115] <= 16'b0000000000000111;
        weights1[2116] <= 16'b0000000000011011;
        weights1[2117] <= 16'b1111111111110111;
        weights1[2118] <= 16'b0000000000011101;
        weights1[2119] <= 16'b0000000000010101;
        weights1[2120] <= 16'b0000000000110000;
        weights1[2121] <= 16'b0000000000001001;
        weights1[2122] <= 16'b0000000000000001;
        weights1[2123] <= 16'b0000000000000001;
        weights1[2124] <= 16'b0000000000010001;
        weights1[2125] <= 16'b0000000000010111;
        weights1[2126] <= 16'b0000000000000111;
        weights1[2127] <= 16'b0000000000000110;
        weights1[2128] <= 16'b1111111111111001;
        weights1[2129] <= 16'b1111111111111000;
        weights1[2130] <= 16'b1111111111101100;
        weights1[2131] <= 16'b1111111111100010;
        weights1[2132] <= 16'b1111111111100000;
        weights1[2133] <= 16'b1111111111011010;
        weights1[2134] <= 16'b0000000000001001;
        weights1[2135] <= 16'b0000000000001101;
        weights1[2136] <= 16'b0000000000011111;
        weights1[2137] <= 16'b0000000000011001;
        weights1[2138] <= 16'b0000000000000100;
        weights1[2139] <= 16'b0000000000101001;
        weights1[2140] <= 16'b0000000000011101;
        weights1[2141] <= 16'b0000000000000011;
        weights1[2142] <= 16'b0000000000011110;
        weights1[2143] <= 16'b0000000000011100;
        weights1[2144] <= 16'b0000000000000110;
        weights1[2145] <= 16'b0000000000100100;
        weights1[2146] <= 16'b0000000001000010;
        weights1[2147] <= 16'b0000000000101010;
        weights1[2148] <= 16'b0000000000011101;
        weights1[2149] <= 16'b0000000000010101;
        weights1[2150] <= 16'b0000000000010000;
        weights1[2151] <= 16'b0000000000001110;
        weights1[2152] <= 16'b0000000000010110;
        weights1[2153] <= 16'b0000000000000110;
        weights1[2154] <= 16'b0000000000000111;
        weights1[2155] <= 16'b0000000000000010;
        weights1[2156] <= 16'b1111111111111000;
        weights1[2157] <= 16'b1111111111110001;
        weights1[2158] <= 16'b1111111111110001;
        weights1[2159] <= 16'b1111111111101001;
        weights1[2160] <= 16'b1111111111101011;
        weights1[2161] <= 16'b1111111111111001;
        weights1[2162] <= 16'b1111111111111100;
        weights1[2163] <= 16'b0000000000001100;
        weights1[2164] <= 16'b0000000000001011;
        weights1[2165] <= 16'b0000000000001111;
        weights1[2166] <= 16'b0000000000011000;
        weights1[2167] <= 16'b0000000000001011;
        weights1[2168] <= 16'b1111111111100110;
        weights1[2169] <= 16'b0000000000001000;
        weights1[2170] <= 16'b1111111111111111;
        weights1[2171] <= 16'b0000000000010111;
        weights1[2172] <= 16'b0000000000001101;
        weights1[2173] <= 16'b0000000000011101;
        weights1[2174] <= 16'b0000000000101001;
        weights1[2175] <= 16'b0000000000011001;
        weights1[2176] <= 16'b0000000000100001;
        weights1[2177] <= 16'b0000000000001001;
        weights1[2178] <= 16'b0000000000000101;
        weights1[2179] <= 16'b0000000000001111;
        weights1[2180] <= 16'b0000000000001000;
        weights1[2181] <= 16'b0000000000001000;
        weights1[2182] <= 16'b0000000000000101;
        weights1[2183] <= 16'b0000000000000100;
        weights1[2184] <= 16'b1111111111111100;
        weights1[2185] <= 16'b0000000000000000;
        weights1[2186] <= 16'b1111111111111100;
        weights1[2187] <= 16'b1111111111111010;
        weights1[2188] <= 16'b1111111111111111;
        weights1[2189] <= 16'b1111111111111111;
        weights1[2190] <= 16'b1111111111111001;
        weights1[2191] <= 16'b0000000000000111;
        weights1[2192] <= 16'b0000000000101001;
        weights1[2193] <= 16'b0000000000011001;
        weights1[2194] <= 16'b0000000000011000;
        weights1[2195] <= 16'b1111111111101000;
        weights1[2196] <= 16'b1111111111110000;
        weights1[2197] <= 16'b1111111111001101;
        weights1[2198] <= 16'b1111111111111101;
        weights1[2199] <= 16'b1111111111101110;
        weights1[2200] <= 16'b0000000000001011;
        weights1[2201] <= 16'b0000000000000111;
        weights1[2202] <= 16'b0000000000110000;
        weights1[2203] <= 16'b0000000000100011;
        weights1[2204] <= 16'b0000000000011110;
        weights1[2205] <= 16'b0000000000100001;
        weights1[2206] <= 16'b0000000000010101;
        weights1[2207] <= 16'b0000000000000010;
        weights1[2208] <= 16'b0000000000000110;
        weights1[2209] <= 16'b0000000000001001;
        weights1[2210] <= 16'b0000000000000101;
        weights1[2211] <= 16'b0000000000000011;
        weights1[2212] <= 16'b1111111111111110;
        weights1[2213] <= 16'b0000000000000111;
        weights1[2214] <= 16'b0000000000001000;
        weights1[2215] <= 16'b0000000000000110;
        weights1[2216] <= 16'b0000000000010101;
        weights1[2217] <= 16'b0000000000000101;
        weights1[2218] <= 16'b0000000000000101;
        weights1[2219] <= 16'b0000000000011101;
        weights1[2220] <= 16'b0000000000011110;
        weights1[2221] <= 16'b0000000000000000;
        weights1[2222] <= 16'b0000000000000010;
        weights1[2223] <= 16'b0000000000011110;
        weights1[2224] <= 16'b0000000000001010;
        weights1[2225] <= 16'b1111111111100011;
        weights1[2226] <= 16'b1111111111110101;
        weights1[2227] <= 16'b1111111111111110;
        weights1[2228] <= 16'b1111111111101110;
        weights1[2229] <= 16'b0000000000010010;
        weights1[2230] <= 16'b1111111111110111;
        weights1[2231] <= 16'b0000000000001000;
        weights1[2232] <= 16'b0000000000001110;
        weights1[2233] <= 16'b0000000000000111;
        weights1[2234] <= 16'b0000000000001111;
        weights1[2235] <= 16'b0000000000000101;
        weights1[2236] <= 16'b0000000000000111;
        weights1[2237] <= 16'b0000000000000101;
        weights1[2238] <= 16'b0000000000001000;
        weights1[2239] <= 16'b0000000000000100;
        weights1[2240] <= 16'b0000000000000000;
        weights1[2241] <= 16'b0000000000000001;
        weights1[2242] <= 16'b0000000000000110;
        weights1[2243] <= 16'b0000000000000101;
        weights1[2244] <= 16'b0000000000010010;
        weights1[2245] <= 16'b1111111111111111;
        weights1[2246] <= 16'b0000000000001111;
        weights1[2247] <= 16'b0000000000010001;
        weights1[2248] <= 16'b0000000000010010;
        weights1[2249] <= 16'b0000000000000111;
        weights1[2250] <= 16'b0000000000001110;
        weights1[2251] <= 16'b0000000000000011;
        weights1[2252] <= 16'b1111111111100111;
        weights1[2253] <= 16'b1111111111101000;
        weights1[2254] <= 16'b1111111111011001;
        weights1[2255] <= 16'b1111111111111101;
        weights1[2256] <= 16'b1111111111000100;
        weights1[2257] <= 16'b1111111111101101;
        weights1[2258] <= 16'b1111111111100011;
        weights1[2259] <= 16'b1111111111110101;
        weights1[2260] <= 16'b1111111111111100;
        weights1[2261] <= 16'b0000000000001000;
        weights1[2262] <= 16'b0000000000000110;
        weights1[2263] <= 16'b0000000000000100;
        weights1[2264] <= 16'b0000000000000100;
        weights1[2265] <= 16'b0000000000000001;
        weights1[2266] <= 16'b0000000000000011;
        weights1[2267] <= 16'b1111111111111111;
        weights1[2268] <= 16'b0000000000000100;
        weights1[2269] <= 16'b0000000000000101;
        weights1[2270] <= 16'b0000000000000100;
        weights1[2271] <= 16'b0000000000000010;
        weights1[2272] <= 16'b0000000000010111;
        weights1[2273] <= 16'b0000000000010001;
        weights1[2274] <= 16'b0000000000011100;
        weights1[2275] <= 16'b0000000000000111;
        weights1[2276] <= 16'b0000000000010001;
        weights1[2277] <= 16'b1111111111111011;
        weights1[2278] <= 16'b1111111111111001;
        weights1[2279] <= 16'b1111111111111100;
        weights1[2280] <= 16'b1111111111110101;
        weights1[2281] <= 16'b1111111111101111;
        weights1[2282] <= 16'b1111111111111000;
        weights1[2283] <= 16'b1111111111100001;
        weights1[2284] <= 16'b1111111111111110;
        weights1[2285] <= 16'b0000000000000011;
        weights1[2286] <= 16'b1111111111110110;
        weights1[2287] <= 16'b1111111111111001;
        weights1[2288] <= 16'b1111111111111000;
        weights1[2289] <= 16'b1111111111111110;
        weights1[2290] <= 16'b1111111111111101;
        weights1[2291] <= 16'b1111111111111100;
        weights1[2292] <= 16'b0000000000000010;
        weights1[2293] <= 16'b1111111111111111;
        weights1[2294] <= 16'b1111111111111111;
        weights1[2295] <= 16'b1111111111111111;
        weights1[2296] <= 16'b0000000000000100;
        weights1[2297] <= 16'b0000000000000110;
        weights1[2298] <= 16'b0000000000000011;
        weights1[2299] <= 16'b0000000000000000;
        weights1[2300] <= 16'b0000000000001010;
        weights1[2301] <= 16'b0000000000000111;
        weights1[2302] <= 16'b0000000000000010;
        weights1[2303] <= 16'b0000000000001110;
        weights1[2304] <= 16'b1111111111111100;
        weights1[2305] <= 16'b0000000000000001;
        weights1[2306] <= 16'b0000000000000010;
        weights1[2307] <= 16'b1111111111111110;
        weights1[2308] <= 16'b0000000000001110;
        weights1[2309] <= 16'b1111111111111011;
        weights1[2310] <= 16'b1111111111110100;
        weights1[2311] <= 16'b1111111111110010;
        weights1[2312] <= 16'b0000000000000010;
        weights1[2313] <= 16'b0000000000000001;
        weights1[2314] <= 16'b1111111111101100;
        weights1[2315] <= 16'b1111111111101000;
        weights1[2316] <= 16'b1111111111101110;
        weights1[2317] <= 16'b1111111111111000;
        weights1[2318] <= 16'b1111111111111111;
        weights1[2319] <= 16'b0000000000000000;
        weights1[2320] <= 16'b1111111111111110;
        weights1[2321] <= 16'b1111111111111110;
        weights1[2322] <= 16'b0000000000000000;
        weights1[2323] <= 16'b0000000000000000;
        weights1[2324] <= 16'b1111111111111111;
        weights1[2325] <= 16'b0000000000000001;
        weights1[2326] <= 16'b0000000000000001;
        weights1[2327] <= 16'b0000000000000001;
        weights1[2328] <= 16'b0000000000000111;
        weights1[2329] <= 16'b0000000000001101;
        weights1[2330] <= 16'b0000000000000100;
        weights1[2331] <= 16'b0000000000000100;
        weights1[2332] <= 16'b0000000000001100;
        weights1[2333] <= 16'b0000000000000000;
        weights1[2334] <= 16'b1111111111111000;
        weights1[2335] <= 16'b1111111111101001;
        weights1[2336] <= 16'b1111111111110001;
        weights1[2337] <= 16'b1111111111101111;
        weights1[2338] <= 16'b1111111111101010;
        weights1[2339] <= 16'b1111111111101010;
        weights1[2340] <= 16'b1111111111101101;
        weights1[2341] <= 16'b1111111111101011;
        weights1[2342] <= 16'b1111111111101010;
        weights1[2343] <= 16'b1111111111101110;
        weights1[2344] <= 16'b1111111111101001;
        weights1[2345] <= 16'b1111111111111011;
        weights1[2346] <= 16'b1111111111110111;
        weights1[2347] <= 16'b1111111111110110;
        weights1[2348] <= 16'b1111111111111111;
        weights1[2349] <= 16'b1111111111111101;
        weights1[2350] <= 16'b0000000000000000;
        weights1[2351] <= 16'b0000000000000000;
        weights1[2352] <= 16'b1111111111111111;
        weights1[2353] <= 16'b1111111111111111;
        weights1[2354] <= 16'b1111111111111111;
        weights1[2355] <= 16'b1111111111111111;
        weights1[2356] <= 16'b1111111111111111;
        weights1[2357] <= 16'b0000000000000000;
        weights1[2358] <= 16'b1111111111111010;
        weights1[2359] <= 16'b1111111111111110;
        weights1[2360] <= 16'b1111111111111111;
        weights1[2361] <= 16'b1111111111110100;
        weights1[2362] <= 16'b1111111111101011;
        weights1[2363] <= 16'b1111111111100110;
        weights1[2364] <= 16'b1111111111100001;
        weights1[2365] <= 16'b1111111111100010;
        weights1[2366] <= 16'b1111111111011111;
        weights1[2367] <= 16'b1111111111101011;
        weights1[2368] <= 16'b0000000000001101;
        weights1[2369] <= 16'b0000000000010101;
        weights1[2370] <= 16'b0000000000100110;
        weights1[2371] <= 16'b0000000000010100;
        weights1[2372] <= 16'b0000000000010011;
        weights1[2373] <= 16'b0000000000000110;
        weights1[2374] <= 16'b0000000000000011;
        weights1[2375] <= 16'b1111111111111101;
        weights1[2376] <= 16'b1111111111111010;
        weights1[2377] <= 16'b1111111111111100;
        weights1[2378] <= 16'b1111111111111111;
        weights1[2379] <= 16'b0000000000000000;
        weights1[2380] <= 16'b1111111111111111;
        weights1[2381] <= 16'b0000000000000000;
        weights1[2382] <= 16'b0000000000000000;
        weights1[2383] <= 16'b1111111111111111;
        weights1[2384] <= 16'b1111111111111011;
        weights1[2385] <= 16'b1111111111111011;
        weights1[2386] <= 16'b1111111111111111;
        weights1[2387] <= 16'b0000000000000011;
        weights1[2388] <= 16'b0000000000000110;
        weights1[2389] <= 16'b1111111111101110;
        weights1[2390] <= 16'b1111111111101110;
        weights1[2391] <= 16'b1111111111100000;
        weights1[2392] <= 16'b1111111111000111;
        weights1[2393] <= 16'b1111111111000000;
        weights1[2394] <= 16'b1111111111000011;
        weights1[2395] <= 16'b1111111111100001;
        weights1[2396] <= 16'b1111111111111011;
        weights1[2397] <= 16'b0000000000101111;
        weights1[2398] <= 16'b0000000000100101;
        weights1[2399] <= 16'b0000000000100001;
        weights1[2400] <= 16'b0000000000010011;
        weights1[2401] <= 16'b0000000000001100;
        weights1[2402] <= 16'b0000000000001101;
        weights1[2403] <= 16'b0000000000000010;
        weights1[2404] <= 16'b1111111111101101;
        weights1[2405] <= 16'b1111111111110111;
        weights1[2406] <= 16'b1111111111111011;
        weights1[2407] <= 16'b1111111111111110;
        weights1[2408] <= 16'b0000000000000000;
        weights1[2409] <= 16'b0000000000000000;
        weights1[2410] <= 16'b0000000000000001;
        weights1[2411] <= 16'b1111111111111011;
        weights1[2412] <= 16'b1111111111110110;
        weights1[2413] <= 16'b1111111111111010;
        weights1[2414] <= 16'b1111111111111011;
        weights1[2415] <= 16'b1111111111111001;
        weights1[2416] <= 16'b0000000000010011;
        weights1[2417] <= 16'b0000000000001001;
        weights1[2418] <= 16'b1111111111011110;
        weights1[2419] <= 16'b1111111111100101;
        weights1[2420] <= 16'b1111111110111111;
        weights1[2421] <= 16'b1111111110011001;
        weights1[2422] <= 16'b1111111110011000;
        weights1[2423] <= 16'b1111111111001111;
        weights1[2424] <= 16'b0000000000011110;
        weights1[2425] <= 16'b0000000000011101;
        weights1[2426] <= 16'b0000000000010010;
        weights1[2427] <= 16'b0000000000001010;
        weights1[2428] <= 16'b0000000000010011;
        weights1[2429] <= 16'b1111111111110111;
        weights1[2430] <= 16'b1111111111110100;
        weights1[2431] <= 16'b1111111111101000;
        weights1[2432] <= 16'b1111111111101011;
        weights1[2433] <= 16'b1111111111110011;
        weights1[2434] <= 16'b1111111111110001;
        weights1[2435] <= 16'b1111111111111000;
        weights1[2436] <= 16'b0000000000000001;
        weights1[2437] <= 16'b0000000000000001;
        weights1[2438] <= 16'b0000000000000011;
        weights1[2439] <= 16'b0000000000000000;
        weights1[2440] <= 16'b1111111111111000;
        weights1[2441] <= 16'b1111111111111111;
        weights1[2442] <= 16'b1111111111111010;
        weights1[2443] <= 16'b1111111111111100;
        weights1[2444] <= 16'b0000000000000110;
        weights1[2445] <= 16'b0000000000000011;
        weights1[2446] <= 16'b1111111111110111;
        weights1[2447] <= 16'b1111111111100100;
        weights1[2448] <= 16'b1111111111001000;
        weights1[2449] <= 16'b1111111101111111;
        weights1[2450] <= 16'b1111111110000101;
        weights1[2451] <= 16'b1111111111000011;
        weights1[2452] <= 16'b1111111111010111;
        weights1[2453] <= 16'b0000000000011001;
        weights1[2454] <= 16'b0000000000001100;
        weights1[2455] <= 16'b0000000000010100;
        weights1[2456] <= 16'b1111111111011110;
        weights1[2457] <= 16'b1111111111101000;
        weights1[2458] <= 16'b0000000000001010;
        weights1[2459] <= 16'b1111111111101001;
        weights1[2460] <= 16'b1111111111100110;
        weights1[2461] <= 16'b1111111111100100;
        weights1[2462] <= 16'b1111111111100110;
        weights1[2463] <= 16'b1111111111110111;
        weights1[2464] <= 16'b0000000000000100;
        weights1[2465] <= 16'b0000000000000100;
        weights1[2466] <= 16'b0000000000000000;
        weights1[2467] <= 16'b0000000000000001;
        weights1[2468] <= 16'b1111111111111001;
        weights1[2469] <= 16'b1111111111111011;
        weights1[2470] <= 16'b1111111111110110;
        weights1[2471] <= 16'b0000000000000001;
        weights1[2472] <= 16'b1111111111111111;
        weights1[2473] <= 16'b0000000000010000;
        weights1[2474] <= 16'b1111111111110111;
        weights1[2475] <= 16'b1111111111110100;
        weights1[2476] <= 16'b1111111111001111;
        weights1[2477] <= 16'b1111111101111001;
        weights1[2478] <= 16'b1111111101100101;
        weights1[2479] <= 16'b1111111110110000;
        weights1[2480] <= 16'b0000000000010001;
        weights1[2481] <= 16'b0000000000000111;
        weights1[2482] <= 16'b0000000000001010;
        weights1[2483] <= 16'b1111111111111001;
        weights1[2484] <= 16'b0000000000001110;
        weights1[2485] <= 16'b1111111111111110;
        weights1[2486] <= 16'b1111111111101010;
        weights1[2487] <= 16'b1111111111110111;
        weights1[2488] <= 16'b1111111111001110;
        weights1[2489] <= 16'b1111111111011111;
        weights1[2490] <= 16'b1111111111100101;
        weights1[2491] <= 16'b1111111111110010;
        weights1[2492] <= 16'b0000000000001000;
        weights1[2493] <= 16'b0000000000000001;
        weights1[2494] <= 16'b0000000000000000;
        weights1[2495] <= 16'b0000000000001010;
        weights1[2496] <= 16'b1111111111110011;
        weights1[2497] <= 16'b1111111111111101;
        weights1[2498] <= 16'b0000000000000100;
        weights1[2499] <= 16'b0000000000000001;
        weights1[2500] <= 16'b0000000000000001;
        weights1[2501] <= 16'b0000000000000001;
        weights1[2502] <= 16'b0000000000010001;
        weights1[2503] <= 16'b1111111111111101;
        weights1[2504] <= 16'b1111111111000001;
        weights1[2505] <= 16'b1111111101100000;
        weights1[2506] <= 16'b1111111101000110;
        weights1[2507] <= 16'b1111111110100000;
        weights1[2508] <= 16'b0000000000110001;
        weights1[2509] <= 16'b0000000000111100;
        weights1[2510] <= 16'b0000000000100111;
        weights1[2511] <= 16'b1111111111111110;
        weights1[2512] <= 16'b0000000000001001;
        weights1[2513] <= 16'b0000000000010010;
        weights1[2514] <= 16'b0000000000000001;
        weights1[2515] <= 16'b1111111111001000;
        weights1[2516] <= 16'b1111111111001010;
        weights1[2517] <= 16'b1111111111010110;
        weights1[2518] <= 16'b1111111111101010;
        weights1[2519] <= 16'b1111111111110100;
        weights1[2520] <= 16'b0000000000000100;
        weights1[2521] <= 16'b1111111111111101;
        weights1[2522] <= 16'b1111111111111111;
        weights1[2523] <= 16'b1111111111111011;
        weights1[2524] <= 16'b0000000000000000;
        weights1[2525] <= 16'b0000000000000010;
        weights1[2526] <= 16'b1111111111111111;
        weights1[2527] <= 16'b1111111111111000;
        weights1[2528] <= 16'b0000000000000011;
        weights1[2529] <= 16'b0000000000011011;
        weights1[2530] <= 16'b0000000000010100;
        weights1[2531] <= 16'b0000000000000110;
        weights1[2532] <= 16'b1111111111010100;
        weights1[2533] <= 16'b1111111101110001;
        weights1[2534] <= 16'b1111111100000100;
        weights1[2535] <= 16'b1111111111000111;
        weights1[2536] <= 16'b0000000000010111;
        weights1[2537] <= 16'b0000000000110011;
        weights1[2538] <= 16'b0000000000010011;
        weights1[2539] <= 16'b0000000000001010;
        weights1[2540] <= 16'b0000000000101111;
        weights1[2541] <= 16'b1111111111111111;
        weights1[2542] <= 16'b1111111111100101;
        weights1[2543] <= 16'b1111111111001000;
        weights1[2544] <= 16'b1111111111001011;
        weights1[2545] <= 16'b1111111111010000;
        weights1[2546] <= 16'b1111111111011110;
        weights1[2547] <= 16'b1111111111101101;
        weights1[2548] <= 16'b1111111111111110;
        weights1[2549] <= 16'b1111111111111011;
        weights1[2550] <= 16'b1111111111111100;
        weights1[2551] <= 16'b0000000000000111;
        weights1[2552] <= 16'b1111111111101001;
        weights1[2553] <= 16'b0000000000011000;
        weights1[2554] <= 16'b0000000000000110;
        weights1[2555] <= 16'b0000000000010101;
        weights1[2556] <= 16'b0000000000010100;
        weights1[2557] <= 16'b0000000000010010;
        weights1[2558] <= 16'b0000000000100011;
        weights1[2559] <= 16'b0000000000100000;
        weights1[2560] <= 16'b1111111111100101;
        weights1[2561] <= 16'b1111111101000010;
        weights1[2562] <= 16'b1111111011110010;
        weights1[2563] <= 16'b1111111111111111;
        weights1[2564] <= 16'b0000000000111100;
        weights1[2565] <= 16'b0000000000101100;
        weights1[2566] <= 16'b0000000000001001;
        weights1[2567] <= 16'b0000000000010111;
        weights1[2568] <= 16'b0000000000000011;
        weights1[2569] <= 16'b0000000000000111;
        weights1[2570] <= 16'b1111111111010100;
        weights1[2571] <= 16'b1111111110111001;
        weights1[2572] <= 16'b1111111110111111;
        weights1[2573] <= 16'b1111111111010011;
        weights1[2574] <= 16'b1111111111100001;
        weights1[2575] <= 16'b1111111111110101;
        weights1[2576] <= 16'b1111111111111111;
        weights1[2577] <= 16'b1111111111111100;
        weights1[2578] <= 16'b1111111111111101;
        weights1[2579] <= 16'b1111111111111110;
        weights1[2580] <= 16'b1111111111111101;
        weights1[2581] <= 16'b0000000000000110;
        weights1[2582] <= 16'b0000000000100010;
        weights1[2583] <= 16'b0000000000000111;
        weights1[2584] <= 16'b1111111111110011;
        weights1[2585] <= 16'b0000000000101001;
        weights1[2586] <= 16'b0000000000000010;
        weights1[2587] <= 16'b0000000000101101;
        weights1[2588] <= 16'b1111111111100100;
        weights1[2589] <= 16'b1111111101000010;
        weights1[2590] <= 16'b1111111101010010;
        weights1[2591] <= 16'b0000000000100011;
        weights1[2592] <= 16'b0000000000100010;
        weights1[2593] <= 16'b0000000000101001;
        weights1[2594] <= 16'b0000000000100101;
        weights1[2595] <= 16'b0000000000000010;
        weights1[2596] <= 16'b0000000000010111;
        weights1[2597] <= 16'b0000000000000010;
        weights1[2598] <= 16'b1111111110111101;
        weights1[2599] <= 16'b1111111110101111;
        weights1[2600] <= 16'b1111111110101111;
        weights1[2601] <= 16'b1111111111010100;
        weights1[2602] <= 16'b1111111111100111;
        weights1[2603] <= 16'b0000000000000000;
        weights1[2604] <= 16'b1111111111111101;
        weights1[2605] <= 16'b1111111111111100;
        weights1[2606] <= 16'b1111111111111100;
        weights1[2607] <= 16'b1111111111111111;
        weights1[2608] <= 16'b1111111111110110;
        weights1[2609] <= 16'b1111111111111110;
        weights1[2610] <= 16'b1111111111111010;
        weights1[2611] <= 16'b1111111111110110;
        weights1[2612] <= 16'b0000000000011010;
        weights1[2613] <= 16'b0000000000001111;
        weights1[2614] <= 16'b0000000000101101;
        weights1[2615] <= 16'b0000000000101010;
        weights1[2616] <= 16'b1111111111011001;
        weights1[2617] <= 16'b1111111101000101;
        weights1[2618] <= 16'b1111111110001101;
        weights1[2619] <= 16'b0000000000001110;
        weights1[2620] <= 16'b0000000000100011;
        weights1[2621] <= 16'b0000000000010100;
        weights1[2622] <= 16'b0000000000011100;
        weights1[2623] <= 16'b0000000000010101;
        weights1[2624] <= 16'b0000000000010001;
        weights1[2625] <= 16'b1111111111111000;
        weights1[2626] <= 16'b1111111110011101;
        weights1[2627] <= 16'b1111111111001101;
        weights1[2628] <= 16'b1111111111010011;
        weights1[2629] <= 16'b1111111111101111;
        weights1[2630] <= 16'b1111111111111111;
        weights1[2631] <= 16'b0000000000011000;
        weights1[2632] <= 16'b1111111111111110;
        weights1[2633] <= 16'b0000000000000101;
        weights1[2634] <= 16'b1111111111111000;
        weights1[2635] <= 16'b0000000000000000;
        weights1[2636] <= 16'b1111111111111000;
        weights1[2637] <= 16'b1111111111110100;
        weights1[2638] <= 16'b1111111111101110;
        weights1[2639] <= 16'b0000000000011011;
        weights1[2640] <= 16'b1111111111111101;
        weights1[2641] <= 16'b0000000000000000;
        weights1[2642] <= 16'b0000000000101010;
        weights1[2643] <= 16'b0000000000110110;
        weights1[2644] <= 16'b1111111111010100;
        weights1[2645] <= 16'b1111111101111000;
        weights1[2646] <= 16'b1111111111010100;
        weights1[2647] <= 16'b0000000000001101;
        weights1[2648] <= 16'b0000000000010111;
        weights1[2649] <= 16'b0000000000100001;
        weights1[2650] <= 16'b0000000000001110;
        weights1[2651] <= 16'b0000000000010001;
        weights1[2652] <= 16'b1111111111100110;
        weights1[2653] <= 16'b1111111110111111;
        weights1[2654] <= 16'b1111111110111011;
        weights1[2655] <= 16'b1111111111000011;
        weights1[2656] <= 16'b1111111111101000;
        weights1[2657] <= 16'b0000000000010110;
        weights1[2658] <= 16'b0000000000100111;
        weights1[2659] <= 16'b0000000000100111;
        weights1[2660] <= 16'b0000000000000100;
        weights1[2661] <= 16'b0000000000000110;
        weights1[2662] <= 16'b1111111111101111;
        weights1[2663] <= 16'b1111111111111110;
        weights1[2664] <= 16'b1111111111111101;
        weights1[2665] <= 16'b0000000000000000;
        weights1[2666] <= 16'b1111111111111000;
        weights1[2667] <= 16'b0000000000000010;
        weights1[2668] <= 16'b0000000000001000;
        weights1[2669] <= 16'b0000000000100001;
        weights1[2670] <= 16'b0000000000100101;
        weights1[2671] <= 16'b0000000000011101;
        weights1[2672] <= 16'b1111111111010000;
        weights1[2673] <= 16'b1111111110101110;
        weights1[2674] <= 16'b1111111111011011;
        weights1[2675] <= 16'b0000000000001011;
        weights1[2676] <= 16'b0000000000011100;
        weights1[2677] <= 16'b0000000000011110;
        weights1[2678] <= 16'b0000000000100000;
        weights1[2679] <= 16'b1111111111101011;
        weights1[2680] <= 16'b0000000000000001;
        weights1[2681] <= 16'b1111111111000011;
        weights1[2682] <= 16'b1111111111000010;
        weights1[2683] <= 16'b1111111111001011;
        weights1[2684] <= 16'b0000000000000001;
        weights1[2685] <= 16'b0000000000110000;
        weights1[2686] <= 16'b0000000000101010;
        weights1[2687] <= 16'b0000000000011111;
        weights1[2688] <= 16'b1111111111111101;
        weights1[2689] <= 16'b0000000000001010;
        weights1[2690] <= 16'b0000000000001010;
        weights1[2691] <= 16'b0000000000010111;
        weights1[2692] <= 16'b0000000000000100;
        weights1[2693] <= 16'b0000000000000111;
        weights1[2694] <= 16'b0000000000000010;
        weights1[2695] <= 16'b0000000000101011;
        weights1[2696] <= 16'b1111111111110100;
        weights1[2697] <= 16'b0000000000001101;
        weights1[2698] <= 16'b0000000000100011;
        weights1[2699] <= 16'b0000000000011110;
        weights1[2700] <= 16'b1111111111011111;
        weights1[2701] <= 16'b1111111111001011;
        weights1[2702] <= 16'b1111111111011001;
        weights1[2703] <= 16'b0000000000000010;
        weights1[2704] <= 16'b0000000000001110;
        weights1[2705] <= 16'b0000000000100011;
        weights1[2706] <= 16'b1111111111111000;
        weights1[2707] <= 16'b1111111111111111;
        weights1[2708] <= 16'b1111111111111010;
        weights1[2709] <= 16'b1111111111000101;
        weights1[2710] <= 16'b1111111111100011;
        weights1[2711] <= 16'b1111111111111011;
        weights1[2712] <= 16'b0000000000110111;
        weights1[2713] <= 16'b0000000000011111;
        weights1[2714] <= 16'b0000000000011101;
        weights1[2715] <= 16'b0000000000001001;
        weights1[2716] <= 16'b1111111111111111;
        weights1[2717] <= 16'b0000000000001111;
        weights1[2718] <= 16'b0000000000001011;
        weights1[2719] <= 16'b1111111111111100;
        weights1[2720] <= 16'b0000000000001010;
        weights1[2721] <= 16'b0000000000001010;
        weights1[2722] <= 16'b0000000000010000;
        weights1[2723] <= 16'b1111111111100111;
        weights1[2724] <= 16'b0000000000001100;
        weights1[2725] <= 16'b0000000000000100;
        weights1[2726] <= 16'b0000000000010100;
        weights1[2727] <= 16'b0000000000100010;
        weights1[2728] <= 16'b1111111111111100;
        weights1[2729] <= 16'b1111111111101000;
        weights1[2730] <= 16'b1111111111111000;
        weights1[2731] <= 16'b1111111111111010;
        weights1[2732] <= 16'b1111111111111011;
        weights1[2733] <= 16'b0000000000000000;
        weights1[2734] <= 16'b1111111111111010;
        weights1[2735] <= 16'b1111111111111110;
        weights1[2736] <= 16'b1111111111011110;
        weights1[2737] <= 16'b1111111111011010;
        weights1[2738] <= 16'b1111111111011011;
        weights1[2739] <= 16'b0000000000001101;
        weights1[2740] <= 16'b0000000000011011;
        weights1[2741] <= 16'b0000000000001011;
        weights1[2742] <= 16'b1111111111111101;
        weights1[2743] <= 16'b1111111111111111;
        weights1[2744] <= 16'b0000000000000000;
        weights1[2745] <= 16'b0000000000001010;
        weights1[2746] <= 16'b0000000000001101;
        weights1[2747] <= 16'b1111111111110100;
        weights1[2748] <= 16'b1111111111110100;
        weights1[2749] <= 16'b1111111111111010;
        weights1[2750] <= 16'b1111111111101000;
        weights1[2751] <= 16'b0000000000000011;
        weights1[2752] <= 16'b0000000000010000;
        weights1[2753] <= 16'b0000000000000101;
        weights1[2754] <= 16'b0000000000001011;
        weights1[2755] <= 16'b0000000000011011;
        weights1[2756] <= 16'b0000000000001100;
        weights1[2757] <= 16'b1111111111101001;
        weights1[2758] <= 16'b1111111111101010;
        weights1[2759] <= 16'b0000000000000100;
        weights1[2760] <= 16'b0000000000001100;
        weights1[2761] <= 16'b0000000000001001;
        weights1[2762] <= 16'b0000000000000011;
        weights1[2763] <= 16'b1111111111111010;
        weights1[2764] <= 16'b1111111111100001;
        weights1[2765] <= 16'b1111111111110001;
        weights1[2766] <= 16'b0000000000000001;
        weights1[2767] <= 16'b0000000000010000;
        weights1[2768] <= 16'b0000000000010001;
        weights1[2769] <= 16'b0000000000010001;
        weights1[2770] <= 16'b0000000000000101;
        weights1[2771] <= 16'b1111111111110110;
        weights1[2772] <= 16'b0000000000001011;
        weights1[2773] <= 16'b0000000000001001;
        weights1[2774] <= 16'b0000000000001100;
        weights1[2775] <= 16'b1111111111111001;
        weights1[2776] <= 16'b0000000000001001;
        weights1[2777] <= 16'b0000000000000010;
        weights1[2778] <= 16'b0000000000010101;
        weights1[2779] <= 16'b0000000000000001;
        weights1[2780] <= 16'b0000000000001101;
        weights1[2781] <= 16'b0000000000001011;
        weights1[2782] <= 16'b0000000000000110;
        weights1[2783] <= 16'b0000000000001001;
        weights1[2784] <= 16'b0000000000000101;
        weights1[2785] <= 16'b0000000000001101;
        weights1[2786] <= 16'b1111111111110010;
        weights1[2787] <= 16'b1111111111111000;
        weights1[2788] <= 16'b0000000000000100;
        weights1[2789] <= 16'b0000000000000010;
        weights1[2790] <= 16'b1111111111110010;
        weights1[2791] <= 16'b0000000000000001;
        weights1[2792] <= 16'b1111111111101011;
        weights1[2793] <= 16'b1111111111110000;
        weights1[2794] <= 16'b0000000000010111;
        weights1[2795] <= 16'b0000000000011111;
        weights1[2796] <= 16'b1111111111111111;
        weights1[2797] <= 16'b1111111111110000;
        weights1[2798] <= 16'b1111111111111011;
        weights1[2799] <= 16'b1111111111111101;
        weights1[2800] <= 16'b0000000000000110;
        weights1[2801] <= 16'b0000000000000010;
        weights1[2802] <= 16'b0000000000000010;
        weights1[2803] <= 16'b1111111111111101;
        weights1[2804] <= 16'b1111111111111110;
        weights1[2805] <= 16'b1111111111111100;
        weights1[2806] <= 16'b0000000000000110;
        weights1[2807] <= 16'b0000000000000100;
        weights1[2808] <= 16'b1111111111110100;
        weights1[2809] <= 16'b1111111111111111;
        weights1[2810] <= 16'b0000000000001010;
        weights1[2811] <= 16'b0000000000000101;
        weights1[2812] <= 16'b0000000000000110;
        weights1[2813] <= 16'b0000000000000011;
        weights1[2814] <= 16'b0000000000001101;
        weights1[2815] <= 16'b0000000000000001;
        weights1[2816] <= 16'b1111111111101111;
        weights1[2817] <= 16'b1111111111111010;
        weights1[2818] <= 16'b1111111111110011;
        weights1[2819] <= 16'b1111111111111100;
        weights1[2820] <= 16'b0000000000000000;
        weights1[2821] <= 16'b1111111111111111;
        weights1[2822] <= 16'b1111111111111010;
        weights1[2823] <= 16'b0000000000000111;
        weights1[2824] <= 16'b0000000000000001;
        weights1[2825] <= 16'b1111111111101101;
        weights1[2826] <= 16'b1111111111111001;
        weights1[2827] <= 16'b1111111111111101;
        weights1[2828] <= 16'b0000000000000101;
        weights1[2829] <= 16'b0000000000000101;
        weights1[2830] <= 16'b0000000000001001;
        weights1[2831] <= 16'b1111111111110110;
        weights1[2832] <= 16'b0000000000000111;
        weights1[2833] <= 16'b0000000000100101;
        weights1[2834] <= 16'b1111111111101111;
        weights1[2835] <= 16'b0000000000010000;
        weights1[2836] <= 16'b1111111111101011;
        weights1[2837] <= 16'b1111111111111010;
        weights1[2838] <= 16'b0000000000000001;
        weights1[2839] <= 16'b0000000000000101;
        weights1[2840] <= 16'b0000000000000011;
        weights1[2841] <= 16'b1111111111110111;
        weights1[2842] <= 16'b0000000000000000;
        weights1[2843] <= 16'b1111111111110111;
        weights1[2844] <= 16'b1111111111111011;
        weights1[2845] <= 16'b1111111111110010;
        weights1[2846] <= 16'b1111111111111001;
        weights1[2847] <= 16'b1111111111111010;
        weights1[2848] <= 16'b0000000000001110;
        weights1[2849] <= 16'b0000000000001011;
        weights1[2850] <= 16'b0000000000000010;
        weights1[2851] <= 16'b1111111111110110;
        weights1[2852] <= 16'b1111111111110000;
        weights1[2853] <= 16'b1111111111110001;
        weights1[2854] <= 16'b1111111111101111;
        weights1[2855] <= 16'b1111111111111001;
        weights1[2856] <= 16'b0000000000000011;
        weights1[2857] <= 16'b1111111111111110;
        weights1[2858] <= 16'b1111111111111010;
        weights1[2859] <= 16'b1111111111110101;
        weights1[2860] <= 16'b0000000000011011;
        weights1[2861] <= 16'b0000000000000001;
        weights1[2862] <= 16'b0000000000000101;
        weights1[2863] <= 16'b1111111111111100;
        weights1[2864] <= 16'b0000000000001010;
        weights1[2865] <= 16'b0000000000000111;
        weights1[2866] <= 16'b0000000000010101;
        weights1[2867] <= 16'b0000000000010010;
        weights1[2868] <= 16'b0000000000000011;
        weights1[2869] <= 16'b1111111111111011;
        weights1[2870] <= 16'b1111111111110010;
        weights1[2871] <= 16'b1111111111101010;
        weights1[2872] <= 16'b1111111111110001;
        weights1[2873] <= 16'b1111111111111011;
        weights1[2874] <= 16'b1111111111111101;
        weights1[2875] <= 16'b1111111111111001;
        weights1[2876] <= 16'b1111111111110100;
        weights1[2877] <= 16'b1111111111101010;
        weights1[2878] <= 16'b1111111111110010;
        weights1[2879] <= 16'b1111111111100111;
        weights1[2880] <= 16'b1111111111110101;
        weights1[2881] <= 16'b1111111111111100;
        weights1[2882] <= 16'b1111111111111011;
        weights1[2883] <= 16'b1111111111111000;
        weights1[2884] <= 16'b0000000000000000;
        weights1[2885] <= 16'b1111111111111011;
        weights1[2886] <= 16'b0000000000000000;
        weights1[2887] <= 16'b0000000000000101;
        weights1[2888] <= 16'b0000000000000010;
        weights1[2889] <= 16'b1111111111111011;
        weights1[2890] <= 16'b1111111111110110;
        weights1[2891] <= 16'b1111111111111110;
        weights1[2892] <= 16'b1111111111111111;
        weights1[2893] <= 16'b1111111111110101;
        weights1[2894] <= 16'b1111111111110110;
        weights1[2895] <= 16'b0000000000001000;
        weights1[2896] <= 16'b0000000000000001;
        weights1[2897] <= 16'b1111111111111000;
        weights1[2898] <= 16'b0000000000000110;
        weights1[2899] <= 16'b1111111111101101;
        weights1[2900] <= 16'b1111111111111111;
        weights1[2901] <= 16'b1111111111111000;
        weights1[2902] <= 16'b0000000000000010;
        weights1[2903] <= 16'b1111111111111110;
        weights1[2904] <= 16'b1111111111101111;
        weights1[2905] <= 16'b1111111111111100;
        weights1[2906] <= 16'b1111111111110110;
        weights1[2907] <= 16'b1111111111101101;
        weights1[2908] <= 16'b0000000000000110;
        weights1[2909] <= 16'b1111111111111111;
        weights1[2910] <= 16'b0000000000001000;
        weights1[2911] <= 16'b0000000000000101;
        weights1[2912] <= 16'b0000000000000101;
        weights1[2913] <= 16'b1111111111110111;
        weights1[2914] <= 16'b1111111111111100;
        weights1[2915] <= 16'b1111111111111111;
        weights1[2916] <= 16'b0000000000000000;
        weights1[2917] <= 16'b1111111111110011;
        weights1[2918] <= 16'b0000000000001001;
        weights1[2919] <= 16'b1111111111101100;
        weights1[2920] <= 16'b1111111111110010;
        weights1[2921] <= 16'b0000000000000101;
        weights1[2922] <= 16'b0000000000000010;
        weights1[2923] <= 16'b0000000000000101;
        weights1[2924] <= 16'b0000000000000111;
        weights1[2925] <= 16'b1111111111111011;
        weights1[2926] <= 16'b1111111111100011;
        weights1[2927] <= 16'b0000000000000010;
        weights1[2928] <= 16'b1111111111110101;
        weights1[2929] <= 16'b1111111111110110;
        weights1[2930] <= 16'b1111111111101111;
        weights1[2931] <= 16'b0000000000000011;
        weights1[2932] <= 16'b1111111111111000;
        weights1[2933] <= 16'b1111111111110001;
        weights1[2934] <= 16'b1111111111110100;
        weights1[2935] <= 16'b0000000000000111;
        weights1[2936] <= 16'b0000000000010001;
        weights1[2937] <= 16'b0000000000001111;
        weights1[2938] <= 16'b0000000000001001;
        weights1[2939] <= 16'b0000000000001100;
        weights1[2940] <= 16'b1111111111111101;
        weights1[2941] <= 16'b1111111111111111;
        weights1[2942] <= 16'b0000000000000110;
        weights1[2943] <= 16'b1111111111111011;
        weights1[2944] <= 16'b1111111111110000;
        weights1[2945] <= 16'b1111111111110100;
        weights1[2946] <= 16'b1111111111111110;
        weights1[2947] <= 16'b0000000000000100;
        weights1[2948] <= 16'b0000000000101111;
        weights1[2949] <= 16'b1111111111110111;
        weights1[2950] <= 16'b1111111111111000;
        weights1[2951] <= 16'b0000000000000100;
        weights1[2952] <= 16'b1111111111110101;
        weights1[2953] <= 16'b1111111111111111;
        weights1[2954] <= 16'b1111111111111011;
        weights1[2955] <= 16'b1111111111110111;
        weights1[2956] <= 16'b1111111111111000;
        weights1[2957] <= 16'b0000000000000001;
        weights1[2958] <= 16'b0000000000001011;
        weights1[2959] <= 16'b0000000000000100;
        weights1[2960] <= 16'b1111111111111011;
        weights1[2961] <= 16'b1111111111011101;
        weights1[2962] <= 16'b1111111111111010;
        weights1[2963] <= 16'b1111111111111110;
        weights1[2964] <= 16'b0000000000001100;
        weights1[2965] <= 16'b1111111111111011;
        weights1[2966] <= 16'b0000000000001000;
        weights1[2967] <= 16'b0000000000001001;
        weights1[2968] <= 16'b1111111111111011;
        weights1[2969] <= 16'b1111111111111001;
        weights1[2970] <= 16'b0000000000000110;
        weights1[2971] <= 16'b1111111111110101;
        weights1[2972] <= 16'b1111111111111011;
        weights1[2973] <= 16'b0000000000001011;
        weights1[2974] <= 16'b0000000000001000;
        weights1[2975] <= 16'b0000000000000011;
        weights1[2976] <= 16'b1111111111111010;
        weights1[2977] <= 16'b1111111111110111;
        weights1[2978] <= 16'b0000000000000001;
        weights1[2979] <= 16'b1111111111101100;
        weights1[2980] <= 16'b1111111111111111;
        weights1[2981] <= 16'b0000000000000111;
        weights1[2982] <= 16'b1111111111111110;
        weights1[2983] <= 16'b0000000000000000;
        weights1[2984] <= 16'b1111111111110110;
        weights1[2985] <= 16'b1111111111110000;
        weights1[2986] <= 16'b1111111111011101;
        weights1[2987] <= 16'b1111111111111101;
        weights1[2988] <= 16'b0000000000010000;
        weights1[2989] <= 16'b0000000000000001;
        weights1[2990] <= 16'b1111111111101110;
        weights1[2991] <= 16'b1111111111111010;
        weights1[2992] <= 16'b1111111111111101;
        weights1[2993] <= 16'b1111111111110100;
        weights1[2994] <= 16'b0000000000000011;
        weights1[2995] <= 16'b0000000000000010;
        weights1[2996] <= 16'b1111111111111001;
        weights1[2997] <= 16'b1111111111111011;
        weights1[2998] <= 16'b0000000000000010;
        weights1[2999] <= 16'b0000000000001000;
        weights1[3000] <= 16'b0000000000000000;
        weights1[3001] <= 16'b1111111111111010;
        weights1[3002] <= 16'b1111111111011011;
        weights1[3003] <= 16'b1111111111111110;
        weights1[3004] <= 16'b0000000000001110;
        weights1[3005] <= 16'b1111111111111000;
        weights1[3006] <= 16'b0000000000001100;
        weights1[3007] <= 16'b0000000000000110;
        weights1[3008] <= 16'b0000000000000000;
        weights1[3009] <= 16'b1111111111111110;
        weights1[3010] <= 16'b1111111111110001;
        weights1[3011] <= 16'b1111111111110111;
        weights1[3012] <= 16'b1111111111110011;
        weights1[3013] <= 16'b0000000000000111;
        weights1[3014] <= 16'b0000000000011001;
        weights1[3015] <= 16'b1111111111110101;
        weights1[3016] <= 16'b1111111111111011;
        weights1[3017] <= 16'b0000000000000111;
        weights1[3018] <= 16'b1111111111110100;
        weights1[3019] <= 16'b1111111111110010;
        weights1[3020] <= 16'b1111111111111000;
        weights1[3021] <= 16'b1111111111110111;
        weights1[3022] <= 16'b1111111111111110;
        weights1[3023] <= 16'b0000000000000010;
        weights1[3024] <= 16'b0000000000000001;
        weights1[3025] <= 16'b1111111111111011;
        weights1[3026] <= 16'b1111111111111110;
        weights1[3027] <= 16'b1111111111111101;
        weights1[3028] <= 16'b1111111111110111;
        weights1[3029] <= 16'b1111111111101100;
        weights1[3030] <= 16'b1111111111110010;
        weights1[3031] <= 16'b1111111111111000;
        weights1[3032] <= 16'b1111111111100110;
        weights1[3033] <= 16'b1111111111111010;
        weights1[3034] <= 16'b1111111111100101;
        weights1[3035] <= 16'b1111111111110111;
        weights1[3036] <= 16'b0000000000010110;
        weights1[3037] <= 16'b0000000000000011;
        weights1[3038] <= 16'b1111111111111000;
        weights1[3039] <= 16'b0000000000000101;
        weights1[3040] <= 16'b0000000000000101;
        weights1[3041] <= 16'b0000000000010110;
        weights1[3042] <= 16'b0000000000001101;
        weights1[3043] <= 16'b1111111111110100;
        weights1[3044] <= 16'b0000000000000110;
        weights1[3045] <= 16'b0000000000001010;
        weights1[3046] <= 16'b0000000000000100;
        weights1[3047] <= 16'b1111111111111001;
        weights1[3048] <= 16'b1111111111111101;
        weights1[3049] <= 16'b0000000000000001;
        weights1[3050] <= 16'b1111111111111101;
        weights1[3051] <= 16'b0000000000000001;
        weights1[3052] <= 16'b0000000000000000;
        weights1[3053] <= 16'b1111111111111100;
        weights1[3054] <= 16'b1111111111110110;
        weights1[3055] <= 16'b0000000000000010;
        weights1[3056] <= 16'b1111111111111001;
        weights1[3057] <= 16'b1111111111111110;
        weights1[3058] <= 16'b1111111111111101;
        weights1[3059] <= 16'b1111111111110011;
        weights1[3060] <= 16'b1111111111110011;
        weights1[3061] <= 16'b1111111111100001;
        weights1[3062] <= 16'b0000000000010001;
        weights1[3063] <= 16'b1111111111110101;
        weights1[3064] <= 16'b1111111111101011;
        weights1[3065] <= 16'b0000000000011011;
        weights1[3066] <= 16'b1111111111100111;
        weights1[3067] <= 16'b0000000000001001;
        weights1[3068] <= 16'b1111111111110111;
        weights1[3069] <= 16'b0000000000000100;
        weights1[3070] <= 16'b0000000000001001;
        weights1[3071] <= 16'b1111111111111100;
        weights1[3072] <= 16'b1111111111110001;
        weights1[3073] <= 16'b0000000000000111;
        weights1[3074] <= 16'b0000000000000101;
        weights1[3075] <= 16'b0000000000000111;
        weights1[3076] <= 16'b0000000000000011;
        weights1[3077] <= 16'b0000000000000011;
        weights1[3078] <= 16'b0000000000000001;
        weights1[3079] <= 16'b1111111111111111;
        weights1[3080] <= 16'b0000000000000000;
        weights1[3081] <= 16'b1111111111111110;
        weights1[3082] <= 16'b0000000000000000;
        weights1[3083] <= 16'b1111111111111111;
        weights1[3084] <= 16'b1111111111111111;
        weights1[3085] <= 16'b1111111111111001;
        weights1[3086] <= 16'b1111111111110111;
        weights1[3087] <= 16'b0000000000010000;
        weights1[3088] <= 16'b0000000000000000;
        weights1[3089] <= 16'b0000000000000011;
        weights1[3090] <= 16'b0000000000000010;
        weights1[3091] <= 16'b1111111111111011;
        weights1[3092] <= 16'b1111111111111110;
        weights1[3093] <= 16'b1111111111111000;
        weights1[3094] <= 16'b1111111111110100;
        weights1[3095] <= 16'b0000000000000000;
        weights1[3096] <= 16'b1111111111110111;
        weights1[3097] <= 16'b0000000000000100;
        weights1[3098] <= 16'b0000000000000000;
        weights1[3099] <= 16'b0000000000000101;
        weights1[3100] <= 16'b0000000000010100;
        weights1[3101] <= 16'b1111111111111011;
        weights1[3102] <= 16'b0000000000010000;
        weights1[3103] <= 16'b0000000000001011;
        weights1[3104] <= 16'b0000000000000100;
        weights1[3105] <= 16'b0000000000001000;
        weights1[3106] <= 16'b0000000000000010;
        weights1[3107] <= 16'b1111111111111111;
        weights1[3108] <= 16'b0000000000000000;
        weights1[3109] <= 16'b0000000000000010;
        weights1[3110] <= 16'b0000000000000101;
        weights1[3111] <= 16'b0000000000001000;
        weights1[3112] <= 16'b0000000000001000;
        weights1[3113] <= 16'b1111111111110010;
        weights1[3114] <= 16'b1111111111110001;
        weights1[3115] <= 16'b1111111111110100;
        weights1[3116] <= 16'b1111111111111100;
        weights1[3117] <= 16'b1111111111111011;
        weights1[3118] <= 16'b0000000000001000;
        weights1[3119] <= 16'b1111111111111000;
        weights1[3120] <= 16'b1111111111111110;
        weights1[3121] <= 16'b0000000000001010;
        weights1[3122] <= 16'b1111111111111100;
        weights1[3123] <= 16'b0000000000000111;
        weights1[3124] <= 16'b0000000000010000;
        weights1[3125] <= 16'b1111111111111011;
        weights1[3126] <= 16'b1111111111111101;
        weights1[3127] <= 16'b0000000000000111;
        weights1[3128] <= 16'b0000000000000100;
        weights1[3129] <= 16'b1111111111110101;
        weights1[3130] <= 16'b0000000000000111;
        weights1[3131] <= 16'b0000000000001000;
        weights1[3132] <= 16'b0000000000000101;
        weights1[3133] <= 16'b0000000000000110;
        weights1[3134] <= 16'b0000000000000001;
        weights1[3135] <= 16'b0000000000000001;
        weights1[3136] <= 16'b1111111111111111;
        weights1[3137] <= 16'b1111111111111111;
        weights1[3138] <= 16'b1111111111111110;
        weights1[3139] <= 16'b0000000000000000;
        weights1[3140] <= 16'b1111111111111110;
        weights1[3141] <= 16'b1111111111111100;
        weights1[3142] <= 16'b0000000000000011;
        weights1[3143] <= 16'b1111111111111110;
        weights1[3144] <= 16'b1111111111111001;
        weights1[3145] <= 16'b1111111111110001;
        weights1[3146] <= 16'b1111111111110010;
        weights1[3147] <= 16'b1111111111110000;
        weights1[3148] <= 16'b1111111111101010;
        weights1[3149] <= 16'b1111111111110001;
        weights1[3150] <= 16'b1111111111101100;
        weights1[3151] <= 16'b1111111111101100;
        weights1[3152] <= 16'b1111111111101001;
        weights1[3153] <= 16'b1111111111101100;
        weights1[3154] <= 16'b1111111111110010;
        weights1[3155] <= 16'b1111111111110110;
        weights1[3156] <= 16'b1111111111110100;
        weights1[3157] <= 16'b1111111111110101;
        weights1[3158] <= 16'b1111111111110111;
        weights1[3159] <= 16'b1111111111111110;
        weights1[3160] <= 16'b1111111111111110;
        weights1[3161] <= 16'b1111111111111111;
        weights1[3162] <= 16'b1111111111111111;
        weights1[3163] <= 16'b1111111111111111;
        weights1[3164] <= 16'b1111111111111111;
        weights1[3165] <= 16'b1111111111111111;
        weights1[3166] <= 16'b1111111111111111;
        weights1[3167] <= 16'b1111111111111111;
        weights1[3168] <= 16'b0000000000000001;
        weights1[3169] <= 16'b0000000000000000;
        weights1[3170] <= 16'b0000000000001100;
        weights1[3171] <= 16'b0000000000000011;
        weights1[3172] <= 16'b1111111111110110;
        weights1[3173] <= 16'b1111111111110110;
        weights1[3174] <= 16'b1111111111110011;
        weights1[3175] <= 16'b1111111111110001;
        weights1[3176] <= 16'b1111111111110011;
        weights1[3177] <= 16'b1111111111100111;
        weights1[3178] <= 16'b1111111111110001;
        weights1[3179] <= 16'b1111111111101100;
        weights1[3180] <= 16'b1111111111110101;
        weights1[3181] <= 16'b1111111111100100;
        weights1[3182] <= 16'b1111111111111000;
        weights1[3183] <= 16'b1111111111101110;
        weights1[3184] <= 16'b1111111111101111;
        weights1[3185] <= 16'b1111111111101111;
        weights1[3186] <= 16'b1111111111110010;
        weights1[3187] <= 16'b1111111111110110;
        weights1[3188] <= 16'b1111111111111010;
        weights1[3189] <= 16'b1111111111111110;
        weights1[3190] <= 16'b1111111111111110;
        weights1[3191] <= 16'b1111111111111110;
        weights1[3192] <= 16'b1111111111111111;
        weights1[3193] <= 16'b1111111111111110;
        weights1[3194] <= 16'b1111111111111111;
        weights1[3195] <= 16'b1111111111111100;
        weights1[3196] <= 16'b1111111111111110;
        weights1[3197] <= 16'b0000000000000001;
        weights1[3198] <= 16'b0000000000000101;
        weights1[3199] <= 16'b0000000000001010;
        weights1[3200] <= 16'b1111111111111101;
        weights1[3201] <= 16'b1111111111110101;
        weights1[3202] <= 16'b1111111111111010;
        weights1[3203] <= 16'b1111111111111100;
        weights1[3204] <= 16'b1111111111111011;
        weights1[3205] <= 16'b1111111111111110;
        weights1[3206] <= 16'b0000000000000101;
        weights1[3207] <= 16'b1111111111110111;
        weights1[3208] <= 16'b1111111111110110;
        weights1[3209] <= 16'b1111111111101011;
        weights1[3210] <= 16'b1111111111110100;
        weights1[3211] <= 16'b1111111111110010;
        weights1[3212] <= 16'b1111111111101010;
        weights1[3213] <= 16'b1111111111100101;
        weights1[3214] <= 16'b1111111111101001;
        weights1[3215] <= 16'b1111111111101111;
        weights1[3216] <= 16'b1111111111110100;
        weights1[3217] <= 16'b1111111111111001;
        weights1[3218] <= 16'b1111111111111100;
        weights1[3219] <= 16'b1111111111111100;
        weights1[3220] <= 16'b0000000000000010;
        weights1[3221] <= 16'b0000000000000000;
        weights1[3222] <= 16'b1111111111111101;
        weights1[3223] <= 16'b1111111111111001;
        weights1[3224] <= 16'b1111111111111010;
        weights1[3225] <= 16'b1111111111111011;
        weights1[3226] <= 16'b0000000000000010;
        weights1[3227] <= 16'b0000000000000111;
        weights1[3228] <= 16'b0000000000000010;
        weights1[3229] <= 16'b1111111111111110;
        weights1[3230] <= 16'b0000000000001111;
        weights1[3231] <= 16'b0000000000000100;
        weights1[3232] <= 16'b1111111111100101;
        weights1[3233] <= 16'b1111111111110111;
        weights1[3234] <= 16'b1111111111011110;
        weights1[3235] <= 16'b1111111111110010;
        weights1[3236] <= 16'b1111111111011011;
        weights1[3237] <= 16'b1111111111010100;
        weights1[3238] <= 16'b1111111111011101;
        weights1[3239] <= 16'b1111111111100111;
        weights1[3240] <= 16'b1111111111001010;
        weights1[3241] <= 16'b1111111111011011;
        weights1[3242] <= 16'b1111111111011101;
        weights1[3243] <= 16'b1111111111100101;
        weights1[3244] <= 16'b1111111111110000;
        weights1[3245] <= 16'b1111111111110101;
        weights1[3246] <= 16'b1111111111110010;
        weights1[3247] <= 16'b1111111111110111;
        weights1[3248] <= 16'b0000000000000010;
        weights1[3249] <= 16'b0000000000000001;
        weights1[3250] <= 16'b1111111111111100;
        weights1[3251] <= 16'b1111111111111100;
        weights1[3252] <= 16'b1111111111110010;
        weights1[3253] <= 16'b0000000000000000;
        weights1[3254] <= 16'b0000000000000001;
        weights1[3255] <= 16'b1111111111111000;
        weights1[3256] <= 16'b1111111111111010;
        weights1[3257] <= 16'b1111111111110110;
        weights1[3258] <= 16'b1111111111011111;
        weights1[3259] <= 16'b1111111111010000;
        weights1[3260] <= 16'b1111111111110011;
        weights1[3261] <= 16'b1111111111010011;
        weights1[3262] <= 16'b0000000000000000;
        weights1[3263] <= 16'b1111111111100110;
        weights1[3264] <= 16'b1111111111100110;
        weights1[3265] <= 16'b0000000000001011;
        weights1[3266] <= 16'b1111111111101011;
        weights1[3267] <= 16'b1111111111100011;
        weights1[3268] <= 16'b0000000000000101;
        weights1[3269] <= 16'b0000000000001011;
        weights1[3270] <= 16'b1111111111100111;
        weights1[3271] <= 16'b1111111111011110;
        weights1[3272] <= 16'b1111111111100110;
        weights1[3273] <= 16'b1111111111111101;
        weights1[3274] <= 16'b1111111111111001;
        weights1[3275] <= 16'b1111111111111001;
        weights1[3276] <= 16'b0000000000000011;
        weights1[3277] <= 16'b1111111111111101;
        weights1[3278] <= 16'b1111111111111000;
        weights1[3279] <= 16'b0000000000000101;
        weights1[3280] <= 16'b0000000000001001;
        weights1[3281] <= 16'b1111111111011110;
        weights1[3282] <= 16'b1111111111100110;
        weights1[3283] <= 16'b1111111111110101;
        weights1[3284] <= 16'b1111111111111011;
        weights1[3285] <= 16'b0000000000001100;
        weights1[3286] <= 16'b1111111111111011;
        weights1[3287] <= 16'b0000000000010010;
        weights1[3288] <= 16'b1111111111101111;
        weights1[3289] <= 16'b1111111111111000;
        weights1[3290] <= 16'b1111111111111110;
        weights1[3291] <= 16'b1111111111101110;
        weights1[3292] <= 16'b0000000000000111;
        weights1[3293] <= 16'b1111111111111100;
        weights1[3294] <= 16'b0000000000000000;
        weights1[3295] <= 16'b1111111111011000;
        weights1[3296] <= 16'b1111111111110111;
        weights1[3297] <= 16'b1111111111100001;
        weights1[3298] <= 16'b1111111111110010;
        weights1[3299] <= 16'b1111111111010101;
        weights1[3300] <= 16'b1111111111111110;
        weights1[3301] <= 16'b1111111111111100;
        weights1[3302] <= 16'b1111111111111001;
        weights1[3303] <= 16'b1111111111111000;
        weights1[3304] <= 16'b1111111111111110;
        weights1[3305] <= 16'b1111111111111111;
        weights1[3306] <= 16'b0000000000000000;
        weights1[3307] <= 16'b0000000000000001;
        weights1[3308] <= 16'b1111111111110011;
        weights1[3309] <= 16'b0000000000000100;
        weights1[3310] <= 16'b1111111111101110;
        weights1[3311] <= 16'b0000000000000101;
        weights1[3312] <= 16'b1111111111110011;
        weights1[3313] <= 16'b1111111111111000;
        weights1[3314] <= 16'b0000000000000100;
        weights1[3315] <= 16'b1111111111011010;
        weights1[3316] <= 16'b1111111111111100;
        weights1[3317] <= 16'b1111111111110111;
        weights1[3318] <= 16'b0000000000001000;
        weights1[3319] <= 16'b1111111111100101;
        weights1[3320] <= 16'b0000000000000110;
        weights1[3321] <= 16'b0000000000000110;
        weights1[3322] <= 16'b1111111111101100;
        weights1[3323] <= 16'b1111111111111011;
        weights1[3324] <= 16'b1111111111100111;
        weights1[3325] <= 16'b1111111111110100;
        weights1[3326] <= 16'b1111111111101100;
        weights1[3327] <= 16'b1111111111011100;
        weights1[3328] <= 16'b1111111111101110;
        weights1[3329] <= 16'b1111111111011110;
        weights1[3330] <= 16'b1111111111100001;
        weights1[3331] <= 16'b1111111111101111;
        weights1[3332] <= 16'b1111111111111111;
        weights1[3333] <= 16'b0000000000000011;
        weights1[3334] <= 16'b0000000000001011;
        weights1[3335] <= 16'b1111111111101010;
        weights1[3336] <= 16'b1111111111101110;
        weights1[3337] <= 16'b1111111111101001;
        weights1[3338] <= 16'b1111111111111101;
        weights1[3339] <= 16'b1111111111110010;
        weights1[3340] <= 16'b0000000000011101;
        weights1[3341] <= 16'b0000000000000010;
        weights1[3342] <= 16'b1111111111011100;
        weights1[3343] <= 16'b1111111111110011;
        weights1[3344] <= 16'b1111111111110111;
        weights1[3345] <= 16'b1111111111111101;
        weights1[3346] <= 16'b1111111111101011;
        weights1[3347] <= 16'b1111111111101011;
        weights1[3348] <= 16'b1111111111111001;
        weights1[3349] <= 16'b1111111111011011;
        weights1[3350] <= 16'b1111111111101111;
        weights1[3351] <= 16'b1111111111101000;
        weights1[3352] <= 16'b1111111111101111;
        weights1[3353] <= 16'b1111111111111111;
        weights1[3354] <= 16'b1111111111101101;
        weights1[3355] <= 16'b1111111111011110;
        weights1[3356] <= 16'b1111111111101010;
        weights1[3357] <= 16'b1111111111010110;
        weights1[3358] <= 16'b1111111111110000;
        weights1[3359] <= 16'b1111111111011111;
        weights1[3360] <= 16'b1111111111111111;
        weights1[3361] <= 16'b1111111111111011;
        weights1[3362] <= 16'b1111111111111110;
        weights1[3363] <= 16'b1111111111111001;
        weights1[3364] <= 16'b1111111111110111;
        weights1[3365] <= 16'b0000000000010110;
        weights1[3366] <= 16'b1111111111110100;
        weights1[3367] <= 16'b1111111111101000;
        weights1[3368] <= 16'b1111111111100101;
        weights1[3369] <= 16'b1111111111100010;
        weights1[3370] <= 16'b1111111111111111;
        weights1[3371] <= 16'b0000000000001000;
        weights1[3372] <= 16'b1111111111101100;
        weights1[3373] <= 16'b1111111111101110;
        weights1[3374] <= 16'b0000000000000011;
        weights1[3375] <= 16'b0000000000011110;
        weights1[3376] <= 16'b1111111111101111;
        weights1[3377] <= 16'b1111111111111000;
        weights1[3378] <= 16'b1111111111100010;
        weights1[3379] <= 16'b0000000000001111;
        weights1[3380] <= 16'b1111111111100001;
        weights1[3381] <= 16'b1111111111111100;
        weights1[3382] <= 16'b1111111111101111;
        weights1[3383] <= 16'b1111111111101011;
        weights1[3384] <= 16'b1111111111100100;
        weights1[3385] <= 16'b1111111111100101;
        weights1[3386] <= 16'b1111111111101000;
        weights1[3387] <= 16'b1111111111100001;
        weights1[3388] <= 16'b0000000000000001;
        weights1[3389] <= 16'b1111111111111100;
        weights1[3390] <= 16'b1111111111110111;
        weights1[3391] <= 16'b1111111111110001;
        weights1[3392] <= 16'b1111111111010111;
        weights1[3393] <= 16'b1111111111101100;
        weights1[3394] <= 16'b1111111111010101;
        weights1[3395] <= 16'b0000000000000000;
        weights1[3396] <= 16'b1111111111010001;
        weights1[3397] <= 16'b1111111111110000;
        weights1[3398] <= 16'b1111111111010110;
        weights1[3399] <= 16'b1111111111101101;
        weights1[3400] <= 16'b1111111111001110;
        weights1[3401] <= 16'b1111111111010100;
        weights1[3402] <= 16'b1111111111100010;
        weights1[3403] <= 16'b1111111111100111;
        weights1[3404] <= 16'b1111111111101110;
        weights1[3405] <= 16'b1111111111111111;
        weights1[3406] <= 16'b1111111111110111;
        weights1[3407] <= 16'b1111111111110111;
        weights1[3408] <= 16'b1111111111100001;
        weights1[3409] <= 16'b1111111111111011;
        weights1[3410] <= 16'b0000000000000000;
        weights1[3411] <= 16'b1111111111101110;
        weights1[3412] <= 16'b1111111111100110;
        weights1[3413] <= 16'b1111111111101101;
        weights1[3414] <= 16'b1111111111100100;
        weights1[3415] <= 16'b1111111111011011;
        weights1[3416] <= 16'b1111111111111011;
        weights1[3417] <= 16'b1111111111110001;
        weights1[3418] <= 16'b1111111111101101;
        weights1[3419] <= 16'b1111111111001111;
        weights1[3420] <= 16'b1111111111011011;
        weights1[3421] <= 16'b1111111111001000;
        weights1[3422] <= 16'b1111111111011011;
        weights1[3423] <= 16'b1111111111100100;
        weights1[3424] <= 16'b1111111110111100;
        weights1[3425] <= 16'b1111111111010110;
        weights1[3426] <= 16'b1111111111000000;
        weights1[3427] <= 16'b1111111111001001;
        weights1[3428] <= 16'b1111111111011111;
        weights1[3429] <= 16'b1111111111011001;
        weights1[3430] <= 16'b1111111111011001;
        weights1[3431] <= 16'b1111111111011000;
        weights1[3432] <= 16'b1111111111001110;
        weights1[3433] <= 16'b1111111111110011;
        weights1[3434] <= 16'b1111111111101001;
        weights1[3435] <= 16'b1111111111010101;
        weights1[3436] <= 16'b1111111111011010;
        weights1[3437] <= 16'b1111111111110000;
        weights1[3438] <= 16'b1111111111100110;
        weights1[3439] <= 16'b1111111111010011;
        weights1[3440] <= 16'b1111111111100111;
        weights1[3441] <= 16'b1111111111011111;
        weights1[3442] <= 16'b1111111111100001;
        weights1[3443] <= 16'b1111111111011101;
        weights1[3444] <= 16'b1111111111111100;
        weights1[3445] <= 16'b1111111111101000;
        weights1[3446] <= 16'b1111111111011100;
        weights1[3447] <= 16'b1111111111010001;
        weights1[3448] <= 16'b1111111111100010;
        weights1[3449] <= 16'b1111111111001011;
        weights1[3450] <= 16'b1111111111010011;
        weights1[3451] <= 16'b1111111111001101;
        weights1[3452] <= 16'b1111111111000100;
        weights1[3453] <= 16'b1111111111010100;
        weights1[3454] <= 16'b1111111111000010;
        weights1[3455] <= 16'b1111111111001010;
        weights1[3456] <= 16'b1111111111010000;
        weights1[3457] <= 16'b1111111111010000;
        weights1[3458] <= 16'b1111111111011000;
        weights1[3459] <= 16'b1111111111000010;
        weights1[3460] <= 16'b1111111111011010;
        weights1[3461] <= 16'b1111111111001100;
        weights1[3462] <= 16'b1111111111010100;
        weights1[3463] <= 16'b1111111111100010;
        weights1[3464] <= 16'b1111111111101111;
        weights1[3465] <= 16'b1111111111001101;
        weights1[3466] <= 16'b1111111111010111;
        weights1[3467] <= 16'b1111111111011001;
        weights1[3468] <= 16'b1111111111100100;
        weights1[3469] <= 16'b1111111111011100;
        weights1[3470] <= 16'b1111111111100010;
        weights1[3471] <= 16'b1111111111011001;
        weights1[3472] <= 16'b1111111111111011;
        weights1[3473] <= 16'b1111111111100110;
        weights1[3474] <= 16'b1111111111011011;
        weights1[3475] <= 16'b1111111111100110;
        weights1[3476] <= 16'b1111111111011001;
        weights1[3477] <= 16'b1111111111010001;
        weights1[3478] <= 16'b1111111111100100;
        weights1[3479] <= 16'b1111111110111011;
        weights1[3480] <= 16'b1111111111001101;
        weights1[3481] <= 16'b1111111110110111;
        weights1[3482] <= 16'b1111111110101011;
        weights1[3483] <= 16'b1111111111010001;
        weights1[3484] <= 16'b1111111110101111;
        weights1[3485] <= 16'b1111111111001001;
        weights1[3486] <= 16'b1111111111000100;
        weights1[3487] <= 16'b1111111111000111;
        weights1[3488] <= 16'b1111111110110100;
        weights1[3489] <= 16'b1111111111010101;
        weights1[3490] <= 16'b1111111111010100;
        weights1[3491] <= 16'b1111111111011110;
        weights1[3492] <= 16'b1111111111101001;
        weights1[3493] <= 16'b1111111111011011;
        weights1[3494] <= 16'b1111111111001001;
        weights1[3495] <= 16'b1111111111010110;
        weights1[3496] <= 16'b1111111111011011;
        weights1[3497] <= 16'b1111111111011111;
        weights1[3498] <= 16'b1111111111100011;
        weights1[3499] <= 16'b1111111111100001;
        weights1[3500] <= 16'b1111111111111101;
        weights1[3501] <= 16'b1111111111101101;
        weights1[3502] <= 16'b1111111111011111;
        weights1[3503] <= 16'b1111111111101011;
        weights1[3504] <= 16'b1111111111001111;
        weights1[3505] <= 16'b1111111111010111;
        weights1[3506] <= 16'b1111111111010001;
        weights1[3507] <= 16'b1111111111000101;
        weights1[3508] <= 16'b1111111111100000;
        weights1[3509] <= 16'b1111111111000000;
        weights1[3510] <= 16'b1111111111010000;
        weights1[3511] <= 16'b1111111111010001;
        weights1[3512] <= 16'b1111111111001011;
        weights1[3513] <= 16'b1111111111001110;
        weights1[3514] <= 16'b1111111111000010;
        weights1[3515] <= 16'b1111111111001000;
        weights1[3516] <= 16'b1111111111000110;
        weights1[3517] <= 16'b1111111111010110;
        weights1[3518] <= 16'b1111111110111000;
        weights1[3519] <= 16'b1111111111001101;
        weights1[3520] <= 16'b1111111111011010;
        weights1[3521] <= 16'b1111111111010100;
        weights1[3522] <= 16'b1111111111011001;
        weights1[3523] <= 16'b1111111111100001;
        weights1[3524] <= 16'b1111111111100110;
        weights1[3525] <= 16'b1111111111100101;
        weights1[3526] <= 16'b1111111111100101;
        weights1[3527] <= 16'b1111111111010111;
        weights1[3528] <= 16'b1111111111111110;
        weights1[3529] <= 16'b1111111111111000;
        weights1[3530] <= 16'b1111111111110000;
        weights1[3531] <= 16'b1111111111101010;
        weights1[3532] <= 16'b1111111111100110;
        weights1[3533] <= 16'b1111111111011111;
        weights1[3534] <= 16'b1111111111101011;
        weights1[3535] <= 16'b1111111111100110;
        weights1[3536] <= 16'b1111111111111001;
        weights1[3537] <= 16'b1111111111011101;
        weights1[3538] <= 16'b1111111111101110;
        weights1[3539] <= 16'b1111111111100111;
        weights1[3540] <= 16'b1111111111010000;
        weights1[3541] <= 16'b1111111111100011;
        weights1[3542] <= 16'b1111111111000001;
        weights1[3543] <= 16'b1111111111001000;
        weights1[3544] <= 16'b1111111111001001;
        weights1[3545] <= 16'b1111111110111000;
        weights1[3546] <= 16'b1111111110111011;
        weights1[3547] <= 16'b1111111111001111;
        weights1[3548] <= 16'b1111111111001011;
        weights1[3549] <= 16'b1111111111011001;
        weights1[3550] <= 16'b1111111111010100;
        weights1[3551] <= 16'b1111111111010110;
        weights1[3552] <= 16'b1111111111001010;
        weights1[3553] <= 16'b1111111111010111;
        weights1[3554] <= 16'b1111111111010101;
        weights1[3555] <= 16'b1111111111010110;
        weights1[3556] <= 16'b1111111111111101;
        weights1[3557] <= 16'b0000000000000110;
        weights1[3558] <= 16'b1111111111110010;
        weights1[3559] <= 16'b0000000000000010;
        weights1[3560] <= 16'b1111111111110100;
        weights1[3561] <= 16'b1111111111010001;
        weights1[3562] <= 16'b0000000000001001;
        weights1[3563] <= 16'b1111111111011110;
        weights1[3564] <= 16'b0000000000000111;
        weights1[3565] <= 16'b1111111111111101;
        weights1[3566] <= 16'b1111111111110001;
        weights1[3567] <= 16'b1111111111110110;
        weights1[3568] <= 16'b1111111111110000;
        weights1[3569] <= 16'b1111111111010110;
        weights1[3570] <= 16'b1111111111101110;
        weights1[3571] <= 16'b1111111111100010;
        weights1[3572] <= 16'b1111111111010101;
        weights1[3573] <= 16'b1111111111011011;
        weights1[3574] <= 16'b1111111111000000;
        weights1[3575] <= 16'b1111111110111101;
        weights1[3576] <= 16'b1111111111001010;
        weights1[3577] <= 16'b1111111111001100;
        weights1[3578] <= 16'b1111111111001111;
        weights1[3579] <= 16'b1111111110110001;
        weights1[3580] <= 16'b1111111111001010;
        weights1[3581] <= 16'b1111111111001000;
        weights1[3582] <= 16'b1111111111010110;
        weights1[3583] <= 16'b1111111111011001;
        weights1[3584] <= 16'b0000000000011000;
        weights1[3585] <= 16'b0000000000001110;
        weights1[3586] <= 16'b0000000000010110;
        weights1[3587] <= 16'b0000000000011011;
        weights1[3588] <= 16'b0000000000001101;
        weights1[3589] <= 16'b1111111111111010;
        weights1[3590] <= 16'b0000000000000100;
        weights1[3591] <= 16'b0000000000010001;
        weights1[3592] <= 16'b0000000000001100;
        weights1[3593] <= 16'b0000000000001001;
        weights1[3594] <= 16'b1111111111110101;
        weights1[3595] <= 16'b1111111111001111;
        weights1[3596] <= 16'b0000000000000100;
        weights1[3597] <= 16'b1111111111110110;
        weights1[3598] <= 16'b1111111111101110;
        weights1[3599] <= 16'b1111111111110101;
        weights1[3600] <= 16'b1111111111110111;
        weights1[3601] <= 16'b1111111111100001;
        weights1[3602] <= 16'b1111111111100001;
        weights1[3603] <= 16'b1111111111101000;
        weights1[3604] <= 16'b1111111111011101;
        weights1[3605] <= 16'b1111111110110110;
        weights1[3606] <= 16'b1111111110110010;
        weights1[3607] <= 16'b1111111111000001;
        weights1[3608] <= 16'b1111111110110101;
        weights1[3609] <= 16'b1111111111010000;
        weights1[3610] <= 16'b1111111111011011;
        weights1[3611] <= 16'b1111111111011001;
        weights1[3612] <= 16'b0000000000011111;
        weights1[3613] <= 16'b0000000000010110;
        weights1[3614] <= 16'b0000000000101011;
        weights1[3615] <= 16'b0000000000101000;
        weights1[3616] <= 16'b0000000000010110;
        weights1[3617] <= 16'b0000000000111010;
        weights1[3618] <= 16'b0000000000110100;
        weights1[3619] <= 16'b0000000000110001;
        weights1[3620] <= 16'b0000000000101100;
        weights1[3621] <= 16'b0000000000001111;
        weights1[3622] <= 16'b0000000000011100;
        weights1[3623] <= 16'b1111111111111111;
        weights1[3624] <= 16'b0000000000000101;
        weights1[3625] <= 16'b0000000000001010;
        weights1[3626] <= 16'b1111111111111110;
        weights1[3627] <= 16'b0000000000001101;
        weights1[3628] <= 16'b1111111111111010;
        weights1[3629] <= 16'b1111111111110010;
        weights1[3630] <= 16'b1111111111100100;
        weights1[3631] <= 16'b0000000000000010;
        weights1[3632] <= 16'b1111111111111000;
        weights1[3633] <= 16'b1111111111101110;
        weights1[3634] <= 16'b1111111111110110;
        weights1[3635] <= 16'b1111111111101100;
        weights1[3636] <= 16'b1111111111110000;
        weights1[3637] <= 16'b1111111111110011;
        weights1[3638] <= 16'b1111111111100101;
        weights1[3639] <= 16'b1111111111110011;
        weights1[3640] <= 16'b0000000000011110;
        weights1[3641] <= 16'b0000000000101000;
        weights1[3642] <= 16'b0000000000101010;
        weights1[3643] <= 16'b0000000000100000;
        weights1[3644] <= 16'b0000000000111111;
        weights1[3645] <= 16'b0000000001000101;
        weights1[3646] <= 16'b0000000000101111;
        weights1[3647] <= 16'b0000000001001011;
        weights1[3648] <= 16'b0000000000110101;
        weights1[3649] <= 16'b0000000000110111;
        weights1[3650] <= 16'b0000000000011001;
        weights1[3651] <= 16'b0000000000110011;
        weights1[3652] <= 16'b0000000001001111;
        weights1[3653] <= 16'b0000000000011001;
        weights1[3654] <= 16'b0000000000100011;
        weights1[3655] <= 16'b0000000000010111;
        weights1[3656] <= 16'b0000000001000001;
        weights1[3657] <= 16'b0000000000010101;
        weights1[3658] <= 16'b0000000000011100;
        weights1[3659] <= 16'b0000000000101000;
        weights1[3660] <= 16'b0000000000011001;
        weights1[3661] <= 16'b0000000000001010;
        weights1[3662] <= 16'b0000000000100000;
        weights1[3663] <= 16'b0000000000101100;
        weights1[3664] <= 16'b0000000000100001;
        weights1[3665] <= 16'b0000000000000110;
        weights1[3666] <= 16'b1111111111110011;
        weights1[3667] <= 16'b0000000000001111;
        weights1[3668] <= 16'b0000000000101000;
        weights1[3669] <= 16'b0000000000101100;
        weights1[3670] <= 16'b0000000000011101;
        weights1[3671] <= 16'b0000000000100000;
        weights1[3672] <= 16'b0000000000100011;
        weights1[3673] <= 16'b0000000000110110;
        weights1[3674] <= 16'b0000000000111011;
        weights1[3675] <= 16'b0000000000111100;
        weights1[3676] <= 16'b0000000001001000;
        weights1[3677] <= 16'b0000000001000101;
        weights1[3678] <= 16'b0000000001000110;
        weights1[3679] <= 16'b0000000001011010;
        weights1[3680] <= 16'b0000000001001111;
        weights1[3681] <= 16'b0000000001001000;
        weights1[3682] <= 16'b0000000000111111;
        weights1[3683] <= 16'b0000000001001000;
        weights1[3684] <= 16'b0000000000101110;
        weights1[3685] <= 16'b0000000000100001;
        weights1[3686] <= 16'b0000000000110100;
        weights1[3687] <= 16'b0000000000101011;
        weights1[3688] <= 16'b0000000000011101;
        weights1[3689] <= 16'b0000000000011111;
        weights1[3690] <= 16'b0000000000100110;
        weights1[3691] <= 16'b0000000000110001;
        weights1[3692] <= 16'b0000000000110100;
        weights1[3693] <= 16'b0000000000011110;
        weights1[3694] <= 16'b0000000000011010;
        weights1[3695] <= 16'b0000000000100111;
        weights1[3696] <= 16'b0000000000010101;
        weights1[3697] <= 16'b0000000000011111;
        weights1[3698] <= 16'b0000000000011110;
        weights1[3699] <= 16'b0000000000111101;
        weights1[3700] <= 16'b0000000000111010;
        weights1[3701] <= 16'b0000000000101101;
        weights1[3702] <= 16'b0000000000110111;
        weights1[3703] <= 16'b0000000000111001;
        weights1[3704] <= 16'b0000000000101101;
        weights1[3705] <= 16'b0000000000101111;
        weights1[3706] <= 16'b0000000000110110;
        weights1[3707] <= 16'b0000000001001011;
        weights1[3708] <= 16'b0000000001001100;
        weights1[3709] <= 16'b0000000001001100;
        weights1[3710] <= 16'b0000000001011101;
        weights1[3711] <= 16'b0000000000110110;
        weights1[3712] <= 16'b0000000001000011;
        weights1[3713] <= 16'b0000000000110001;
        weights1[3714] <= 16'b0000000001001000;
        weights1[3715] <= 16'b0000000000111010;
        weights1[3716] <= 16'b0000000001000101;
        weights1[3717] <= 16'b0000000000100010;
        weights1[3718] <= 16'b0000000000100111;
        weights1[3719] <= 16'b0000000000110000;
        weights1[3720] <= 16'b0000000000111101;
        weights1[3721] <= 16'b0000000000101011;
        weights1[3722] <= 16'b0000000000110001;
        weights1[3723] <= 16'b0000000000100100;
        weights1[3724] <= 16'b0000000000000111;
        weights1[3725] <= 16'b0000000000010001;
        weights1[3726] <= 16'b0000000000101011;
        weights1[3727] <= 16'b0000000000110010;
        weights1[3728] <= 16'b0000000000100000;
        weights1[3729] <= 16'b0000000000100001;
        weights1[3730] <= 16'b0000000000100110;
        weights1[3731] <= 16'b0000000000100110;
        weights1[3732] <= 16'b0000000000100111;
        weights1[3733] <= 16'b0000000000100000;
        weights1[3734] <= 16'b0000000000101100;
        weights1[3735] <= 16'b0000000000011100;
        weights1[3736] <= 16'b0000000000010011;
        weights1[3737] <= 16'b0000000000100111;
        weights1[3738] <= 16'b0000000000101110;
        weights1[3739] <= 16'b0000000000101001;
        weights1[3740] <= 16'b0000000000111100;
        weights1[3741] <= 16'b0000000001010001;
        weights1[3742] <= 16'b0000000001000111;
        weights1[3743] <= 16'b0000000001001011;
        weights1[3744] <= 16'b0000000000101110;
        weights1[3745] <= 16'b0000000000111011;
        weights1[3746] <= 16'b0000000000110000;
        weights1[3747] <= 16'b0000000001100000;
        weights1[3748] <= 16'b0000000001001110;
        weights1[3749] <= 16'b0000000001000010;
        weights1[3750] <= 16'b0000000000101100;
        weights1[3751] <= 16'b0000000000100001;
        weights1[3752] <= 16'b0000000000001011;
        weights1[3753] <= 16'b0000000000001110;
        weights1[3754] <= 16'b0000000000001110;
        weights1[3755] <= 16'b0000000000010100;
        weights1[3756] <= 16'b0000000000010110;
        weights1[3757] <= 16'b0000000000100111;
        weights1[3758] <= 16'b0000000000010000;
        weights1[3759] <= 16'b0000000000100000;
        weights1[3760] <= 16'b0000000000110000;
        weights1[3761] <= 16'b0000000000010111;
        weights1[3762] <= 16'b1111111111111001;
        weights1[3763] <= 16'b0000000000010101;
        weights1[3764] <= 16'b0000000000010110;
        weights1[3765] <= 16'b0000000000001011;
        weights1[3766] <= 16'b0000000000011001;
        weights1[3767] <= 16'b0000000000100100;
        weights1[3768] <= 16'b0000000000011110;
        weights1[3769] <= 16'b0000000000101101;
        weights1[3770] <= 16'b0000000000111001;
        weights1[3771] <= 16'b0000000001000100;
        weights1[3772] <= 16'b0000000000110011;
        weights1[3773] <= 16'b0000000000111100;
        weights1[3774] <= 16'b0000000001000110;
        weights1[3775] <= 16'b0000000000111011;
        weights1[3776] <= 16'b0000000001000100;
        weights1[3777] <= 16'b0000000000110111;
        weights1[3778] <= 16'b0000000000100111;
        weights1[3779] <= 16'b0000000000011110;
        weights1[3780] <= 16'b0000000000000010;
        weights1[3781] <= 16'b0000000000000101;
        weights1[3782] <= 16'b0000000000001011;
        weights1[3783] <= 16'b0000000000001100;
        weights1[3784] <= 16'b0000000000001000;
        weights1[3785] <= 16'b0000000000011000;
        weights1[3786] <= 16'b0000000000011010;
        weights1[3787] <= 16'b0000000000001100;
        weights1[3788] <= 16'b0000000000100000;
        weights1[3789] <= 16'b0000000000100000;
        weights1[3790] <= 16'b0000000000011011;
        weights1[3791] <= 16'b0000000000100101;
        weights1[3792] <= 16'b0000000000100011;
        weights1[3793] <= 16'b0000000000000110;
        weights1[3794] <= 16'b0000000000001011;
        weights1[3795] <= 16'b0000000000010111;
        weights1[3796] <= 16'b0000000000010111;
        weights1[3797] <= 16'b0000000000000110;
        weights1[3798] <= 16'b0000000000100111;
        weights1[3799] <= 16'b0000000000111100;
        weights1[3800] <= 16'b0000000001000010;
        weights1[3801] <= 16'b0000000000111111;
        weights1[3802] <= 16'b0000000001000010;
        weights1[3803] <= 16'b0000000000100010;
        weights1[3804] <= 16'b0000000000111110;
        weights1[3805] <= 16'b0000000000110011;
        weights1[3806] <= 16'b0000000000011001;
        weights1[3807] <= 16'b0000000000010000;
        weights1[3808] <= 16'b0000000000000011;
        weights1[3809] <= 16'b0000000000000100;
        weights1[3810] <= 16'b0000000000001100;
        weights1[3811] <= 16'b0000000000000101;
        weights1[3812] <= 16'b0000000000000011;
        weights1[3813] <= 16'b0000000000000100;
        weights1[3814] <= 16'b0000000000000011;
        weights1[3815] <= 16'b0000000000000111;
        weights1[3816] <= 16'b0000000000000101;
        weights1[3817] <= 16'b0000000000000010;
        weights1[3818] <= 16'b1111111111110001;
        weights1[3819] <= 16'b1111111111111011;
        weights1[3820] <= 16'b0000000000010011;
        weights1[3821] <= 16'b0000000000100110;
        weights1[3822] <= 16'b0000000000010101;
        weights1[3823] <= 16'b0000000000000111;
        weights1[3824] <= 16'b0000000000011000;
        weights1[3825] <= 16'b1111111111111010;
        weights1[3826] <= 16'b1111111111111100;
        weights1[3827] <= 16'b0000000000000001;
        weights1[3828] <= 16'b0000000000010001;
        weights1[3829] <= 16'b0000000000001000;
        weights1[3830] <= 16'b0000000000100100;
        weights1[3831] <= 16'b0000000000010111;
        weights1[3832] <= 16'b0000000000110011;
        weights1[3833] <= 16'b0000000000110011;
        weights1[3834] <= 16'b0000000000010100;
        weights1[3835] <= 16'b0000000000001001;
        weights1[3836] <= 16'b0000000000000000;
        weights1[3837] <= 16'b0000000000000001;
        weights1[3838] <= 16'b1111111111110110;
        weights1[3839] <= 16'b1111111111101101;
        weights1[3840] <= 16'b1111111111101101;
        weights1[3841] <= 16'b1111111111111100;
        weights1[3842] <= 16'b0000000000000000;
        weights1[3843] <= 16'b1111111111101011;
        weights1[3844] <= 16'b0000000000001000;
        weights1[3845] <= 16'b0000000000000001;
        weights1[3846] <= 16'b0000000000000101;
        weights1[3847] <= 16'b1111111111111111;
        weights1[3848] <= 16'b1111111111101111;
        weights1[3849] <= 16'b1111111111111111;
        weights1[3850] <= 16'b1111111111111101;
        weights1[3851] <= 16'b0000000000000110;
        weights1[3852] <= 16'b0000000000000110;
        weights1[3853] <= 16'b1111111111110110;
        weights1[3854] <= 16'b0000000000000000;
        weights1[3855] <= 16'b1111111111101000;
        weights1[3856] <= 16'b0000000000000100;
        weights1[3857] <= 16'b1111111111110001;
        weights1[3858] <= 16'b0000000000000000;
        weights1[3859] <= 16'b0000000000001111;
        weights1[3860] <= 16'b0000000000100101;
        weights1[3861] <= 16'b0000000000100011;
        weights1[3862] <= 16'b0000000000001001;
        weights1[3863] <= 16'b0000000000000100;
        weights1[3864] <= 16'b1111111111111110;
        weights1[3865] <= 16'b1111111111111111;
        weights1[3866] <= 16'b1111111111110111;
        weights1[3867] <= 16'b1111111111110000;
        weights1[3868] <= 16'b1111111111110011;
        weights1[3869] <= 16'b1111111111110001;
        weights1[3870] <= 16'b1111111111110010;
        weights1[3871] <= 16'b1111111111110011;
        weights1[3872] <= 16'b1111111111110011;
        weights1[3873] <= 16'b1111111111101111;
        weights1[3874] <= 16'b1111111111101011;
        weights1[3875] <= 16'b1111111111101001;
        weights1[3876] <= 16'b0000000000000110;
        weights1[3877] <= 16'b1111111111111011;
        weights1[3878] <= 16'b0000000000010111;
        weights1[3879] <= 16'b0000000000000011;
        weights1[3880] <= 16'b1111111111111010;
        weights1[3881] <= 16'b1111111111111010;
        weights1[3882] <= 16'b1111111111111001;
        weights1[3883] <= 16'b1111111111111001;
        weights1[3884] <= 16'b0000000000001110;
        weights1[3885] <= 16'b1111111111101110;
        weights1[3886] <= 16'b0000000000001001;
        weights1[3887] <= 16'b0000000000000110;
        weights1[3888] <= 16'b0000000000001001;
        weights1[3889] <= 16'b0000000000010000;
        weights1[3890] <= 16'b0000000000000001;
        weights1[3891] <= 16'b0000000000000000;
        weights1[3892] <= 16'b0000000000000001;
        weights1[3893] <= 16'b1111111111111100;
        weights1[3894] <= 16'b1111111111111100;
        weights1[3895] <= 16'b1111111111110011;
        weights1[3896] <= 16'b1111111111111010;
        weights1[3897] <= 16'b1111111111101111;
        weights1[3898] <= 16'b1111111111101001;
        weights1[3899] <= 16'b1111111111101001;
        weights1[3900] <= 16'b1111111111100110;
        weights1[3901] <= 16'b1111111111100011;
        weights1[3902] <= 16'b1111111111101111;
        weights1[3903] <= 16'b1111111111101101;
        weights1[3904] <= 16'b1111111111110001;
        weights1[3905] <= 16'b1111111111111000;
        weights1[3906] <= 16'b1111111111110001;
        weights1[3907] <= 16'b1111111111100101;
        weights1[3908] <= 16'b1111111111101001;
        weights1[3909] <= 16'b1111111111111111;
        weights1[3910] <= 16'b0000000000000101;
        weights1[3911] <= 16'b0000000000001101;
        weights1[3912] <= 16'b1111111111110101;
        weights1[3913] <= 16'b0000000000000110;
        weights1[3914] <= 16'b0000000000000011;
        weights1[3915] <= 16'b0000000000000100;
        weights1[3916] <= 16'b1111111111111101;
        weights1[3917] <= 16'b1111111111111111;
        weights1[3918] <= 16'b1111111111111011;
        weights1[3919] <= 16'b0000000000000001;
        weights1[3920] <= 16'b0000000000000001;
        weights1[3921] <= 16'b0000000000000001;
        weights1[3922] <= 16'b0000000000000000;
        weights1[3923] <= 16'b0000000000000101;
        weights1[3924] <= 16'b0000000000001001;
        weights1[3925] <= 16'b0000000000001101;
        weights1[3926] <= 16'b0000000000000110;
        weights1[3927] <= 16'b0000000000010110;
        weights1[3928] <= 16'b0000000000100101;
        weights1[3929] <= 16'b0000000000001100;
        weights1[3930] <= 16'b0000000000000011;
        weights1[3931] <= 16'b1111111111110111;
        weights1[3932] <= 16'b1111111111101110;
        weights1[3933] <= 16'b1111111111010011;
        weights1[3934] <= 16'b1111111111011110;
        weights1[3935] <= 16'b1111111111011011;
        weights1[3936] <= 16'b1111111111011000;
        weights1[3937] <= 16'b1111111111100011;
        weights1[3938] <= 16'b1111111111101010;
        weights1[3939] <= 16'b1111111111110010;
        weights1[3940] <= 16'b1111111111111001;
        weights1[3941] <= 16'b1111111111111010;
        weights1[3942] <= 16'b1111111111111011;
        weights1[3943] <= 16'b0000000000000000;
        weights1[3944] <= 16'b0000000000000000;
        weights1[3945] <= 16'b0000000000000000;
        weights1[3946] <= 16'b0000000000000000;
        weights1[3947] <= 16'b0000000000000000;
        weights1[3948] <= 16'b0000000000000010;
        weights1[3949] <= 16'b0000000000000100;
        weights1[3950] <= 16'b0000000000001010;
        weights1[3951] <= 16'b0000000000000101;
        weights1[3952] <= 16'b0000000000010010;
        weights1[3953] <= 16'b0000000000011111;
        weights1[3954] <= 16'b0000000000100100;
        weights1[3955] <= 16'b0000000000100001;
        weights1[3956] <= 16'b0000000000100001;
        weights1[3957] <= 16'b0000000000000111;
        weights1[3958] <= 16'b0000000000000101;
        weights1[3959] <= 16'b1111111111111101;
        weights1[3960] <= 16'b1111111111110001;
        weights1[3961] <= 16'b1111111111101000;
        weights1[3962] <= 16'b1111111111100111;
        weights1[3963] <= 16'b1111111111100010;
        weights1[3964] <= 16'b1111111111011100;
        weights1[3965] <= 16'b1111111111011001;
        weights1[3966] <= 16'b1111111111011011;
        weights1[3967] <= 16'b1111111111100001;
        weights1[3968] <= 16'b1111111111110011;
        weights1[3969] <= 16'b1111111111110101;
        weights1[3970] <= 16'b1111111111111011;
        weights1[3971] <= 16'b1111111111111100;
        weights1[3972] <= 16'b1111111111111111;
        weights1[3973] <= 16'b0000000000000000;
        weights1[3974] <= 16'b0000000000000000;
        weights1[3975] <= 16'b0000000000000000;
        weights1[3976] <= 16'b0000000000000110;
        weights1[3977] <= 16'b0000000000001001;
        weights1[3978] <= 16'b0000000000001011;
        weights1[3979] <= 16'b0000000000010100;
        weights1[3980] <= 16'b0000000000010100;
        weights1[3981] <= 16'b0000000000100100;
        weights1[3982] <= 16'b0000000000100000;
        weights1[3983] <= 16'b0000000000010110;
        weights1[3984] <= 16'b0000000000010011;
        weights1[3985] <= 16'b0000000000001000;
        weights1[3986] <= 16'b0000000000001100;
        weights1[3987] <= 16'b0000000000001010;
        weights1[3988] <= 16'b0000000000000110;
        weights1[3989] <= 16'b1111111111101001;
        weights1[3990] <= 16'b1111111111100010;
        weights1[3991] <= 16'b1111111111100000;
        weights1[3992] <= 16'b1111111111101000;
        weights1[3993] <= 16'b1111111111001111;
        weights1[3994] <= 16'b1111111111000100;
        weights1[3995] <= 16'b1111111111010000;
        weights1[3996] <= 16'b1111111111011111;
        weights1[3997] <= 16'b1111111111110100;
        weights1[3998] <= 16'b1111111111111011;
        weights1[3999] <= 16'b1111111111111101;
        weights1[4000] <= 16'b0000000000000000;
        weights1[4001] <= 16'b0000000000000001;
        weights1[4002] <= 16'b0000000000000000;
        weights1[4003] <= 16'b0000000000000000;
        weights1[4004] <= 16'b0000000000001100;
        weights1[4005] <= 16'b0000000000011000;
        weights1[4006] <= 16'b0000000000011000;
        weights1[4007] <= 16'b0000000000001111;
        weights1[4008] <= 16'b0000000000100010;
        weights1[4009] <= 16'b0000000000011010;
        weights1[4010] <= 16'b0000000000100111;
        weights1[4011] <= 16'b0000000000100001;
        weights1[4012] <= 16'b0000000000010101;
        weights1[4013] <= 16'b0000000000000011;
        weights1[4014] <= 16'b0000000000010110;
        weights1[4015] <= 16'b1111111111111100;
        weights1[4016] <= 16'b1111111111100110;
        weights1[4017] <= 16'b1111111111100101;
        weights1[4018] <= 16'b1111111111100110;
        weights1[4019] <= 16'b1111111110111110;
        weights1[4020] <= 16'b1111111111100100;
        weights1[4021] <= 16'b1111111111010010;
        weights1[4022] <= 16'b1111111110110010;
        weights1[4023] <= 16'b1111111111001000;
        weights1[4024] <= 16'b1111111111100001;
        weights1[4025] <= 16'b1111111111110000;
        weights1[4026] <= 16'b1111111111110111;
        weights1[4027] <= 16'b1111111111111001;
        weights1[4028] <= 16'b0000000000000000;
        weights1[4029] <= 16'b0000000000000000;
        weights1[4030] <= 16'b0000000000000000;
        weights1[4031] <= 16'b0000000000000000;
        weights1[4032] <= 16'b0000000000001100;
        weights1[4033] <= 16'b0000000000011100;
        weights1[4034] <= 16'b0000000000010011;
        weights1[4035] <= 16'b0000000000010011;
        weights1[4036] <= 16'b0000000000010001;
        weights1[4037] <= 16'b0000000000010100;
        weights1[4038] <= 16'b0000000000010101;
        weights1[4039] <= 16'b0000000000011000;
        weights1[4040] <= 16'b0000000000011100;
        weights1[4041] <= 16'b0000000000001100;
        weights1[4042] <= 16'b0000000000010111;
        weights1[4043] <= 16'b0000000000011010;
        weights1[4044] <= 16'b0000000000010110;
        weights1[4045] <= 16'b0000000000011010;
        weights1[4046] <= 16'b0000000000000001;
        weights1[4047] <= 16'b1111111111100100;
        weights1[4048] <= 16'b1111111111000000;
        weights1[4049] <= 16'b1111111110101000;
        weights1[4050] <= 16'b1111111110100111;
        weights1[4051] <= 16'b1111111111000010;
        weights1[4052] <= 16'b1111111111011010;
        weights1[4053] <= 16'b1111111111101101;
        weights1[4054] <= 16'b1111111111110011;
        weights1[4055] <= 16'b1111111111110110;
        weights1[4056] <= 16'b1111111111111110;
        weights1[4057] <= 16'b0000000000000000;
        weights1[4058] <= 16'b0000000000000000;
        weights1[4059] <= 16'b0000000000000000;
        weights1[4060] <= 16'b0000000000001100;
        weights1[4061] <= 16'b0000000000011101;
        weights1[4062] <= 16'b0000000000010110;
        weights1[4063] <= 16'b0000000000011000;
        weights1[4064] <= 16'b0000000000001010;
        weights1[4065] <= 16'b0000000000011110;
        weights1[4066] <= 16'b0000000000001110;
        weights1[4067] <= 16'b0000000000010111;
        weights1[4068] <= 16'b0000000000010111;
        weights1[4069] <= 16'b0000000000000001;
        weights1[4070] <= 16'b0000000000011011;
        weights1[4071] <= 16'b0000000000010011;
        weights1[4072] <= 16'b0000000000001111;
        weights1[4073] <= 16'b0000000000010010;
        weights1[4074] <= 16'b1111111111111001;
        weights1[4075] <= 16'b0000000000000110;
        weights1[4076] <= 16'b1111111111111001;
        weights1[4077] <= 16'b1111111110110101;
        weights1[4078] <= 16'b1111111110101001;
        weights1[4079] <= 16'b1111111110101111;
        weights1[4080] <= 16'b1111111111011000;
        weights1[4081] <= 16'b1111111111110001;
        weights1[4082] <= 16'b1111111111110010;
        weights1[4083] <= 16'b1111111111110100;
        weights1[4084] <= 16'b1111111111111011;
        weights1[4085] <= 16'b1111111111111011;
        weights1[4086] <= 16'b1111111111111100;
        weights1[4087] <= 16'b0000000000000000;
        weights1[4088] <= 16'b0000000000001101;
        weights1[4089] <= 16'b0000000000010101;
        weights1[4090] <= 16'b0000000000011110;
        weights1[4091] <= 16'b0000000000011111;
        weights1[4092] <= 16'b0000000000010100;
        weights1[4093] <= 16'b0000000000011001;
        weights1[4094] <= 16'b0000000000011011;
        weights1[4095] <= 16'b0000000000101110;
        weights1[4096] <= 16'b0000000000010001;
        weights1[4097] <= 16'b0000000000001101;
        weights1[4098] <= 16'b0000000000100010;
        weights1[4099] <= 16'b0000000000100000;
        weights1[4100] <= 16'b0000000000001100;
        weights1[4101] <= 16'b0000000000010010;
        weights1[4102] <= 16'b1111111111110101;
        weights1[4103] <= 16'b0000000000000011;
        weights1[4104] <= 16'b1111111111110000;
        weights1[4105] <= 16'b1111111111000100;
        weights1[4106] <= 16'b1111111101111010;
        weights1[4107] <= 16'b1111111110010100;
        weights1[4108] <= 16'b1111111111011010;
        weights1[4109] <= 16'b1111111111101001;
        weights1[4110] <= 16'b1111111111101100;
        weights1[4111] <= 16'b1111111111110010;
        weights1[4112] <= 16'b1111111111110010;
        weights1[4113] <= 16'b1111111111110111;
        weights1[4114] <= 16'b1111111111111011;
        weights1[4115] <= 16'b0000000000000000;
        weights1[4116] <= 16'b0000000000010101;
        weights1[4117] <= 16'b0000000000100010;
        weights1[4118] <= 16'b0000000000101000;
        weights1[4119] <= 16'b0000000000010000;
        weights1[4120] <= 16'b0000000000001111;
        weights1[4121] <= 16'b1111111111110111;
        weights1[4122] <= 16'b0000000000000101;
        weights1[4123] <= 16'b1111111111101010;
        weights1[4124] <= 16'b1111111111111101;
        weights1[4125] <= 16'b0000000000010000;
        weights1[4126] <= 16'b0000000000010001;
        weights1[4127] <= 16'b0000000000110101;
        weights1[4128] <= 16'b0000000000011101;
        weights1[4129] <= 16'b0000000000000010;
        weights1[4130] <= 16'b0000000000010011;
        weights1[4131] <= 16'b0000000000001011;
        weights1[4132] <= 16'b0000000000001101;
        weights1[4133] <= 16'b1111111110111001;
        weights1[4134] <= 16'b1111111101100010;
        weights1[4135] <= 16'b1111111110010111;
        weights1[4136] <= 16'b1111111111010010;
        weights1[4137] <= 16'b1111111111101011;
        weights1[4138] <= 16'b1111111111101111;
        weights1[4139] <= 16'b1111111111101111;
        weights1[4140] <= 16'b1111111111110100;
        weights1[4141] <= 16'b1111111111110011;
        weights1[4142] <= 16'b1111111111111011;
        weights1[4143] <= 16'b0000000000000000;
        weights1[4144] <= 16'b0000000000011110;
        weights1[4145] <= 16'b0000000000100000;
        weights1[4146] <= 16'b0000000000000010;
        weights1[4147] <= 16'b0000000000001000;
        weights1[4148] <= 16'b0000000000000100;
        weights1[4149] <= 16'b1111111111111000;
        weights1[4150] <= 16'b1111111111111100;
        weights1[4151] <= 16'b0000000000001100;
        weights1[4152] <= 16'b1111111111110100;
        weights1[4153] <= 16'b0000000000000111;
        weights1[4154] <= 16'b0000000000111111;
        weights1[4155] <= 16'b0000000000100100;
        weights1[4156] <= 16'b0000000000101000;
        weights1[4157] <= 16'b0000000000110011;
        weights1[4158] <= 16'b0000000000101110;
        weights1[4159] <= 16'b0000000000001101;
        weights1[4160] <= 16'b1111111111101001;
        weights1[4161] <= 16'b1111111111010011;
        weights1[4162] <= 16'b1111111101110111;
        weights1[4163] <= 16'b1111111110101111;
        weights1[4164] <= 16'b1111111111001010;
        weights1[4165] <= 16'b1111111111011100;
        weights1[4166] <= 16'b1111111111100101;
        weights1[4167] <= 16'b1111111111101000;
        weights1[4168] <= 16'b1111111111101111;
        weights1[4169] <= 16'b1111111111110010;
        weights1[4170] <= 16'b1111111111110110;
        weights1[4171] <= 16'b1111111111111001;
        weights1[4172] <= 16'b0000000000010011;
        weights1[4173] <= 16'b0000000000010000;
        weights1[4174] <= 16'b0000000000010000;
        weights1[4175] <= 16'b0000000000000011;
        weights1[4176] <= 16'b0000000000000110;
        weights1[4177] <= 16'b0000000000001110;
        weights1[4178] <= 16'b1111111111110101;
        weights1[4179] <= 16'b1111111111101010;
        weights1[4180] <= 16'b1111111111101111;
        weights1[4181] <= 16'b0000000000011000;
        weights1[4182] <= 16'b0000000000101100;
        weights1[4183] <= 16'b0000000000011100;
        weights1[4184] <= 16'b0000000000101000;
        weights1[4185] <= 16'b0000000000111111;
        weights1[4186] <= 16'b0000000000101010;
        weights1[4187] <= 16'b0000000000011111;
        weights1[4188] <= 16'b1111111111010101;
        weights1[4189] <= 16'b1111111110110110;
        weights1[4190] <= 16'b1111111101111010;
        weights1[4191] <= 16'b1111111110111011;
        weights1[4192] <= 16'b1111111111000110;
        weights1[4193] <= 16'b1111111111011010;
        weights1[4194] <= 16'b1111111111100001;
        weights1[4195] <= 16'b1111111111011100;
        weights1[4196] <= 16'b1111111111011111;
        weights1[4197] <= 16'b1111111111110001;
        weights1[4198] <= 16'b1111111111110110;
        weights1[4199] <= 16'b1111111111111111;
        weights1[4200] <= 16'b0000000000011010;
        weights1[4201] <= 16'b0000000000100100;
        weights1[4202] <= 16'b0000000000011111;
        weights1[4203] <= 16'b0000000000000010;
        weights1[4204] <= 16'b1111111111111001;
        weights1[4205] <= 16'b1111111111110010;
        weights1[4206] <= 16'b1111111111110110;
        weights1[4207] <= 16'b1111111111110111;
        weights1[4208] <= 16'b1111111111111001;
        weights1[4209] <= 16'b1111111111111001;
        weights1[4210] <= 16'b0000000000101001;
        weights1[4211] <= 16'b0000000000101111;
        weights1[4212] <= 16'b0000000000101111;
        weights1[4213] <= 16'b0000000000110110;
        weights1[4214] <= 16'b0000000000100011;
        weights1[4215] <= 16'b0000000000000001;
        weights1[4216] <= 16'b1111111111101000;
        weights1[4217] <= 16'b1111111110111011;
        weights1[4218] <= 16'b1111111110010101;
        weights1[4219] <= 16'b1111111111000101;
        weights1[4220] <= 16'b1111111111000100;
        weights1[4221] <= 16'b1111111111011101;
        weights1[4222] <= 16'b1111111111100111;
        weights1[4223] <= 16'b1111111111011100;
        weights1[4224] <= 16'b1111111111100001;
        weights1[4225] <= 16'b1111111111110100;
        weights1[4226] <= 16'b1111111111111001;
        weights1[4227] <= 16'b1111111111110111;
        weights1[4228] <= 16'b0000000000011011;
        weights1[4229] <= 16'b0000000000010100;
        weights1[4230] <= 16'b0000000000001000;
        weights1[4231] <= 16'b0000000000001000;
        weights1[4232] <= 16'b1111111111111101;
        weights1[4233] <= 16'b0000000000000001;
        weights1[4234] <= 16'b1111111111100101;
        weights1[4235] <= 16'b1111111111110010;
        weights1[4236] <= 16'b1111111111100110;
        weights1[4237] <= 16'b1111111111101010;
        weights1[4238] <= 16'b0000000000000010;
        weights1[4239] <= 16'b0000000000100100;
        weights1[4240] <= 16'b0000000000011101;
        weights1[4241] <= 16'b0000000000111101;
        weights1[4242] <= 16'b0000000000110100;
        weights1[4243] <= 16'b1111111111111100;
        weights1[4244] <= 16'b1111111111011100;
        weights1[4245] <= 16'b1111111111001110;
        weights1[4246] <= 16'b1111111110101101;
        weights1[4247] <= 16'b1111111111000111;
        weights1[4248] <= 16'b1111111111010010;
        weights1[4249] <= 16'b1111111111001100;
        weights1[4250] <= 16'b1111111111100011;
        weights1[4251] <= 16'b1111111111101011;
        weights1[4252] <= 16'b1111111111101001;
        weights1[4253] <= 16'b1111111111111100;
        weights1[4254] <= 16'b1111111111101110;
        weights1[4255] <= 16'b1111111111110110;
        weights1[4256] <= 16'b0000000000011100;
        weights1[4257] <= 16'b0000000000010001;
        weights1[4258] <= 16'b1111111111111110;
        weights1[4259] <= 16'b1111111111111010;
        weights1[4260] <= 16'b1111111111110110;
        weights1[4261] <= 16'b1111111111110000;
        weights1[4262] <= 16'b1111111111101101;
        weights1[4263] <= 16'b1111111111011011;
        weights1[4264] <= 16'b1111111111100000;
        weights1[4265] <= 16'b1111111111110100;
        weights1[4266] <= 16'b1111111111111011;
        weights1[4267] <= 16'b0000000000010100;
        weights1[4268] <= 16'b0000000000100010;
        weights1[4269] <= 16'b0000000000101001;
        weights1[4270] <= 16'b0000000000010110;
        weights1[4271] <= 16'b0000000000000000;
        weights1[4272] <= 16'b1111111111001001;
        weights1[4273] <= 16'b1111111111011110;
        weights1[4274] <= 16'b1111111111100001;
        weights1[4275] <= 16'b1111111111110001;
        weights1[4276] <= 16'b1111111111110101;
        weights1[4277] <= 16'b1111111111100001;
        weights1[4278] <= 16'b1111111111100001;
        weights1[4279] <= 16'b1111111111100001;
        weights1[4280] <= 16'b1111111111101101;
        weights1[4281] <= 16'b1111111111110101;
        weights1[4282] <= 16'b1111111111101110;
        weights1[4283] <= 16'b1111111111110101;
        weights1[4284] <= 16'b0000000000001110;
        weights1[4285] <= 16'b0000000000000000;
        weights1[4286] <= 16'b0000000000000111;
        weights1[4287] <= 16'b1111111111111001;
        weights1[4288] <= 16'b1111111111110101;
        weights1[4289] <= 16'b1111111111101110;
        weights1[4290] <= 16'b1111111111111001;
        weights1[4291] <= 16'b1111111111011011;
        weights1[4292] <= 16'b1111111111101111;
        weights1[4293] <= 16'b1111111111110111;
        weights1[4294] <= 16'b0000000000000011;
        weights1[4295] <= 16'b0000000000101101;
        weights1[4296] <= 16'b0000000000100111;
        weights1[4297] <= 16'b0000000000010000;
        weights1[4298] <= 16'b0000000000010000;
        weights1[4299] <= 16'b1111111111110011;
        weights1[4300] <= 16'b1111111111011010;
        weights1[4301] <= 16'b1111111111111010;
        weights1[4302] <= 16'b1111111111010001;
        weights1[4303] <= 16'b1111111111101110;
        weights1[4304] <= 16'b1111111111010001;
        weights1[4305] <= 16'b1111111111101110;
        weights1[4306] <= 16'b1111111111100100;
        weights1[4307] <= 16'b1111111111111011;
        weights1[4308] <= 16'b1111111111101010;
        weights1[4309] <= 16'b1111111111101001;
        weights1[4310] <= 16'b1111111111101101;
        weights1[4311] <= 16'b1111111111111100;
        weights1[4312] <= 16'b0000000000001010;
        weights1[4313] <= 16'b1111111111111000;
        weights1[4314] <= 16'b1111111111110101;
        weights1[4315] <= 16'b1111111111110000;
        weights1[4316] <= 16'b1111111111101000;
        weights1[4317] <= 16'b1111111111101011;
        weights1[4318] <= 16'b1111111111100100;
        weights1[4319] <= 16'b1111111111011101;
        weights1[4320] <= 16'b1111111111101101;
        weights1[4321] <= 16'b0000000000000011;
        weights1[4322] <= 16'b1111111111111100;
        weights1[4323] <= 16'b0000000000001001;
        weights1[4324] <= 16'b0000000000011111;
        weights1[4325] <= 16'b0000000000001011;
        weights1[4326] <= 16'b0000000000000110;
        weights1[4327] <= 16'b1111111111110100;
        weights1[4328] <= 16'b1111111111101000;
        weights1[4329] <= 16'b1111111111100101;
        weights1[4330] <= 16'b1111111111011010;
        weights1[4331] <= 16'b1111111111111101;
        weights1[4332] <= 16'b1111111111100011;
        weights1[4333] <= 16'b1111111111110010;
        weights1[4334] <= 16'b1111111111100101;
        weights1[4335] <= 16'b1111111111111010;
        weights1[4336] <= 16'b1111111111111100;
        weights1[4337] <= 16'b1111111111110010;
        weights1[4338] <= 16'b1111111111101101;
        weights1[4339] <= 16'b1111111111110110;
        weights1[4340] <= 16'b0000000000001001;
        weights1[4341] <= 16'b1111111111110001;
        weights1[4342] <= 16'b0000000000000101;
        weights1[4343] <= 16'b1111111111110110;
        weights1[4344] <= 16'b1111111111110111;
        weights1[4345] <= 16'b1111111111100111;
        weights1[4346] <= 16'b1111111111110110;
        weights1[4347] <= 16'b1111111111111000;
        weights1[4348] <= 16'b1111111111111010;
        weights1[4349] <= 16'b1111111111111111;
        weights1[4350] <= 16'b1111111111111010;
        weights1[4351] <= 16'b0000000000001101;
        weights1[4352] <= 16'b1111111111111101;
        weights1[4353] <= 16'b0000000000011001;
        weights1[4354] <= 16'b1111111111110110;
        weights1[4355] <= 16'b1111111111100100;
        weights1[4356] <= 16'b1111111111011011;
        weights1[4357] <= 16'b1111111111101010;
        weights1[4358] <= 16'b1111111111011100;
        weights1[4359] <= 16'b1111111111110111;
        weights1[4360] <= 16'b1111111111110000;
        weights1[4361] <= 16'b1111111111111010;
        weights1[4362] <= 16'b1111111111110111;
        weights1[4363] <= 16'b1111111111100010;
        weights1[4364] <= 16'b0000000000010111;
        weights1[4365] <= 16'b0000000000001011;
        weights1[4366] <= 16'b0000000000000100;
        weights1[4367] <= 16'b1111111111101011;
        weights1[4368] <= 16'b0000000000001100;
        weights1[4369] <= 16'b1111111111111000;
        weights1[4370] <= 16'b1111111111111100;
        weights1[4371] <= 16'b1111111111101100;
        weights1[4372] <= 16'b1111111111101101;
        weights1[4373] <= 16'b1111111111111000;
        weights1[4374] <= 16'b1111111111110010;
        weights1[4375] <= 16'b1111111111111011;
        weights1[4376] <= 16'b0000000000010001;
        weights1[4377] <= 16'b1111111111111000;
        weights1[4378] <= 16'b1111111111111110;
        weights1[4379] <= 16'b0000000000000011;
        weights1[4380] <= 16'b0000000000000110;
        weights1[4381] <= 16'b0000000000000000;
        weights1[4382] <= 16'b0000000000001010;
        weights1[4383] <= 16'b1111111111100010;
        weights1[4384] <= 16'b1111111111110111;
        weights1[4385] <= 16'b1111111111011010;
        weights1[4386] <= 16'b1111111111100011;
        weights1[4387] <= 16'b0000000000001100;
        weights1[4388] <= 16'b1111111111111110;
        weights1[4389] <= 16'b0000000000010010;
        weights1[4390] <= 16'b0000000000010000;
        weights1[4391] <= 16'b1111111111111100;
        weights1[4392] <= 16'b0000000000001000;
        weights1[4393] <= 16'b0000000000001010;
        weights1[4394] <= 16'b1111111111111111;
        weights1[4395] <= 16'b1111111111111101;
        weights1[4396] <= 16'b0000000000001100;
        weights1[4397] <= 16'b0000000000000001;
        weights1[4398] <= 16'b0000000000000110;
        weights1[4399] <= 16'b0000000000001010;
        weights1[4400] <= 16'b0000000000001010;
        weights1[4401] <= 16'b1111111111110011;
        weights1[4402] <= 16'b1111111111101111;
        weights1[4403] <= 16'b0000000000001010;
        weights1[4404] <= 16'b1111111111110100;
        weights1[4405] <= 16'b0000000000000010;
        weights1[4406] <= 16'b1111111111110001;
        weights1[4407] <= 16'b1111111111101010;
        weights1[4408] <= 16'b1111111111110001;
        weights1[4409] <= 16'b1111111111110101;
        weights1[4410] <= 16'b0000000000000001;
        weights1[4411] <= 16'b1111111111101101;
        weights1[4412] <= 16'b1111111111111010;
        weights1[4413] <= 16'b0000000000000110;
        weights1[4414] <= 16'b1111111111111001;
        weights1[4415] <= 16'b0000000000001101;
        weights1[4416] <= 16'b1111111111101000;
        weights1[4417] <= 16'b0000000000010110;
        weights1[4418] <= 16'b0000000000011110;
        weights1[4419] <= 16'b0000000000010100;
        weights1[4420] <= 16'b1111111111101110;
        weights1[4421] <= 16'b0000000000000010;
        weights1[4422] <= 16'b1111111111110010;
        weights1[4423] <= 16'b1111111111110011;
        weights1[4424] <= 16'b0000000000001011;
        weights1[4425] <= 16'b0000000000001001;
        weights1[4426] <= 16'b0000000000001111;
        weights1[4427] <= 16'b0000000000000010;
        weights1[4428] <= 16'b1111111111111100;
        weights1[4429] <= 16'b0000000000010001;
        weights1[4430] <= 16'b0000000000001100;
        weights1[4431] <= 16'b1111111111110010;
        weights1[4432] <= 16'b1111111111111110;
        weights1[4433] <= 16'b0000000000000110;
        weights1[4434] <= 16'b1111111111111011;
        weights1[4435] <= 16'b1111111111110110;
        weights1[4436] <= 16'b1111111111110000;
        weights1[4437] <= 16'b0000000000000101;
        weights1[4438] <= 16'b0000000000010101;
        weights1[4439] <= 16'b0000000000001011;
        weights1[4440] <= 16'b1111111111110000;
        weights1[4441] <= 16'b1111111111110100;
        weights1[4442] <= 16'b1111111111111010;
        weights1[4443] <= 16'b1111111111110101;
        weights1[4444] <= 16'b0000000000000001;
        weights1[4445] <= 16'b0000000000001111;
        weights1[4446] <= 16'b0000000000100111;
        weights1[4447] <= 16'b0000000000100011;
        weights1[4448] <= 16'b0000000000000011;
        weights1[4449] <= 16'b1111111111101101;
        weights1[4450] <= 16'b1111111111110100;
        weights1[4451] <= 16'b1111111111111010;
        weights1[4452] <= 16'b0000000000001011;
        weights1[4453] <= 16'b0000000000010001;
        weights1[4454] <= 16'b0000000000100010;
        weights1[4455] <= 16'b0000000000001000;
        weights1[4456] <= 16'b0000000000001101;
        weights1[4457] <= 16'b0000000000000100;
        weights1[4458] <= 16'b1111111111111000;
        weights1[4459] <= 16'b1111111111101010;
        weights1[4460] <= 16'b1111111111111000;
        weights1[4461] <= 16'b1111111111100101;
        weights1[4462] <= 16'b0000000000000100;
        weights1[4463] <= 16'b1111111111101000;
        weights1[4464] <= 16'b1111111111101010;
        weights1[4465] <= 16'b1111111111111110;
        weights1[4466] <= 16'b1111111111101101;
        weights1[4467] <= 16'b0000000000001101;
        weights1[4468] <= 16'b1111111111110011;
        weights1[4469] <= 16'b1111111111101110;
        weights1[4470] <= 16'b0000000000000011;
        weights1[4471] <= 16'b0000000000000001;
        weights1[4472] <= 16'b1111111111101110;
        weights1[4473] <= 16'b1111111111110101;
        weights1[4474] <= 16'b0000000000000010;
        weights1[4475] <= 16'b0000000000000011;
        weights1[4476] <= 16'b1111111111111001;
        weights1[4477] <= 16'b1111111111111000;
        weights1[4478] <= 16'b1111111111110100;
        weights1[4479] <= 16'b1111111111110101;
        weights1[4480] <= 16'b0000000000010010;
        weights1[4481] <= 16'b0000000000010110;
        weights1[4482] <= 16'b0000000000010011;
        weights1[4483] <= 16'b0000000000001011;
        weights1[4484] <= 16'b0000000000000110;
        weights1[4485] <= 16'b0000000000000110;
        weights1[4486] <= 16'b1111111111110010;
        weights1[4487] <= 16'b0000000000000101;
        weights1[4488] <= 16'b0000000000000001;
        weights1[4489] <= 16'b0000000000000001;
        weights1[4490] <= 16'b0000000000000001;
        weights1[4491] <= 16'b1111111111110100;
        weights1[4492] <= 16'b1111111111110100;
        weights1[4493] <= 16'b1111111111111010;
        weights1[4494] <= 16'b0000000000001001;
        weights1[4495] <= 16'b0000000000000100;
        weights1[4496] <= 16'b1111111111111010;
        weights1[4497] <= 16'b0000000000001011;
        weights1[4498] <= 16'b1111111111100011;
        weights1[4499] <= 16'b1111111111101011;
        weights1[4500] <= 16'b1111111111111100;
        weights1[4501] <= 16'b1111111111111001;
        weights1[4502] <= 16'b0000000000001101;
        weights1[4503] <= 16'b1111111111111110;
        weights1[4504] <= 16'b1111111111110101;
        weights1[4505] <= 16'b0000000000000110;
        weights1[4506] <= 16'b1111111111110100;
        weights1[4507] <= 16'b1111111111111000;
        weights1[4508] <= 16'b0000000000010100;
        weights1[4509] <= 16'b0000000000010000;
        weights1[4510] <= 16'b0000000000001001;
        weights1[4511] <= 16'b1111111111111111;
        weights1[4512] <= 16'b1111111111101010;
        weights1[4513] <= 16'b1111111111101001;
        weights1[4514] <= 16'b1111111111110110;
        weights1[4515] <= 16'b0000000000000100;
        weights1[4516] <= 16'b1111111111110101;
        weights1[4517] <= 16'b0000000000000000;
        weights1[4518] <= 16'b0000000000000100;
        weights1[4519] <= 16'b1111111111110100;
        weights1[4520] <= 16'b1111111111101111;
        weights1[4521] <= 16'b1111111111100000;
        weights1[4522] <= 16'b0000000000000010;
        weights1[4523] <= 16'b0000000000010000;
        weights1[4524] <= 16'b1111111111110010;
        weights1[4525] <= 16'b1111111111111110;
        weights1[4526] <= 16'b0000000000000100;
        weights1[4527] <= 16'b1111111111110011;
        weights1[4528] <= 16'b1111111111101010;
        weights1[4529] <= 16'b1111111111011110;
        weights1[4530] <= 16'b1111111111101111;
        weights1[4531] <= 16'b1111111111100110;
        weights1[4532] <= 16'b1111111111110110;
        weights1[4533] <= 16'b1111111111111001;
        weights1[4534] <= 16'b1111111111111000;
        weights1[4535] <= 16'b1111111111111000;
        weights1[4536] <= 16'b0000000000001100;
        weights1[4537] <= 16'b0000000000011001;
        weights1[4538] <= 16'b0000000000000101;
        weights1[4539] <= 16'b0000000000001011;
        weights1[4540] <= 16'b1111111111111111;
        weights1[4541] <= 16'b1111111111110011;
        weights1[4542] <= 16'b1111111111110100;
        weights1[4543] <= 16'b1111111111110110;
        weights1[4544] <= 16'b1111111111111000;
        weights1[4545] <= 16'b0000000000000101;
        weights1[4546] <= 16'b1111111111110100;
        weights1[4547] <= 16'b0000000000001010;
        weights1[4548] <= 16'b0000000000000110;
        weights1[4549] <= 16'b1111111111110111;
        weights1[4550] <= 16'b1111111111101101;
        weights1[4551] <= 16'b1111111111110010;
        weights1[4552] <= 16'b1111111111101010;
        weights1[4553] <= 16'b1111111111110010;
        weights1[4554] <= 16'b0000000000001011;
        weights1[4555] <= 16'b1111111111111000;
        weights1[4556] <= 16'b0000000000011110;
        weights1[4557] <= 16'b1111111111111010;
        weights1[4558] <= 16'b1111111111011100;
        weights1[4559] <= 16'b1111111111111010;
        weights1[4560] <= 16'b0000000000000000;
        weights1[4561] <= 16'b1111111111111001;
        weights1[4562] <= 16'b1111111111110111;
        weights1[4563] <= 16'b1111111111111010;
        weights1[4564] <= 16'b0000000000000101;
        weights1[4565] <= 16'b0000000000001011;
        weights1[4566] <= 16'b0000000000001111;
        weights1[4567] <= 16'b0000000000001001;
        weights1[4568] <= 16'b0000000000001000;
        weights1[4569] <= 16'b0000000000000110;
        weights1[4570] <= 16'b0000000000001010;
        weights1[4571] <= 16'b1111111111110001;
        weights1[4572] <= 16'b1111111111111011;
        weights1[4573] <= 16'b0000000000000110;
        weights1[4574] <= 16'b0000000000010000;
        weights1[4575] <= 16'b0000000000000100;
        weights1[4576] <= 16'b1111111111111001;
        weights1[4577] <= 16'b1111111111111010;
        weights1[4578] <= 16'b1111111111111100;
        weights1[4579] <= 16'b0000000000011100;
        weights1[4580] <= 16'b1111111111110100;
        weights1[4581] <= 16'b0000000000001001;
        weights1[4582] <= 16'b1111111111101000;
        weights1[4583] <= 16'b1111111111111011;
        weights1[4584] <= 16'b1111111111110111;
        weights1[4585] <= 16'b1111111111110011;
        weights1[4586] <= 16'b1111111111111001;
        weights1[4587] <= 16'b1111111111101100;
        weights1[4588] <= 16'b1111111111111111;
        weights1[4589] <= 16'b1111111111111011;
        weights1[4590] <= 16'b0000000000000010;
        weights1[4591] <= 16'b0000000000000000;
        weights1[4592] <= 16'b0000000000000100;
        weights1[4593] <= 16'b0000000000001011;
        weights1[4594] <= 16'b0000000000000100;
        weights1[4595] <= 16'b0000000000000100;
        weights1[4596] <= 16'b1111111111111110;
        weights1[4597] <= 16'b0000000000000010;
        weights1[4598] <= 16'b1111111111111011;
        weights1[4599] <= 16'b0000000000000110;
        weights1[4600] <= 16'b0000000000011001;
        weights1[4601] <= 16'b0000000000000010;
        weights1[4602] <= 16'b1111111111111110;
        weights1[4603] <= 16'b1111111111110101;
        weights1[4604] <= 16'b1111111111100011;
        weights1[4605] <= 16'b0000000000000010;
        weights1[4606] <= 16'b1111111111101011;
        weights1[4607] <= 16'b1111111111110010;
        weights1[4608] <= 16'b1111111111101000;
        weights1[4609] <= 16'b1111111111111101;
        weights1[4610] <= 16'b1111111111100010;
        weights1[4611] <= 16'b1111111111111001;
        weights1[4612] <= 16'b1111111111101111;
        weights1[4613] <= 16'b1111111111111101;
        weights1[4614] <= 16'b1111111111110001;
        weights1[4615] <= 16'b1111111111111110;
        weights1[4616] <= 16'b1111111111111101;
        weights1[4617] <= 16'b1111111111111100;
        weights1[4618] <= 16'b0000000000000100;
        weights1[4619] <= 16'b0000000000000100;
        weights1[4620] <= 16'b1111111111111101;
        weights1[4621] <= 16'b0000000000001110;
        weights1[4622] <= 16'b0000000000010000;
        weights1[4623] <= 16'b0000000000001010;
        weights1[4624] <= 16'b0000000000001000;
        weights1[4625] <= 16'b0000000000001100;
        weights1[4626] <= 16'b0000000000000010;
        weights1[4627] <= 16'b0000000000000110;
        weights1[4628] <= 16'b1111111111111111;
        weights1[4629] <= 16'b1111111111100101;
        weights1[4630] <= 16'b1111111111111111;
        weights1[4631] <= 16'b1111111111101000;
        weights1[4632] <= 16'b1111111111110111;
        weights1[4633] <= 16'b1111111111110101;
        weights1[4634] <= 16'b1111111111111110;
        weights1[4635] <= 16'b1111111111110101;
        weights1[4636] <= 16'b0000000000001111;
        weights1[4637] <= 16'b0000000000010101;
        weights1[4638] <= 16'b0000000000001010;
        weights1[4639] <= 16'b1111111111111110;
        weights1[4640] <= 16'b1111111111101111;
        weights1[4641] <= 16'b1111111111111111;
        weights1[4642] <= 16'b1111111111111000;
        weights1[4643] <= 16'b1111111111111010;
        weights1[4644] <= 16'b1111111111111111;
        weights1[4645] <= 16'b0000000000000001;
        weights1[4646] <= 16'b1111111111111101;
        weights1[4647] <= 16'b0000000000000001;
        weights1[4648] <= 16'b0000000000000001;
        weights1[4649] <= 16'b0000000000000110;
        weights1[4650] <= 16'b0000000000010010;
        weights1[4651] <= 16'b0000000000010001;
        weights1[4652] <= 16'b0000000000000100;
        weights1[4653] <= 16'b0000000000000011;
        weights1[4654] <= 16'b0000000000010110;
        weights1[4655] <= 16'b0000000000001001;
        weights1[4656] <= 16'b0000000000000011;
        weights1[4657] <= 16'b1111111111111101;
        weights1[4658] <= 16'b0000000000011100;
        weights1[4659] <= 16'b1111111111110100;
        weights1[4660] <= 16'b0000000000001100;
        weights1[4661] <= 16'b0000000000001101;
        weights1[4662] <= 16'b1111111111110001;
        weights1[4663] <= 16'b1111111111110001;
        weights1[4664] <= 16'b0000000000000111;
        weights1[4665] <= 16'b0000000000011000;
        weights1[4666] <= 16'b0000000000010011;
        weights1[4667] <= 16'b0000000000010011;
        weights1[4668] <= 16'b0000000000000110;
        weights1[4669] <= 16'b0000000000010011;
        weights1[4670] <= 16'b1111111111111011;
        weights1[4671] <= 16'b1111111111111010;
        weights1[4672] <= 16'b0000000000000000;
        weights1[4673] <= 16'b0000000000000000;
        weights1[4674] <= 16'b1111111111111110;
        weights1[4675] <= 16'b1111111111111111;
        weights1[4676] <= 16'b0000000000000101;
        weights1[4677] <= 16'b0000000000000110;
        weights1[4678] <= 16'b0000000000001100;
        weights1[4679] <= 16'b0000000000010001;
        weights1[4680] <= 16'b0000000000010001;
        weights1[4681] <= 16'b0000000000010011;
        weights1[4682] <= 16'b0000000000001111;
        weights1[4683] <= 16'b0000000000000110;
        weights1[4684] <= 16'b0000000000001011;
        weights1[4685] <= 16'b0000000000000100;
        weights1[4686] <= 16'b0000000000001101;
        weights1[4687] <= 16'b1111111111111111;
        weights1[4688] <= 16'b0000000000001001;
        weights1[4689] <= 16'b0000000000001111;
        weights1[4690] <= 16'b1111111111111100;
        weights1[4691] <= 16'b0000000000010000;
        weights1[4692] <= 16'b0000000000001111;
        weights1[4693] <= 16'b0000000000010011;
        weights1[4694] <= 16'b0000000000010010;
        weights1[4695] <= 16'b0000000000000010;
        weights1[4696] <= 16'b0000000000000110;
        weights1[4697] <= 16'b0000000000000011;
        weights1[4698] <= 16'b1111111111111101;
        weights1[4699] <= 16'b1111111111111011;
        weights1[4700] <= 16'b0000000000000000;
        weights1[4701] <= 16'b0000000000000001;
        weights1[4702] <= 16'b1111111111111111;
        weights1[4703] <= 16'b1111111111111111;
        weights1[4704] <= 16'b0000000000000000;
        weights1[4705] <= 16'b0000000000000000;
        weights1[4706] <= 16'b0000000000000000;
        weights1[4707] <= 16'b0000000000000000;
        weights1[4708] <= 16'b0000000000000000;
        weights1[4709] <= 16'b0000000000000000;
        weights1[4710] <= 16'b0000000000000000;
        weights1[4711] <= 16'b0000000000000000;
        weights1[4712] <= 16'b0000000000000000;
        weights1[4713] <= 16'b0000000000000000;
        weights1[4714] <= 16'b0000000000000000;
        weights1[4715] <= 16'b0000000000000000;
        weights1[4716] <= 16'b0000000000000000;
        weights1[4717] <= 16'b0000000000000000;
        weights1[4718] <= 16'b0000000000000000;
        weights1[4719] <= 16'b0000000000000000;
        weights1[4720] <= 16'b0000000000000000;
        weights1[4721] <= 16'b0000000000000000;
        weights1[4722] <= 16'b0000000000000000;
        weights1[4723] <= 16'b0000000000000000;
        weights1[4724] <= 16'b0000000000000000;
        weights1[4725] <= 16'b0000000000000000;
        weights1[4726] <= 16'b0000000000000000;
        weights1[4727] <= 16'b0000000000000000;
        weights1[4728] <= 16'b0000000000000000;
        weights1[4729] <= 16'b0000000000000000;
        weights1[4730] <= 16'b0000000000000000;
        weights1[4731] <= 16'b0000000000000000;
        weights1[4732] <= 16'b0000000000000000;
        weights1[4733] <= 16'b0000000000000000;
        weights1[4734] <= 16'b0000000000000000;
        weights1[4735] <= 16'b0000000000000000;
        weights1[4736] <= 16'b0000000000000000;
        weights1[4737] <= 16'b0000000000000000;
        weights1[4738] <= 16'b0000000000000000;
        weights1[4739] <= 16'b0000000000000000;
        weights1[4740] <= 16'b0000000000000000;
        weights1[4741] <= 16'b0000000000000000;
        weights1[4742] <= 16'b0000000000000000;
        weights1[4743] <= 16'b0000000000000000;
        weights1[4744] <= 16'b0000000000000000;
        weights1[4745] <= 16'b0000000000000000;
        weights1[4746] <= 16'b0000000000000000;
        weights1[4747] <= 16'b0000000000000000;
        weights1[4748] <= 16'b0000000000000000;
        weights1[4749] <= 16'b0000000000000000;
        weights1[4750] <= 16'b0000000000000000;
        weights1[4751] <= 16'b0000000000000000;
        weights1[4752] <= 16'b0000000000000000;
        weights1[4753] <= 16'b0000000000000000;
        weights1[4754] <= 16'b0000000000000000;
        weights1[4755] <= 16'b0000000000000000;
        weights1[4756] <= 16'b0000000000000000;
        weights1[4757] <= 16'b0000000000000000;
        weights1[4758] <= 16'b0000000000000000;
        weights1[4759] <= 16'b0000000000000000;
        weights1[4760] <= 16'b0000000000000000;
        weights1[4761] <= 16'b0000000000000000;
        weights1[4762] <= 16'b0000000000000000;
        weights1[4763] <= 16'b0000000000000000;
        weights1[4764] <= 16'b0000000000000000;
        weights1[4765] <= 16'b0000000000000000;
        weights1[4766] <= 16'b0000000000000000;
        weights1[4767] <= 16'b0000000000000000;
        weights1[4768] <= 16'b0000000000000000;
        weights1[4769] <= 16'b0000000000000000;
        weights1[4770] <= 16'b0000000000000000;
        weights1[4771] <= 16'b0000000000000000;
        weights1[4772] <= 16'b0000000000000000;
        weights1[4773] <= 16'b0000000000000000;
        weights1[4774] <= 16'b0000000000000000;
        weights1[4775] <= 16'b0000000000000000;
        weights1[4776] <= 16'b0000000000000000;
        weights1[4777] <= 16'b0000000000000000;
        weights1[4778] <= 16'b0000000000000000;
        weights1[4779] <= 16'b0000000000000000;
        weights1[4780] <= 16'b0000000000000000;
        weights1[4781] <= 16'b0000000000000000;
        weights1[4782] <= 16'b0000000000000000;
        weights1[4783] <= 16'b0000000000000000;
        weights1[4784] <= 16'b0000000000000000;
        weights1[4785] <= 16'b0000000000000000;
        weights1[4786] <= 16'b0000000000000000;
        weights1[4787] <= 16'b0000000000000000;
        weights1[4788] <= 16'b0000000000000000;
        weights1[4789] <= 16'b0000000000000000;
        weights1[4790] <= 16'b0000000000000000;
        weights1[4791] <= 16'b0000000000000000;
        weights1[4792] <= 16'b0000000000000000;
        weights1[4793] <= 16'b0000000000000000;
        weights1[4794] <= 16'b0000000000000000;
        weights1[4795] <= 16'b0000000000000000;
        weights1[4796] <= 16'b0000000000000000;
        weights1[4797] <= 16'b0000000000000000;
        weights1[4798] <= 16'b0000000000000000;
        weights1[4799] <= 16'b0000000000000000;
        weights1[4800] <= 16'b0000000000000000;
        weights1[4801] <= 16'b0000000000000000;
        weights1[4802] <= 16'b0000000000000000;
        weights1[4803] <= 16'b0000000000000000;
        weights1[4804] <= 16'b0000000000000000;
        weights1[4805] <= 16'b0000000000000000;
        weights1[4806] <= 16'b0000000000000000;
        weights1[4807] <= 16'b0000000000000000;
        weights1[4808] <= 16'b0000000000000000;
        weights1[4809] <= 16'b0000000000000000;
        weights1[4810] <= 16'b0000000000000000;
        weights1[4811] <= 16'b0000000000000000;
        weights1[4812] <= 16'b0000000000000000;
        weights1[4813] <= 16'b0000000000000000;
        weights1[4814] <= 16'b0000000000000000;
        weights1[4815] <= 16'b0000000000000000;
        weights1[4816] <= 16'b0000000000000000;
        weights1[4817] <= 16'b0000000000000000;
        weights1[4818] <= 16'b0000000000000000;
        weights1[4819] <= 16'b0000000000000000;
        weights1[4820] <= 16'b0000000000000000;
        weights1[4821] <= 16'b0000000000000000;
        weights1[4822] <= 16'b0000000000000000;
        weights1[4823] <= 16'b0000000000000000;
        weights1[4824] <= 16'b0000000000000000;
        weights1[4825] <= 16'b0000000000000000;
        weights1[4826] <= 16'b0000000000000000;
        weights1[4827] <= 16'b0000000000000000;
        weights1[4828] <= 16'b0000000000000000;
        weights1[4829] <= 16'b0000000000000000;
        weights1[4830] <= 16'b0000000000000000;
        weights1[4831] <= 16'b0000000000000000;
        weights1[4832] <= 16'b0000000000000000;
        weights1[4833] <= 16'b0000000000000000;
        weights1[4834] <= 16'b0000000000000000;
        weights1[4835] <= 16'b0000000000000000;
        weights1[4836] <= 16'b0000000000000000;
        weights1[4837] <= 16'b0000000000000000;
        weights1[4838] <= 16'b0000000000000000;
        weights1[4839] <= 16'b0000000000000000;
        weights1[4840] <= 16'b0000000000000000;
        weights1[4841] <= 16'b0000000000000000;
        weights1[4842] <= 16'b0000000000000000;
        weights1[4843] <= 16'b0000000000000000;
        weights1[4844] <= 16'b0000000000000000;
        weights1[4845] <= 16'b0000000000000000;
        weights1[4846] <= 16'b0000000000000000;
        weights1[4847] <= 16'b0000000000000000;
        weights1[4848] <= 16'b0000000000000000;
        weights1[4849] <= 16'b0000000000000000;
        weights1[4850] <= 16'b0000000000000000;
        weights1[4851] <= 16'b0000000000000000;
        weights1[4852] <= 16'b0000000000000000;
        weights1[4853] <= 16'b0000000000000000;
        weights1[4854] <= 16'b0000000000000000;
        weights1[4855] <= 16'b0000000000000000;
        weights1[4856] <= 16'b0000000000000000;
        weights1[4857] <= 16'b0000000000000000;
        weights1[4858] <= 16'b0000000000000000;
        weights1[4859] <= 16'b0000000000000000;
        weights1[4860] <= 16'b0000000000000000;
        weights1[4861] <= 16'b0000000000000000;
        weights1[4862] <= 16'b0000000000000000;
        weights1[4863] <= 16'b0000000000000000;
        weights1[4864] <= 16'b0000000000000000;
        weights1[4865] <= 16'b0000000000000000;
        weights1[4866] <= 16'b0000000000000000;
        weights1[4867] <= 16'b0000000000000000;
        weights1[4868] <= 16'b0000000000000000;
        weights1[4869] <= 16'b0000000000000000;
        weights1[4870] <= 16'b0000000000000000;
        weights1[4871] <= 16'b0000000000000000;
        weights1[4872] <= 16'b0000000000000000;
        weights1[4873] <= 16'b0000000000000000;
        weights1[4874] <= 16'b0000000000000000;
        weights1[4875] <= 16'b0000000000000000;
        weights1[4876] <= 16'b0000000000000000;
        weights1[4877] <= 16'b0000000000000000;
        weights1[4878] <= 16'b0000000000000000;
        weights1[4879] <= 16'b0000000000000000;
        weights1[4880] <= 16'b0000000000000000;
        weights1[4881] <= 16'b0000000000000000;
        weights1[4882] <= 16'b0000000000000000;
        weights1[4883] <= 16'b0000000000000000;
        weights1[4884] <= 16'b0000000000000000;
        weights1[4885] <= 16'b0000000000000000;
        weights1[4886] <= 16'b0000000000000000;
        weights1[4887] <= 16'b0000000000000000;
        weights1[4888] <= 16'b0000000000000000;
        weights1[4889] <= 16'b0000000000000000;
        weights1[4890] <= 16'b0000000000000000;
        weights1[4891] <= 16'b0000000000000000;
        weights1[4892] <= 16'b0000000000000000;
        weights1[4893] <= 16'b0000000000000000;
        weights1[4894] <= 16'b0000000000000000;
        weights1[4895] <= 16'b0000000000000000;
        weights1[4896] <= 16'b0000000000000000;
        weights1[4897] <= 16'b0000000000000000;
        weights1[4898] <= 16'b0000000000000000;
        weights1[4899] <= 16'b0000000000000000;
        weights1[4900] <= 16'b0000000000000000;
        weights1[4901] <= 16'b0000000000000000;
        weights1[4902] <= 16'b0000000000000000;
        weights1[4903] <= 16'b0000000000000000;
        weights1[4904] <= 16'b0000000000000000;
        weights1[4905] <= 16'b0000000000000000;
        weights1[4906] <= 16'b0000000000000000;
        weights1[4907] <= 16'b0000000000000000;
        weights1[4908] <= 16'b0000000000000000;
        weights1[4909] <= 16'b0000000000000000;
        weights1[4910] <= 16'b0000000000000000;
        weights1[4911] <= 16'b0000000000000000;
        weights1[4912] <= 16'b0000000000000000;
        weights1[4913] <= 16'b0000000000000000;
        weights1[4914] <= 16'b0000000000000000;
        weights1[4915] <= 16'b0000000000000000;
        weights1[4916] <= 16'b0000000000000000;
        weights1[4917] <= 16'b0000000000000000;
        weights1[4918] <= 16'b0000000000000000;
        weights1[4919] <= 16'b0000000000000000;
        weights1[4920] <= 16'b0000000000000000;
        weights1[4921] <= 16'b0000000000000000;
        weights1[4922] <= 16'b0000000000000000;
        weights1[4923] <= 16'b0000000000000000;
        weights1[4924] <= 16'b0000000000000000;
        weights1[4925] <= 16'b0000000000000000;
        weights1[4926] <= 16'b0000000000000000;
        weights1[4927] <= 16'b0000000000000000;
        weights1[4928] <= 16'b0000000000000000;
        weights1[4929] <= 16'b0000000000000000;
        weights1[4930] <= 16'b0000000000000000;
        weights1[4931] <= 16'b0000000000000000;
        weights1[4932] <= 16'b0000000000000000;
        weights1[4933] <= 16'b0000000000000000;
        weights1[4934] <= 16'b0000000000000000;
        weights1[4935] <= 16'b0000000000000000;
        weights1[4936] <= 16'b0000000000000000;
        weights1[4937] <= 16'b0000000000000000;
        weights1[4938] <= 16'b0000000000000000;
        weights1[4939] <= 16'b0000000000000000;
        weights1[4940] <= 16'b0000000000000000;
        weights1[4941] <= 16'b0000000000000000;
        weights1[4942] <= 16'b0000000000000000;
        weights1[4943] <= 16'b0000000000000000;
        weights1[4944] <= 16'b0000000000000000;
        weights1[4945] <= 16'b0000000000000000;
        weights1[4946] <= 16'b0000000000000000;
        weights1[4947] <= 16'b0000000000000000;
        weights1[4948] <= 16'b0000000000000000;
        weights1[4949] <= 16'b0000000000000000;
        weights1[4950] <= 16'b0000000000000000;
        weights1[4951] <= 16'b0000000000000000;
        weights1[4952] <= 16'b0000000000000000;
        weights1[4953] <= 16'b0000000000000000;
        weights1[4954] <= 16'b0000000000000000;
        weights1[4955] <= 16'b0000000000000000;
        weights1[4956] <= 16'b0000000000000000;
        weights1[4957] <= 16'b0000000000000000;
        weights1[4958] <= 16'b0000000000000000;
        weights1[4959] <= 16'b0000000000000000;
        weights1[4960] <= 16'b0000000000000000;
        weights1[4961] <= 16'b0000000000000000;
        weights1[4962] <= 16'b0000000000000000;
        weights1[4963] <= 16'b0000000000000000;
        weights1[4964] <= 16'b0000000000000000;
        weights1[4965] <= 16'b0000000000000000;
        weights1[4966] <= 16'b0000000000000000;
        weights1[4967] <= 16'b0000000000000000;
        weights1[4968] <= 16'b0000000000000000;
        weights1[4969] <= 16'b0000000000000000;
        weights1[4970] <= 16'b0000000000000000;
        weights1[4971] <= 16'b0000000000000000;
        weights1[4972] <= 16'b0000000000000000;
        weights1[4973] <= 16'b0000000000000000;
        weights1[4974] <= 16'b0000000000000000;
        weights1[4975] <= 16'b0000000000000000;
        weights1[4976] <= 16'b0000000000000000;
        weights1[4977] <= 16'b0000000000000000;
        weights1[4978] <= 16'b0000000000000000;
        weights1[4979] <= 16'b0000000000000000;
        weights1[4980] <= 16'b0000000000000000;
        weights1[4981] <= 16'b0000000000000000;
        weights1[4982] <= 16'b0000000000000000;
        weights1[4983] <= 16'b0000000000000000;
        weights1[4984] <= 16'b0000000000000000;
        weights1[4985] <= 16'b0000000000000000;
        weights1[4986] <= 16'b0000000000000000;
        weights1[4987] <= 16'b0000000000000000;
        weights1[4988] <= 16'b0000000000000000;
        weights1[4989] <= 16'b0000000000000000;
        weights1[4990] <= 16'b0000000000000000;
        weights1[4991] <= 16'b0000000000000000;
        weights1[4992] <= 16'b0000000000000000;
        weights1[4993] <= 16'b0000000000000000;
        weights1[4994] <= 16'b0000000000000000;
        weights1[4995] <= 16'b0000000000000000;
        weights1[4996] <= 16'b0000000000000000;
        weights1[4997] <= 16'b0000000000000000;
        weights1[4998] <= 16'b0000000000000000;
        weights1[4999] <= 16'b0000000000000000;
        weights1[5000] <= 16'b0000000000000000;
        weights1[5001] <= 16'b0000000000000000;
        weights1[5002] <= 16'b0000000000000000;
        weights1[5003] <= 16'b0000000000000000;
        weights1[5004] <= 16'b0000000000000000;
        weights1[5005] <= 16'b0000000000000000;
        weights1[5006] <= 16'b0000000000000000;
        weights1[5007] <= 16'b0000000000000000;
        weights1[5008] <= 16'b0000000000000000;
        weights1[5009] <= 16'b0000000000000000;
        weights1[5010] <= 16'b0000000000000000;
        weights1[5011] <= 16'b0000000000000000;
        weights1[5012] <= 16'b0000000000000000;
        weights1[5013] <= 16'b0000000000000000;
        weights1[5014] <= 16'b0000000000000000;
        weights1[5015] <= 16'b0000000000000000;
        weights1[5016] <= 16'b0000000000000000;
        weights1[5017] <= 16'b0000000000000000;
        weights1[5018] <= 16'b0000000000000000;
        weights1[5019] <= 16'b0000000000000000;
        weights1[5020] <= 16'b0000000000000000;
        weights1[5021] <= 16'b0000000000000000;
        weights1[5022] <= 16'b0000000000000000;
        weights1[5023] <= 16'b0000000000000000;
        weights1[5024] <= 16'b0000000000000000;
        weights1[5025] <= 16'b0000000000000000;
        weights1[5026] <= 16'b0000000000000000;
        weights1[5027] <= 16'b0000000000000000;
        weights1[5028] <= 16'b0000000000000000;
        weights1[5029] <= 16'b0000000000000000;
        weights1[5030] <= 16'b0000000000000000;
        weights1[5031] <= 16'b0000000000000000;
        weights1[5032] <= 16'b0000000000000000;
        weights1[5033] <= 16'b0000000000000000;
        weights1[5034] <= 16'b0000000000000000;
        weights1[5035] <= 16'b0000000000000000;
        weights1[5036] <= 16'b0000000000000000;
        weights1[5037] <= 16'b0000000000000000;
        weights1[5038] <= 16'b0000000000000000;
        weights1[5039] <= 16'b0000000000000000;
        weights1[5040] <= 16'b0000000000000000;
        weights1[5041] <= 16'b0000000000000000;
        weights1[5042] <= 16'b0000000000000000;
        weights1[5043] <= 16'b0000000000000000;
        weights1[5044] <= 16'b0000000000000000;
        weights1[5045] <= 16'b0000000000000000;
        weights1[5046] <= 16'b0000000000000000;
        weights1[5047] <= 16'b0000000000000000;
        weights1[5048] <= 16'b0000000000000000;
        weights1[5049] <= 16'b0000000000000000;
        weights1[5050] <= 16'b0000000000000000;
        weights1[5051] <= 16'b0000000000000000;
        weights1[5052] <= 16'b0000000000000000;
        weights1[5053] <= 16'b0000000000000000;
        weights1[5054] <= 16'b0000000000000000;
        weights1[5055] <= 16'b0000000000000000;
        weights1[5056] <= 16'b0000000000000000;
        weights1[5057] <= 16'b0000000000000000;
        weights1[5058] <= 16'b0000000000000000;
        weights1[5059] <= 16'b0000000000000000;
        weights1[5060] <= 16'b0000000000000000;
        weights1[5061] <= 16'b0000000000000000;
        weights1[5062] <= 16'b0000000000000000;
        weights1[5063] <= 16'b0000000000000000;
        weights1[5064] <= 16'b0000000000000000;
        weights1[5065] <= 16'b0000000000000000;
        weights1[5066] <= 16'b0000000000000000;
        weights1[5067] <= 16'b0000000000000000;
        weights1[5068] <= 16'b0000000000000000;
        weights1[5069] <= 16'b0000000000000000;
        weights1[5070] <= 16'b0000000000000000;
        weights1[5071] <= 16'b0000000000000000;
        weights1[5072] <= 16'b0000000000000000;
        weights1[5073] <= 16'b0000000000000000;
        weights1[5074] <= 16'b0000000000000000;
        weights1[5075] <= 16'b0000000000000000;
        weights1[5076] <= 16'b0000000000000000;
        weights1[5077] <= 16'b0000000000000000;
        weights1[5078] <= 16'b0000000000000000;
        weights1[5079] <= 16'b0000000000000000;
        weights1[5080] <= 16'b0000000000000000;
        weights1[5081] <= 16'b0000000000000000;
        weights1[5082] <= 16'b0000000000000000;
        weights1[5083] <= 16'b0000000000000000;
        weights1[5084] <= 16'b0000000000000000;
        weights1[5085] <= 16'b0000000000000000;
        weights1[5086] <= 16'b0000000000000000;
        weights1[5087] <= 16'b0000000000000000;
        weights1[5088] <= 16'b0000000000000000;
        weights1[5089] <= 16'b0000000000000000;
        weights1[5090] <= 16'b0000000000000000;
        weights1[5091] <= 16'b0000000000000000;
        weights1[5092] <= 16'b0000000000000000;
        weights1[5093] <= 16'b0000000000000000;
        weights1[5094] <= 16'b0000000000000000;
        weights1[5095] <= 16'b0000000000000000;
        weights1[5096] <= 16'b0000000000000000;
        weights1[5097] <= 16'b0000000000000000;
        weights1[5098] <= 16'b0000000000000000;
        weights1[5099] <= 16'b0000000000000000;
        weights1[5100] <= 16'b0000000000000000;
        weights1[5101] <= 16'b0000000000000000;
        weights1[5102] <= 16'b0000000000000000;
        weights1[5103] <= 16'b0000000000000000;
        weights1[5104] <= 16'b0000000000000000;
        weights1[5105] <= 16'b0000000000000000;
        weights1[5106] <= 16'b0000000000000000;
        weights1[5107] <= 16'b0000000000000000;
        weights1[5108] <= 16'b0000000000000000;
        weights1[5109] <= 16'b0000000000000000;
        weights1[5110] <= 16'b0000000000000000;
        weights1[5111] <= 16'b0000000000000000;
        weights1[5112] <= 16'b0000000000000000;
        weights1[5113] <= 16'b0000000000000000;
        weights1[5114] <= 16'b0000000000000000;
        weights1[5115] <= 16'b0000000000000000;
        weights1[5116] <= 16'b0000000000000000;
        weights1[5117] <= 16'b0000000000000000;
        weights1[5118] <= 16'b0000000000000000;
        weights1[5119] <= 16'b0000000000000000;
        weights1[5120] <= 16'b0000000000000000;
        weights1[5121] <= 16'b0000000000000000;
        weights1[5122] <= 16'b0000000000000000;
        weights1[5123] <= 16'b0000000000000000;
        weights1[5124] <= 16'b0000000000000000;
        weights1[5125] <= 16'b0000000000000000;
        weights1[5126] <= 16'b0000000000000000;
        weights1[5127] <= 16'b0000000000000000;
        weights1[5128] <= 16'b0000000000000000;
        weights1[5129] <= 16'b0000000000000000;
        weights1[5130] <= 16'b0000000000000000;
        weights1[5131] <= 16'b0000000000000000;
        weights1[5132] <= 16'b0000000000000000;
        weights1[5133] <= 16'b0000000000000000;
        weights1[5134] <= 16'b0000000000000000;
        weights1[5135] <= 16'b0000000000000000;
        weights1[5136] <= 16'b0000000000000000;
        weights1[5137] <= 16'b0000000000000000;
        weights1[5138] <= 16'b0000000000000000;
        weights1[5139] <= 16'b0000000000000000;
        weights1[5140] <= 16'b0000000000000000;
        weights1[5141] <= 16'b0000000000000000;
        weights1[5142] <= 16'b0000000000000000;
        weights1[5143] <= 16'b0000000000000000;
        weights1[5144] <= 16'b0000000000000000;
        weights1[5145] <= 16'b0000000000000000;
        weights1[5146] <= 16'b0000000000000000;
        weights1[5147] <= 16'b0000000000000000;
        weights1[5148] <= 16'b0000000000000000;
        weights1[5149] <= 16'b0000000000000000;
        weights1[5150] <= 16'b0000000000000000;
        weights1[5151] <= 16'b0000000000000000;
        weights1[5152] <= 16'b0000000000000000;
        weights1[5153] <= 16'b0000000000000000;
        weights1[5154] <= 16'b0000000000000000;
        weights1[5155] <= 16'b0000000000000000;
        weights1[5156] <= 16'b0000000000000000;
        weights1[5157] <= 16'b0000000000000000;
        weights1[5158] <= 16'b0000000000000000;
        weights1[5159] <= 16'b0000000000000000;
        weights1[5160] <= 16'b0000000000000000;
        weights1[5161] <= 16'b0000000000000000;
        weights1[5162] <= 16'b0000000000000000;
        weights1[5163] <= 16'b0000000000000000;
        weights1[5164] <= 16'b0000000000000000;
        weights1[5165] <= 16'b0000000000000000;
        weights1[5166] <= 16'b0000000000000000;
        weights1[5167] <= 16'b0000000000000000;
        weights1[5168] <= 16'b0000000000000000;
        weights1[5169] <= 16'b0000000000000000;
        weights1[5170] <= 16'b0000000000000000;
        weights1[5171] <= 16'b0000000000000000;
        weights1[5172] <= 16'b0000000000000000;
        weights1[5173] <= 16'b0000000000000000;
        weights1[5174] <= 16'b0000000000000000;
        weights1[5175] <= 16'b0000000000000000;
        weights1[5176] <= 16'b0000000000000000;
        weights1[5177] <= 16'b0000000000000000;
        weights1[5178] <= 16'b0000000000000000;
        weights1[5179] <= 16'b0000000000000000;
        weights1[5180] <= 16'b0000000000000000;
        weights1[5181] <= 16'b0000000000000000;
        weights1[5182] <= 16'b0000000000000000;
        weights1[5183] <= 16'b0000000000000000;
        weights1[5184] <= 16'b0000000000000000;
        weights1[5185] <= 16'b0000000000000000;
        weights1[5186] <= 16'b0000000000000000;
        weights1[5187] <= 16'b0000000000000000;
        weights1[5188] <= 16'b0000000000000000;
        weights1[5189] <= 16'b0000000000000000;
        weights1[5190] <= 16'b0000000000000000;
        weights1[5191] <= 16'b0000000000000000;
        weights1[5192] <= 16'b0000000000000000;
        weights1[5193] <= 16'b0000000000000000;
        weights1[5194] <= 16'b0000000000000000;
        weights1[5195] <= 16'b0000000000000000;
        weights1[5196] <= 16'b0000000000000000;
        weights1[5197] <= 16'b0000000000000000;
        weights1[5198] <= 16'b0000000000000000;
        weights1[5199] <= 16'b0000000000000000;
        weights1[5200] <= 16'b0000000000000000;
        weights1[5201] <= 16'b0000000000000000;
        weights1[5202] <= 16'b0000000000000000;
        weights1[5203] <= 16'b0000000000000000;
        weights1[5204] <= 16'b0000000000000000;
        weights1[5205] <= 16'b0000000000000000;
        weights1[5206] <= 16'b0000000000000000;
        weights1[5207] <= 16'b0000000000000000;
        weights1[5208] <= 16'b0000000000000000;
        weights1[5209] <= 16'b0000000000000000;
        weights1[5210] <= 16'b0000000000000000;
        weights1[5211] <= 16'b0000000000000000;
        weights1[5212] <= 16'b0000000000000000;
        weights1[5213] <= 16'b0000000000000000;
        weights1[5214] <= 16'b0000000000000000;
        weights1[5215] <= 16'b0000000000000000;
        weights1[5216] <= 16'b0000000000000000;
        weights1[5217] <= 16'b0000000000000000;
        weights1[5218] <= 16'b0000000000000000;
        weights1[5219] <= 16'b0000000000000000;
        weights1[5220] <= 16'b0000000000000000;
        weights1[5221] <= 16'b0000000000000000;
        weights1[5222] <= 16'b0000000000000000;
        weights1[5223] <= 16'b0000000000000000;
        weights1[5224] <= 16'b0000000000000000;
        weights1[5225] <= 16'b0000000000000000;
        weights1[5226] <= 16'b0000000000000000;
        weights1[5227] <= 16'b0000000000000000;
        weights1[5228] <= 16'b0000000000000000;
        weights1[5229] <= 16'b0000000000000000;
        weights1[5230] <= 16'b0000000000000000;
        weights1[5231] <= 16'b0000000000000000;
        weights1[5232] <= 16'b0000000000000000;
        weights1[5233] <= 16'b0000000000000000;
        weights1[5234] <= 16'b0000000000000000;
        weights1[5235] <= 16'b0000000000000000;
        weights1[5236] <= 16'b0000000000000000;
        weights1[5237] <= 16'b0000000000000000;
        weights1[5238] <= 16'b0000000000000000;
        weights1[5239] <= 16'b0000000000000000;
        weights1[5240] <= 16'b0000000000000000;
        weights1[5241] <= 16'b0000000000000000;
        weights1[5242] <= 16'b0000000000000000;
        weights1[5243] <= 16'b0000000000000000;
        weights1[5244] <= 16'b0000000000000000;
        weights1[5245] <= 16'b0000000000000000;
        weights1[5246] <= 16'b0000000000000000;
        weights1[5247] <= 16'b0000000000000000;
        weights1[5248] <= 16'b0000000000000000;
        weights1[5249] <= 16'b0000000000000000;
        weights1[5250] <= 16'b0000000000000000;
        weights1[5251] <= 16'b0000000000000000;
        weights1[5252] <= 16'b0000000000000000;
        weights1[5253] <= 16'b0000000000000000;
        weights1[5254] <= 16'b0000000000000000;
        weights1[5255] <= 16'b0000000000000000;
        weights1[5256] <= 16'b0000000000000000;
        weights1[5257] <= 16'b0000000000000000;
        weights1[5258] <= 16'b0000000000000000;
        weights1[5259] <= 16'b0000000000000000;
        weights1[5260] <= 16'b0000000000000000;
        weights1[5261] <= 16'b0000000000000000;
        weights1[5262] <= 16'b0000000000000000;
        weights1[5263] <= 16'b0000000000000000;
        weights1[5264] <= 16'b0000000000000000;
        weights1[5265] <= 16'b0000000000000000;
        weights1[5266] <= 16'b0000000000000000;
        weights1[5267] <= 16'b0000000000000000;
        weights1[5268] <= 16'b0000000000000000;
        weights1[5269] <= 16'b0000000000000000;
        weights1[5270] <= 16'b0000000000000000;
        weights1[5271] <= 16'b0000000000000000;
        weights1[5272] <= 16'b0000000000000000;
        weights1[5273] <= 16'b0000000000000000;
        weights1[5274] <= 16'b0000000000000000;
        weights1[5275] <= 16'b0000000000000000;
        weights1[5276] <= 16'b0000000000000000;
        weights1[5277] <= 16'b0000000000000000;
        weights1[5278] <= 16'b0000000000000000;
        weights1[5279] <= 16'b0000000000000000;
        weights1[5280] <= 16'b0000000000000000;
        weights1[5281] <= 16'b0000000000000000;
        weights1[5282] <= 16'b0000000000000000;
        weights1[5283] <= 16'b0000000000000000;
        weights1[5284] <= 16'b0000000000000000;
        weights1[5285] <= 16'b0000000000000000;
        weights1[5286] <= 16'b0000000000000000;
        weights1[5287] <= 16'b0000000000000000;
        weights1[5288] <= 16'b0000000000000000;
        weights1[5289] <= 16'b0000000000000000;
        weights1[5290] <= 16'b0000000000000000;
        weights1[5291] <= 16'b0000000000000000;
        weights1[5292] <= 16'b0000000000000000;
        weights1[5293] <= 16'b0000000000000000;
        weights1[5294] <= 16'b0000000000000000;
        weights1[5295] <= 16'b0000000000000000;
        weights1[5296] <= 16'b0000000000000000;
        weights1[5297] <= 16'b0000000000000000;
        weights1[5298] <= 16'b0000000000000000;
        weights1[5299] <= 16'b0000000000000000;
        weights1[5300] <= 16'b0000000000000000;
        weights1[5301] <= 16'b0000000000000000;
        weights1[5302] <= 16'b0000000000000000;
        weights1[5303] <= 16'b0000000000000000;
        weights1[5304] <= 16'b0000000000000000;
        weights1[5305] <= 16'b0000000000000000;
        weights1[5306] <= 16'b0000000000000000;
        weights1[5307] <= 16'b0000000000000000;
        weights1[5308] <= 16'b0000000000000000;
        weights1[5309] <= 16'b0000000000000000;
        weights1[5310] <= 16'b0000000000000000;
        weights1[5311] <= 16'b0000000000000000;
        weights1[5312] <= 16'b0000000000000000;
        weights1[5313] <= 16'b0000000000000000;
        weights1[5314] <= 16'b0000000000000000;
        weights1[5315] <= 16'b0000000000000000;
        weights1[5316] <= 16'b0000000000000000;
        weights1[5317] <= 16'b0000000000000000;
        weights1[5318] <= 16'b0000000000000000;
        weights1[5319] <= 16'b0000000000000000;
        weights1[5320] <= 16'b0000000000000000;
        weights1[5321] <= 16'b0000000000000000;
        weights1[5322] <= 16'b0000000000000000;
        weights1[5323] <= 16'b0000000000000000;
        weights1[5324] <= 16'b0000000000000000;
        weights1[5325] <= 16'b0000000000000000;
        weights1[5326] <= 16'b0000000000000000;
        weights1[5327] <= 16'b0000000000000000;
        weights1[5328] <= 16'b0000000000000000;
        weights1[5329] <= 16'b0000000000000000;
        weights1[5330] <= 16'b0000000000000000;
        weights1[5331] <= 16'b0000000000000000;
        weights1[5332] <= 16'b0000000000000000;
        weights1[5333] <= 16'b0000000000000000;
        weights1[5334] <= 16'b0000000000000000;
        weights1[5335] <= 16'b0000000000000000;
        weights1[5336] <= 16'b0000000000000000;
        weights1[5337] <= 16'b0000000000000000;
        weights1[5338] <= 16'b0000000000000000;
        weights1[5339] <= 16'b0000000000000000;
        weights1[5340] <= 16'b0000000000000000;
        weights1[5341] <= 16'b0000000000000000;
        weights1[5342] <= 16'b0000000000000000;
        weights1[5343] <= 16'b0000000000000000;
        weights1[5344] <= 16'b0000000000000000;
        weights1[5345] <= 16'b0000000000000000;
        weights1[5346] <= 16'b0000000000000000;
        weights1[5347] <= 16'b0000000000000000;
        weights1[5348] <= 16'b0000000000000000;
        weights1[5349] <= 16'b0000000000000000;
        weights1[5350] <= 16'b0000000000000000;
        weights1[5351] <= 16'b0000000000000000;
        weights1[5352] <= 16'b0000000000000000;
        weights1[5353] <= 16'b0000000000000000;
        weights1[5354] <= 16'b0000000000000000;
        weights1[5355] <= 16'b0000000000000000;
        weights1[5356] <= 16'b0000000000000000;
        weights1[5357] <= 16'b0000000000000000;
        weights1[5358] <= 16'b0000000000000000;
        weights1[5359] <= 16'b0000000000000000;
        weights1[5360] <= 16'b0000000000000000;
        weights1[5361] <= 16'b0000000000000000;
        weights1[5362] <= 16'b0000000000000000;
        weights1[5363] <= 16'b0000000000000000;
        weights1[5364] <= 16'b0000000000000000;
        weights1[5365] <= 16'b0000000000000000;
        weights1[5366] <= 16'b0000000000000000;
        weights1[5367] <= 16'b0000000000000000;
        weights1[5368] <= 16'b0000000000000000;
        weights1[5369] <= 16'b0000000000000000;
        weights1[5370] <= 16'b0000000000000000;
        weights1[5371] <= 16'b0000000000000000;
        weights1[5372] <= 16'b0000000000000000;
        weights1[5373] <= 16'b0000000000000000;
        weights1[5374] <= 16'b0000000000000000;
        weights1[5375] <= 16'b0000000000000000;
        weights1[5376] <= 16'b0000000000000000;
        weights1[5377] <= 16'b0000000000000000;
        weights1[5378] <= 16'b0000000000000000;
        weights1[5379] <= 16'b0000000000000000;
        weights1[5380] <= 16'b0000000000000000;
        weights1[5381] <= 16'b0000000000000000;
        weights1[5382] <= 16'b0000000000000000;
        weights1[5383] <= 16'b0000000000000000;
        weights1[5384] <= 16'b0000000000000000;
        weights1[5385] <= 16'b0000000000000000;
        weights1[5386] <= 16'b0000000000000000;
        weights1[5387] <= 16'b0000000000000000;
        weights1[5388] <= 16'b0000000000000000;
        weights1[5389] <= 16'b0000000000000000;
        weights1[5390] <= 16'b0000000000000000;
        weights1[5391] <= 16'b0000000000000000;
        weights1[5392] <= 16'b0000000000000000;
        weights1[5393] <= 16'b0000000000000000;
        weights1[5394] <= 16'b0000000000000000;
        weights1[5395] <= 16'b0000000000000000;
        weights1[5396] <= 16'b0000000000000000;
        weights1[5397] <= 16'b0000000000000000;
        weights1[5398] <= 16'b0000000000000000;
        weights1[5399] <= 16'b0000000000000000;
        weights1[5400] <= 16'b0000000000000000;
        weights1[5401] <= 16'b0000000000000000;
        weights1[5402] <= 16'b0000000000000000;
        weights1[5403] <= 16'b0000000000000000;
        weights1[5404] <= 16'b0000000000000000;
        weights1[5405] <= 16'b0000000000000000;
        weights1[5406] <= 16'b0000000000000000;
        weights1[5407] <= 16'b0000000000000000;
        weights1[5408] <= 16'b0000000000000000;
        weights1[5409] <= 16'b0000000000000000;
        weights1[5410] <= 16'b0000000000000000;
        weights1[5411] <= 16'b0000000000000000;
        weights1[5412] <= 16'b0000000000000000;
        weights1[5413] <= 16'b0000000000000000;
        weights1[5414] <= 16'b0000000000000000;
        weights1[5415] <= 16'b0000000000000000;
        weights1[5416] <= 16'b0000000000000000;
        weights1[5417] <= 16'b0000000000000000;
        weights1[5418] <= 16'b0000000000000000;
        weights1[5419] <= 16'b0000000000000000;
        weights1[5420] <= 16'b0000000000000000;
        weights1[5421] <= 16'b0000000000000000;
        weights1[5422] <= 16'b0000000000000000;
        weights1[5423] <= 16'b0000000000000000;
        weights1[5424] <= 16'b0000000000000000;
        weights1[5425] <= 16'b0000000000000000;
        weights1[5426] <= 16'b0000000000000000;
        weights1[5427] <= 16'b0000000000000000;
        weights1[5428] <= 16'b0000000000000000;
        weights1[5429] <= 16'b0000000000000000;
        weights1[5430] <= 16'b0000000000000000;
        weights1[5431] <= 16'b0000000000000000;
        weights1[5432] <= 16'b0000000000000000;
        weights1[5433] <= 16'b0000000000000000;
        weights1[5434] <= 16'b0000000000000000;
        weights1[5435] <= 16'b0000000000000000;
        weights1[5436] <= 16'b0000000000000000;
        weights1[5437] <= 16'b0000000000000000;
        weights1[5438] <= 16'b0000000000000000;
        weights1[5439] <= 16'b0000000000000000;
        weights1[5440] <= 16'b0000000000000000;
        weights1[5441] <= 16'b0000000000000000;
        weights1[5442] <= 16'b0000000000000000;
        weights1[5443] <= 16'b0000000000000000;
        weights1[5444] <= 16'b0000000000000000;
        weights1[5445] <= 16'b0000000000000000;
        weights1[5446] <= 16'b0000000000000000;
        weights1[5447] <= 16'b0000000000000000;
        weights1[5448] <= 16'b0000000000000000;
        weights1[5449] <= 16'b0000000000000000;
        weights1[5450] <= 16'b0000000000000000;
        weights1[5451] <= 16'b0000000000000000;
        weights1[5452] <= 16'b0000000000000000;
        weights1[5453] <= 16'b0000000000000000;
        weights1[5454] <= 16'b0000000000000000;
        weights1[5455] <= 16'b0000000000000000;
        weights1[5456] <= 16'b0000000000000000;
        weights1[5457] <= 16'b0000000000000000;
        weights1[5458] <= 16'b0000000000000000;
        weights1[5459] <= 16'b0000000000000000;
        weights1[5460] <= 16'b0000000000000000;
        weights1[5461] <= 16'b0000000000000000;
        weights1[5462] <= 16'b0000000000000000;
        weights1[5463] <= 16'b0000000000000000;
        weights1[5464] <= 16'b0000000000000000;
        weights1[5465] <= 16'b0000000000000000;
        weights1[5466] <= 16'b0000000000000000;
        weights1[5467] <= 16'b0000000000000000;
        weights1[5468] <= 16'b0000000000000000;
        weights1[5469] <= 16'b0000000000000000;
        weights1[5470] <= 16'b0000000000000000;
        weights1[5471] <= 16'b0000000000000000;
        weights1[5472] <= 16'b0000000000000000;
        weights1[5473] <= 16'b0000000000000000;
        weights1[5474] <= 16'b0000000000000000;
        weights1[5475] <= 16'b0000000000000000;
        weights1[5476] <= 16'b0000000000000000;
        weights1[5477] <= 16'b0000000000000000;
        weights1[5478] <= 16'b0000000000000000;
        weights1[5479] <= 16'b0000000000000000;
        weights1[5480] <= 16'b0000000000000000;
        weights1[5481] <= 16'b0000000000000000;
        weights1[5482] <= 16'b0000000000000000;
        weights1[5483] <= 16'b0000000000000000;
        weights1[5484] <= 16'b0000000000000000;
        weights1[5485] <= 16'b0000000000000000;
        weights1[5486] <= 16'b0000000000000000;
        weights1[5487] <= 16'b0000000000000000;
        weights1[5488] <= 16'b0000000000000000;
        weights1[5489] <= 16'b0000000000000000;
        weights1[5490] <= 16'b0000000000000000;
        weights1[5491] <= 16'b0000000000000010;
        weights1[5492] <= 16'b1111111111111111;
        weights1[5493] <= 16'b1111111111111101;
        weights1[5494] <= 16'b1111111111111000;
        weights1[5495] <= 16'b1111111111110011;
        weights1[5496] <= 16'b1111111111111010;
        weights1[5497] <= 16'b1111111111110010;
        weights1[5498] <= 16'b1111111111011110;
        weights1[5499] <= 16'b1111111111101111;
        weights1[5500] <= 16'b1111111111111110;
        weights1[5501] <= 16'b1111111111111111;
        weights1[5502] <= 16'b0000000000001001;
        weights1[5503] <= 16'b0000000000000101;
        weights1[5504] <= 16'b1111111111110111;
        weights1[5505] <= 16'b1111111111111101;
        weights1[5506] <= 16'b1111111111110100;
        weights1[5507] <= 16'b1111111111101100;
        weights1[5508] <= 16'b1111111111110111;
        weights1[5509] <= 16'b0000000000000000;
        weights1[5510] <= 16'b0000000000000100;
        weights1[5511] <= 16'b0000000000000011;
        weights1[5512] <= 16'b0000000000000000;
        weights1[5513] <= 16'b0000000000000010;
        weights1[5514] <= 16'b0000000000000011;
        weights1[5515] <= 16'b0000000000000000;
        weights1[5516] <= 16'b0000000000000001;
        weights1[5517] <= 16'b0000000000000001;
        weights1[5518] <= 16'b0000000000000001;
        weights1[5519] <= 16'b1111111111111101;
        weights1[5520] <= 16'b1111111111111000;
        weights1[5521] <= 16'b1111111111111011;
        weights1[5522] <= 16'b1111111111111000;
        weights1[5523] <= 16'b1111111111110011;
        weights1[5524] <= 16'b1111111111111100;
        weights1[5525] <= 16'b1111111111111011;
        weights1[5526] <= 16'b1111111111101110;
        weights1[5527] <= 16'b1111111111111111;
        weights1[5528] <= 16'b1111111111111111;
        weights1[5529] <= 16'b1111111111110101;
        weights1[5530] <= 16'b0000000000000011;
        weights1[5531] <= 16'b1111111111110001;
        weights1[5532] <= 16'b1111111111110110;
        weights1[5533] <= 16'b1111111111111010;
        weights1[5534] <= 16'b0000000000000101;
        weights1[5535] <= 16'b1111111111110101;
        weights1[5536] <= 16'b1111111111110110;
        weights1[5537] <= 16'b1111111111111101;
        weights1[5538] <= 16'b1111111111111100;
        weights1[5539] <= 16'b0000000000000000;
        weights1[5540] <= 16'b1111111111111110;
        weights1[5541] <= 16'b0000000000000101;
        weights1[5542] <= 16'b0000000000000010;
        weights1[5543] <= 16'b0000000000000011;
        weights1[5544] <= 16'b0000000000000001;
        weights1[5545] <= 16'b0000000000000001;
        weights1[5546] <= 16'b1111111111111100;
        weights1[5547] <= 16'b1111111111111100;
        weights1[5548] <= 16'b1111111111110011;
        weights1[5549] <= 16'b1111111111110000;
        weights1[5550] <= 16'b1111111111110000;
        weights1[5551] <= 16'b1111111111110011;
        weights1[5552] <= 16'b1111111111110011;
        weights1[5553] <= 16'b1111111111110101;
        weights1[5554] <= 16'b1111111111111101;
        weights1[5555] <= 16'b1111111111111010;
        weights1[5556] <= 16'b1111111111111000;
        weights1[5557] <= 16'b0000000000000001;
        weights1[5558] <= 16'b1111111111110110;
        weights1[5559] <= 16'b0000000000000010;
        weights1[5560] <= 16'b1111111111110010;
        weights1[5561] <= 16'b1111111111110101;
        weights1[5562] <= 16'b1111111111111111;
        weights1[5563] <= 16'b0000000000000010;
        weights1[5564] <= 16'b0000000000000011;
        weights1[5565] <= 16'b1111111111111110;
        weights1[5566] <= 16'b1111111111111010;
        weights1[5567] <= 16'b1111111111111110;
        weights1[5568] <= 16'b1111111111111110;
        weights1[5569] <= 16'b0000000000000001;
        weights1[5570] <= 16'b0000000000000010;
        weights1[5571] <= 16'b0000000000000010;
        weights1[5572] <= 16'b0000000000000001;
        weights1[5573] <= 16'b0000000000000001;
        weights1[5574] <= 16'b0000000000000010;
        weights1[5575] <= 16'b1111111111111001;
        weights1[5576] <= 16'b1111111111111000;
        weights1[5577] <= 16'b1111111111110000;
        weights1[5578] <= 16'b1111111111101001;
        weights1[5579] <= 16'b1111111111111101;
        weights1[5580] <= 16'b1111111111101011;
        weights1[5581] <= 16'b0000000000000101;
        weights1[5582] <= 16'b1111111111111100;
        weights1[5583] <= 16'b0000000000001011;
        weights1[5584] <= 16'b1111111111111011;
        weights1[5585] <= 16'b0000000000011110;
        weights1[5586] <= 16'b0000000000000110;
        weights1[5587] <= 16'b0000000000000000;
        weights1[5588] <= 16'b1111111111111011;
        weights1[5589] <= 16'b1111111111110101;
        weights1[5590] <= 16'b0000000000000000;
        weights1[5591] <= 16'b1111111111110111;
        weights1[5592] <= 16'b0000000000001010;
        weights1[5593] <= 16'b1111111111111100;
        weights1[5594] <= 16'b0000000000000001;
        weights1[5595] <= 16'b1111111111101000;
        weights1[5596] <= 16'b1111111111101001;
        weights1[5597] <= 16'b1111111111110011;
        weights1[5598] <= 16'b1111111111110010;
        weights1[5599] <= 16'b0000000000000001;
        weights1[5600] <= 16'b0000000000000000;
        weights1[5601] <= 16'b0000000000000000;
        weights1[5602] <= 16'b1111111111111101;
        weights1[5603] <= 16'b1111111111101111;
        weights1[5604] <= 16'b0000000000000011;
        weights1[5605] <= 16'b1111111111110100;
        weights1[5606] <= 16'b1111111111110100;
        weights1[5607] <= 16'b1111111111110011;
        weights1[5608] <= 16'b0000000000000011;
        weights1[5609] <= 16'b1111111111110010;
        weights1[5610] <= 16'b1111111111100111;
        weights1[5611] <= 16'b1111111111100110;
        weights1[5612] <= 16'b0000000000000100;
        weights1[5613] <= 16'b1111111111111110;
        weights1[5614] <= 16'b1111111111101011;
        weights1[5615] <= 16'b1111111111111111;
        weights1[5616] <= 16'b1111111111110101;
        weights1[5617] <= 16'b0000000000001101;
        weights1[5618] <= 16'b0000000000000110;
        weights1[5619] <= 16'b1111111111111111;
        weights1[5620] <= 16'b1111111111101100;
        weights1[5621] <= 16'b1111111111101110;
        weights1[5622] <= 16'b1111111111111000;
        weights1[5623] <= 16'b0000000000010111;
        weights1[5624] <= 16'b1111111111111100;
        weights1[5625] <= 16'b1111111111101110;
        weights1[5626] <= 16'b1111111111110111;
        weights1[5627] <= 16'b1111111111111000;
        weights1[5628] <= 16'b1111111111111110;
        weights1[5629] <= 16'b1111111111111001;
        weights1[5630] <= 16'b1111111111111101;
        weights1[5631] <= 16'b1111111111110010;
        weights1[5632] <= 16'b1111111111110010;
        weights1[5633] <= 16'b1111111111100110;
        weights1[5634] <= 16'b1111111111110111;
        weights1[5635] <= 16'b1111111111101111;
        weights1[5636] <= 16'b1111111111110011;
        weights1[5637] <= 16'b0000000000000101;
        weights1[5638] <= 16'b1111111111111001;
        weights1[5639] <= 16'b0000000000000111;
        weights1[5640] <= 16'b1111111111111111;
        weights1[5641] <= 16'b0000000000010001;
        weights1[5642] <= 16'b1111111111111010;
        weights1[5643] <= 16'b1111111111110101;
        weights1[5644] <= 16'b1111111111111101;
        weights1[5645] <= 16'b1111111111110001;
        weights1[5646] <= 16'b1111111111101011;
        weights1[5647] <= 16'b1111111111111101;
        weights1[5648] <= 16'b1111111111011010;
        weights1[5649] <= 16'b1111111111110101;
        weights1[5650] <= 16'b1111111111111000;
        weights1[5651] <= 16'b1111111111110100;
        weights1[5652] <= 16'b1111111111111011;
        weights1[5653] <= 16'b1111111111111110;
        weights1[5654] <= 16'b1111111111110000;
        weights1[5655] <= 16'b1111111111110101;
        weights1[5656] <= 16'b1111111111111001;
        weights1[5657] <= 16'b1111111111111010;
        weights1[5658] <= 16'b0000000000001011;
        weights1[5659] <= 16'b1111111111110001;
        weights1[5660] <= 16'b0000000000000010;
        weights1[5661] <= 16'b0000000000000110;
        weights1[5662] <= 16'b0000000000010011;
        weights1[5663] <= 16'b1111111111110100;
        weights1[5664] <= 16'b1111111111111101;
        weights1[5665] <= 16'b0000000000001010;
        weights1[5666] <= 16'b0000000000000000;
        weights1[5667] <= 16'b0000000000000011;
        weights1[5668] <= 16'b1111111111111101;
        weights1[5669] <= 16'b1111111111111010;
        weights1[5670] <= 16'b0000000000010101;
        weights1[5671] <= 16'b0000000000001001;
        weights1[5672] <= 16'b0000000000001011;
        weights1[5673] <= 16'b0000000000001001;
        weights1[5674] <= 16'b0000000000000001;
        weights1[5675] <= 16'b1111111111101110;
        weights1[5676] <= 16'b1111111111110111;
        weights1[5677] <= 16'b1111111111111100;
        weights1[5678] <= 16'b1111111111110101;
        weights1[5679] <= 16'b0000000000000111;
        weights1[5680] <= 16'b1111111111111110;
        weights1[5681] <= 16'b1111111111111111;
        weights1[5682] <= 16'b1111111111110111;
        weights1[5683] <= 16'b1111111111110010;
        weights1[5684] <= 16'b1111111111111101;
        weights1[5685] <= 16'b1111111111110100;
        weights1[5686] <= 16'b1111111111111000;
        weights1[5687] <= 16'b1111111111111101;
        weights1[5688] <= 16'b1111111111111110;
        weights1[5689] <= 16'b1111111111111110;
        weights1[5690] <= 16'b0000000000000101;
        weights1[5691] <= 16'b0000000000000001;
        weights1[5692] <= 16'b1111111111111111;
        weights1[5693] <= 16'b1111111111101111;
        weights1[5694] <= 16'b1111111111111010;
        weights1[5695] <= 16'b0000000000001101;
        weights1[5696] <= 16'b1111111111111111;
        weights1[5697] <= 16'b1111111111111100;
        weights1[5698] <= 16'b1111111111110110;
        weights1[5699] <= 16'b1111111111111001;
        weights1[5700] <= 16'b1111111111111000;
        weights1[5701] <= 16'b0000000000000000;
        weights1[5702] <= 16'b0000000000000110;
        weights1[5703] <= 16'b1111111111111110;
        weights1[5704] <= 16'b0000000000010010;
        weights1[5705] <= 16'b0000000000001101;
        weights1[5706] <= 16'b0000000000001100;
        weights1[5707] <= 16'b1111111111110110;
        weights1[5708] <= 16'b1111111111111101;
        weights1[5709] <= 16'b0000000000001111;
        weights1[5710] <= 16'b1111111111101101;
        weights1[5711] <= 16'b1111111111111100;
        weights1[5712] <= 16'b1111111111111000;
        weights1[5713] <= 16'b1111111111110100;
        weights1[5714] <= 16'b1111111111111100;
        weights1[5715] <= 16'b1111111111111101;
        weights1[5716] <= 16'b1111111111110111;
        weights1[5717] <= 16'b1111111111111011;
        weights1[5718] <= 16'b0000000000000100;
        weights1[5719] <= 16'b0000000000000110;
        weights1[5720] <= 16'b1111111111110000;
        weights1[5721] <= 16'b1111111111111010;
        weights1[5722] <= 16'b1111111111111000;
        weights1[5723] <= 16'b1111111111110001;
        weights1[5724] <= 16'b0000000000000101;
        weights1[5725] <= 16'b1111111111111100;
        weights1[5726] <= 16'b0000000000010100;
        weights1[5727] <= 16'b0000000000001111;
        weights1[5728] <= 16'b0000000000010110;
        weights1[5729] <= 16'b0000000000100111;
        weights1[5730] <= 16'b0000000000001101;
        weights1[5731] <= 16'b0000000000001010;
        weights1[5732] <= 16'b0000000000000110;
        weights1[5733] <= 16'b0000000000100111;
        weights1[5734] <= 16'b0000000000010110;
        weights1[5735] <= 16'b0000000000010010;
        weights1[5736] <= 16'b0000000000011001;
        weights1[5737] <= 16'b0000000000001101;
        weights1[5738] <= 16'b0000000000000110;
        weights1[5739] <= 16'b0000000000110000;
        weights1[5740] <= 16'b1111111111110110;
        weights1[5741] <= 16'b0000000000000000;
        weights1[5742] <= 16'b1111111111111111;
        weights1[5743] <= 16'b1111111111110101;
        weights1[5744] <= 16'b1111111111111101;
        weights1[5745] <= 16'b0000000000000010;
        weights1[5746] <= 16'b1111111111110001;
        weights1[5747] <= 16'b1111111111111011;
        weights1[5748] <= 16'b1111111111111110;
        weights1[5749] <= 16'b0000000000000000;
        weights1[5750] <= 16'b1111111111111011;
        weights1[5751] <= 16'b1111111111110010;
        weights1[5752] <= 16'b1111111111111000;
        weights1[5753] <= 16'b1111111111111011;
        weights1[5754] <= 16'b0000000000000000;
        weights1[5755] <= 16'b0000000000011001;
        weights1[5756] <= 16'b0000000000000011;
        weights1[5757] <= 16'b0000000000001110;
        weights1[5758] <= 16'b0000000000000110;
        weights1[5759] <= 16'b0000000000011100;
        weights1[5760] <= 16'b0000000000000111;
        weights1[5761] <= 16'b0000000000100001;
        weights1[5762] <= 16'b1111111111111101;
        weights1[5763] <= 16'b0000000000100010;
        weights1[5764] <= 16'b0000000000111000;
        weights1[5765] <= 16'b0000000000101101;
        weights1[5766] <= 16'b0000000000011111;
        weights1[5767] <= 16'b0000000001000000;
        weights1[5768] <= 16'b1111111111101110;
        weights1[5769] <= 16'b0000000000000011;
        weights1[5770] <= 16'b1111111111110110;
        weights1[5771] <= 16'b1111111111110010;
        weights1[5772] <= 16'b1111111111110101;
        weights1[5773] <= 16'b0000000000010110;
        weights1[5774] <= 16'b1111111111111001;
        weights1[5775] <= 16'b0000000000001010;
        weights1[5776] <= 16'b1111111111110011;
        weights1[5777] <= 16'b0000000000000011;
        weights1[5778] <= 16'b1111111111110000;
        weights1[5779] <= 16'b0000000000001000;
        weights1[5780] <= 16'b1111111111101111;
        weights1[5781] <= 16'b1111111111111100;
        weights1[5782] <= 16'b0000000000000000;
        weights1[5783] <= 16'b0000000000010010;
        weights1[5784] <= 16'b0000000000001011;
        weights1[5785] <= 16'b0000000000001101;
        weights1[5786] <= 16'b0000000000100001;
        weights1[5787] <= 16'b0000000000100000;
        weights1[5788] <= 16'b0000000000001000;
        weights1[5789] <= 16'b1111111111111111;
        weights1[5790] <= 16'b1111111111101010;
        weights1[5791] <= 16'b0000000000100001;
        weights1[5792] <= 16'b0000000001011000;
        weights1[5793] <= 16'b0000000000111110;
        weights1[5794] <= 16'b0000000000110101;
        weights1[5795] <= 16'b0000000000110011;
        weights1[5796] <= 16'b1111111111110011;
        weights1[5797] <= 16'b1111111111110111;
        weights1[5798] <= 16'b0000000000000111;
        weights1[5799] <= 16'b1111111111111101;
        weights1[5800] <= 16'b1111111111110011;
        weights1[5801] <= 16'b0000000000000001;
        weights1[5802] <= 16'b0000000000001101;
        weights1[5803] <= 16'b1111111111110001;
        weights1[5804] <= 16'b0000000000001010;
        weights1[5805] <= 16'b0000000000000010;
        weights1[5806] <= 16'b1111111111111111;
        weights1[5807] <= 16'b1111111111100100;
        weights1[5808] <= 16'b1111111111100001;
        weights1[5809] <= 16'b1111111111111000;
        weights1[5810] <= 16'b1111111111110011;
        weights1[5811] <= 16'b0000000000001001;
        weights1[5812] <= 16'b0000000000011101;
        weights1[5813] <= 16'b0000000000100101;
        weights1[5814] <= 16'b0000000000110110;
        weights1[5815] <= 16'b0000000000110110;
        weights1[5816] <= 16'b0000000000111110;
        weights1[5817] <= 16'b0000000001010000;
        weights1[5818] <= 16'b0000000000110011;
        weights1[5819] <= 16'b0000000001010101;
        weights1[5820] <= 16'b0000000000111001;
        weights1[5821] <= 16'b0000000000111100;
        weights1[5822] <= 16'b0000000000101001;
        weights1[5823] <= 16'b0000000000010110;
        weights1[5824] <= 16'b1111111111111010;
        weights1[5825] <= 16'b1111111111110111;
        weights1[5826] <= 16'b0000000000001100;
        weights1[5827] <= 16'b1111111111111001;
        weights1[5828] <= 16'b1111111111110111;
        weights1[5829] <= 16'b0000000000001010;
        weights1[5830] <= 16'b0000000000000111;
        weights1[5831] <= 16'b0000000000001001;
        weights1[5832] <= 16'b0000000000010110;
        weights1[5833] <= 16'b0000000000010001;
        weights1[5834] <= 16'b0000000000001100;
        weights1[5835] <= 16'b1111111111111000;
        weights1[5836] <= 16'b1111111111101000;
        weights1[5837] <= 16'b1111111110110010;
        weights1[5838] <= 16'b1111111111001000;
        weights1[5839] <= 16'b1111111111110110;
        weights1[5840] <= 16'b0000000000000010;
        weights1[5841] <= 16'b0000000000011100;
        weights1[5842] <= 16'b0000000000101000;
        weights1[5843] <= 16'b0000000000101000;
        weights1[5844] <= 16'b0000000001001111;
        weights1[5845] <= 16'b0000000001001101;
        weights1[5846] <= 16'b0000000001011100;
        weights1[5847] <= 16'b0000000000100101;
        weights1[5848] <= 16'b0000000000111100;
        weights1[5849] <= 16'b0000000000110010;
        weights1[5850] <= 16'b0000000000010010;
        weights1[5851] <= 16'b0000000000010010;
        weights1[5852] <= 16'b0000000000000001;
        weights1[5853] <= 16'b1111111111111000;
        weights1[5854] <= 16'b0000000000000100;
        weights1[5855] <= 16'b0000000000001001;
        weights1[5856] <= 16'b1111111111111001;
        weights1[5857] <= 16'b1111111111111000;
        weights1[5858] <= 16'b0000000000000100;
        weights1[5859] <= 16'b0000000000000000;
        weights1[5860] <= 16'b0000000000010010;
        weights1[5861] <= 16'b0000000000000110;
        weights1[5862] <= 16'b0000000000010111;
        weights1[5863] <= 16'b0000000000100100;
        weights1[5864] <= 16'b1111111111101000;
        weights1[5865] <= 16'b1111111111000101;
        weights1[5866] <= 16'b1111111101111110;
        weights1[5867] <= 16'b1111111110001011;
        weights1[5868] <= 16'b1111111110011100;
        weights1[5869] <= 16'b1111111110101000;
        weights1[5870] <= 16'b1111111111011110;
        weights1[5871] <= 16'b1111111111101100;
        weights1[5872] <= 16'b1111111111111101;
        weights1[5873] <= 16'b0000000000001100;
        weights1[5874] <= 16'b1111111111111010;
        weights1[5875] <= 16'b0000000000001101;
        weights1[5876] <= 16'b1111111111110110;
        weights1[5877] <= 16'b0000000000000110;
        weights1[5878] <= 16'b1111111111101000;
        weights1[5879] <= 16'b1111111111101101;
        weights1[5880] <= 16'b0000000000001100;
        weights1[5881] <= 16'b0000000000000010;
        weights1[5882] <= 16'b0000000000000010;
        weights1[5883] <= 16'b0000000000001001;
        weights1[5884] <= 16'b1111111111110111;
        weights1[5885] <= 16'b1111111111110101;
        weights1[5886] <= 16'b1111111111110101;
        weights1[5887] <= 16'b0000000000000000;
        weights1[5888] <= 16'b0000000000001001;
        weights1[5889] <= 16'b0000000000000111;
        weights1[5890] <= 16'b0000000000000110;
        weights1[5891] <= 16'b0000000000010110;
        weights1[5892] <= 16'b0000000000011111;
        weights1[5893] <= 16'b0000000000000010;
        weights1[5894] <= 16'b1111111111010111;
        weights1[5895] <= 16'b1111111110001100;
        weights1[5896] <= 16'b1111111101001010;
        weights1[5897] <= 16'b1111111101001111;
        weights1[5898] <= 16'b1111111101000000;
        weights1[5899] <= 16'b1111111101110101;
        weights1[5900] <= 16'b1111111101101100;
        weights1[5901] <= 16'b1111111110011100;
        weights1[5902] <= 16'b1111111110100100;
        weights1[5903] <= 16'b1111111110101011;
        weights1[5904] <= 16'b1111111110110000;
        weights1[5905] <= 16'b1111111111001100;
        weights1[5906] <= 16'b1111111110111110;
        weights1[5907] <= 16'b1111111110111010;
        weights1[5908] <= 16'b0000000000001001;
        weights1[5909] <= 16'b0000000000010111;
        weights1[5910] <= 16'b0000000000010001;
        weights1[5911] <= 16'b1111111111111100;
        weights1[5912] <= 16'b1111111111111110;
        weights1[5913] <= 16'b1111111111111000;
        weights1[5914] <= 16'b0000000000001010;
        weights1[5915] <= 16'b0000000000001000;
        weights1[5916] <= 16'b0000000000000111;
        weights1[5917] <= 16'b0000000000000011;
        weights1[5918] <= 16'b0000000000001111;
        weights1[5919] <= 16'b0000000000011000;
        weights1[5920] <= 16'b0000000000000110;
        weights1[5921] <= 16'b0000000000010100;
        weights1[5922] <= 16'b0000000000101011;
        weights1[5923] <= 16'b1111111111100100;
        weights1[5924] <= 16'b1111111110011011;
        weights1[5925] <= 16'b1111111101101000;
        weights1[5926] <= 16'b1111111100101110;
        weights1[5927] <= 16'b1111111100010010;
        weights1[5928] <= 16'b1111111100111001;
        weights1[5929] <= 16'b1111111101110100;
        weights1[5930] <= 16'b1111111101100110;
        weights1[5931] <= 16'b1111111110100000;
        weights1[5932] <= 16'b1111111110100111;
        weights1[5933] <= 16'b1111111110110001;
        weights1[5934] <= 16'b1111111111000001;
        weights1[5935] <= 16'b1111111110101011;
        weights1[5936] <= 16'b0000000000001001;
        weights1[5937] <= 16'b0000000000001001;
        weights1[5938] <= 16'b0000000000001100;
        weights1[5939] <= 16'b1111111111111101;
        weights1[5940] <= 16'b0000000000000111;
        weights1[5941] <= 16'b1111111111101110;
        weights1[5942] <= 16'b1111111111111111;
        weights1[5943] <= 16'b0000000000001101;
        weights1[5944] <= 16'b0000000000001111;
        weights1[5945] <= 16'b0000000000000110;
        weights1[5946] <= 16'b1111111111110101;
        weights1[5947] <= 16'b1111111111111000;
        weights1[5948] <= 16'b0000000000010001;
        weights1[5949] <= 16'b0000000000001011;
        weights1[5950] <= 16'b0000000000001011;
        weights1[5951] <= 16'b0000000000001110;
        weights1[5952] <= 16'b1111111111111111;
        weights1[5953] <= 16'b1111111111011011;
        weights1[5954] <= 16'b1111111110011100;
        weights1[5955] <= 16'b1111111101001011;
        weights1[5956] <= 16'b1111111100110101;
        weights1[5957] <= 16'b1111111101100000;
        weights1[5958] <= 16'b1111111101111101;
        weights1[5959] <= 16'b1111111110010101;
        weights1[5960] <= 16'b1111111110110001;
        weights1[5961] <= 16'b1111111110110000;
        weights1[5962] <= 16'b1111111110111011;
        weights1[5963] <= 16'b1111111110110111;
        weights1[5964] <= 16'b0000000000000011;
        weights1[5965] <= 16'b1111111111111100;
        weights1[5966] <= 16'b0000000000000111;
        weights1[5967] <= 16'b0000000000001100;
        weights1[5968] <= 16'b0000000000001001;
        weights1[5969] <= 16'b0000000000001110;
        weights1[5970] <= 16'b1111111111110101;
        weights1[5971] <= 16'b0000000000000010;
        weights1[5972] <= 16'b1111111111111001;
        weights1[5973] <= 16'b0000000000000001;
        weights1[5974] <= 16'b1111111111111110;
        weights1[5975] <= 16'b0000000000001000;
        weights1[5976] <= 16'b1111111111110111;
        weights1[5977] <= 16'b1111111111111010;
        weights1[5978] <= 16'b0000000000010000;
        weights1[5979] <= 16'b0000000000011010;
        weights1[5980] <= 16'b0000000000001010;
        weights1[5981] <= 16'b0000000000010101;
        weights1[5982] <= 16'b0000000000100001;
        weights1[5983] <= 16'b1111111111000010;
        weights1[5984] <= 16'b1111111101101000;
        weights1[5985] <= 16'b1111111101110001;
        weights1[5986] <= 16'b1111111110000110;
        weights1[5987] <= 16'b1111111110010001;
        weights1[5988] <= 16'b1111111110011110;
        weights1[5989] <= 16'b1111111110111001;
        weights1[5990] <= 16'b1111111111000110;
        weights1[5991] <= 16'b1111111111001000;
        weights1[5992] <= 16'b1111111111111111;
        weights1[5993] <= 16'b0000000000000100;
        weights1[5994] <= 16'b0000000000001000;
        weights1[5995] <= 16'b0000000000010011;
        weights1[5996] <= 16'b0000000000001100;
        weights1[5997] <= 16'b1111111111111111;
        weights1[5998] <= 16'b0000000000000001;
        weights1[5999] <= 16'b1111111111100110;
        weights1[6000] <= 16'b0000000000000000;
        weights1[6001] <= 16'b1111111111110010;
        weights1[6002] <= 16'b0000000000000000;
        weights1[6003] <= 16'b1111111111111011;
        weights1[6004] <= 16'b0000000000010010;
        weights1[6005] <= 16'b1111111111111010;
        weights1[6006] <= 16'b0000000000010001;
        weights1[6007] <= 16'b0000000000010101;
        weights1[6008] <= 16'b0000000000011011;
        weights1[6009] <= 16'b0000000000001101;
        weights1[6010] <= 16'b0000000000100011;
        weights1[6011] <= 16'b0000000000010011;
        weights1[6012] <= 16'b1111111111001100;
        weights1[6013] <= 16'b1111111110001010;
        weights1[6014] <= 16'b1111111110000100;
        weights1[6015] <= 16'b1111111110011000;
        weights1[6016] <= 16'b1111111110101110;
        weights1[6017] <= 16'b1111111110111100;
        weights1[6018] <= 16'b1111111111001000;
        weights1[6019] <= 16'b1111111111000111;
        weights1[6020] <= 16'b1111111111110010;
        weights1[6021] <= 16'b0000000000010000;
        weights1[6022] <= 16'b1111111111111111;
        weights1[6023] <= 16'b0000000000000100;
        weights1[6024] <= 16'b1111111111111000;
        weights1[6025] <= 16'b0000000000010010;
        weights1[6026] <= 16'b0000000000000010;
        weights1[6027] <= 16'b0000000000010100;
        weights1[6028] <= 16'b1111111111111110;
        weights1[6029] <= 16'b0000000000000011;
        weights1[6030] <= 16'b1111111111111110;
        weights1[6031] <= 16'b1111111111101111;
        weights1[6032] <= 16'b0000000000000000;
        weights1[6033] <= 16'b0000000000001001;
        weights1[6034] <= 16'b0000000000000111;
        weights1[6035] <= 16'b0000000000001110;
        weights1[6036] <= 16'b0000000000011001;
        weights1[6037] <= 16'b0000000000001111;
        weights1[6038] <= 16'b0000000000100101;
        weights1[6039] <= 16'b0000000000101110;
        weights1[6040] <= 16'b1111111111111001;
        weights1[6041] <= 16'b1111111111000110;
        weights1[6042] <= 16'b1111111110100101;
        weights1[6043] <= 16'b1111111110100010;
        weights1[6044] <= 16'b1111111110110011;
        weights1[6045] <= 16'b1111111110111101;
        weights1[6046] <= 16'b1111111111001011;
        weights1[6047] <= 16'b1111111111010001;
        weights1[6048] <= 16'b1111111111111110;
        weights1[6049] <= 16'b0000000000001001;
        weights1[6050] <= 16'b0000000000000110;
        weights1[6051] <= 16'b1111111111111110;
        weights1[6052] <= 16'b1111111111110001;
        weights1[6053] <= 16'b1111111111111001;
        weights1[6054] <= 16'b0000000000001000;
        weights1[6055] <= 16'b1111111111111100;
        weights1[6056] <= 16'b0000000000000001;
        weights1[6057] <= 16'b1111111111110101;
        weights1[6058] <= 16'b1111111111111110;
        weights1[6059] <= 16'b0000000000000101;
        weights1[6060] <= 16'b0000000000000110;
        weights1[6061] <= 16'b0000000000010000;
        weights1[6062] <= 16'b0000000000001011;
        weights1[6063] <= 16'b0000000000001000;
        weights1[6064] <= 16'b0000000000101000;
        weights1[6065] <= 16'b0000000000000101;
        weights1[6066] <= 16'b0000000000010011;
        weights1[6067] <= 16'b0000000000101000;
        weights1[6068] <= 16'b0000000000001110;
        weights1[6069] <= 16'b1111111111100110;
        weights1[6070] <= 16'b1111111110111110;
        weights1[6071] <= 16'b1111111110111010;
        weights1[6072] <= 16'b1111111110111110;
        weights1[6073] <= 16'b1111111111001111;
        weights1[6074] <= 16'b1111111111001111;
        weights1[6075] <= 16'b1111111111010010;
        weights1[6076] <= 16'b1111111111111111;
        weights1[6077] <= 16'b1111111111111110;
        weights1[6078] <= 16'b0000000000001001;
        weights1[6079] <= 16'b0000000000000110;
        weights1[6080] <= 16'b1111111111111100;
        weights1[6081] <= 16'b1111111111110111;
        weights1[6082] <= 16'b0000000000001010;
        weights1[6083] <= 16'b0000000000001010;
        weights1[6084] <= 16'b0000000000000100;
        weights1[6085] <= 16'b1111111111111101;
        weights1[6086] <= 16'b1111111111111111;
        weights1[6087] <= 16'b0000000000000000;
        weights1[6088] <= 16'b1111111111101100;
        weights1[6089] <= 16'b1111111111111110;
        weights1[6090] <= 16'b1111111111111101;
        weights1[6091] <= 16'b0000000000001010;
        weights1[6092] <= 16'b0000000000011001;
        weights1[6093] <= 16'b0000000000011100;
        weights1[6094] <= 16'b0000000000000100;
        weights1[6095] <= 16'b0000000000010110;
        weights1[6096] <= 16'b0000000000000100;
        weights1[6097] <= 16'b1111111111110110;
        weights1[6098] <= 16'b1111111111100011;
        weights1[6099] <= 16'b1111111111001010;
        weights1[6100] <= 16'b1111111111001111;
        weights1[6101] <= 16'b1111111111010101;
        weights1[6102] <= 16'b1111111111010110;
        weights1[6103] <= 16'b1111111111011100;
        weights1[6104] <= 16'b1111111111111111;
        weights1[6105] <= 16'b0000000000000010;
        weights1[6106] <= 16'b0000000000000101;
        weights1[6107] <= 16'b0000000000000100;
        weights1[6108] <= 16'b0000000000001000;
        weights1[6109] <= 16'b0000000000001011;
        weights1[6110] <= 16'b1111111111111111;
        weights1[6111] <= 16'b0000000000001111;
        weights1[6112] <= 16'b0000000000000011;
        weights1[6113] <= 16'b0000000000001000;
        weights1[6114] <= 16'b0000000000001000;
        weights1[6115] <= 16'b0000000000000101;
        weights1[6116] <= 16'b0000000000000111;
        weights1[6117] <= 16'b0000000000000011;
        weights1[6118] <= 16'b0000000000000111;
        weights1[6119] <= 16'b1111111111110011;
        weights1[6120] <= 16'b1111111111111111;
        weights1[6121] <= 16'b0000000000011110;
        weights1[6122] <= 16'b0000000000100000;
        weights1[6123] <= 16'b0000000000100011;
        weights1[6124] <= 16'b0000000000010001;
        weights1[6125] <= 16'b0000000000011000;
        weights1[6126] <= 16'b1111111111100111;
        weights1[6127] <= 16'b1111111111001100;
        weights1[6128] <= 16'b1111111111011010;
        weights1[6129] <= 16'b1111111111010011;
        weights1[6130] <= 16'b1111111111100001;
        weights1[6131] <= 16'b1111111111100011;
        weights1[6132] <= 16'b0000000000000101;
        weights1[6133] <= 16'b0000000000001011;
        weights1[6134] <= 16'b0000000000001100;
        weights1[6135] <= 16'b0000000000011000;
        weights1[6136] <= 16'b0000000000000100;
        weights1[6137] <= 16'b0000000000000110;
        weights1[6138] <= 16'b0000000000001110;
        weights1[6139] <= 16'b0000000000011000;
        weights1[6140] <= 16'b0000000000001010;
        weights1[6141] <= 16'b0000000000001000;
        weights1[6142] <= 16'b0000000000001001;
        weights1[6143] <= 16'b0000000000010100;
        weights1[6144] <= 16'b0000000000010110;
        weights1[6145] <= 16'b0000000000000000;
        weights1[6146] <= 16'b1111111111111111;
        weights1[6147] <= 16'b0000000000010001;
        weights1[6148] <= 16'b0000000000001111;
        weights1[6149] <= 16'b0000000000000011;
        weights1[6150] <= 16'b0000000000010111;
        weights1[6151] <= 16'b0000000000100111;
        weights1[6152] <= 16'b0000000000100101;
        weights1[6153] <= 16'b1111111111111100;
        weights1[6154] <= 16'b1111111111100101;
        weights1[6155] <= 16'b1111111111011000;
        weights1[6156] <= 16'b1111111111001111;
        weights1[6157] <= 16'b1111111111011011;
        weights1[6158] <= 16'b1111111111100100;
        weights1[6159] <= 16'b1111111111101110;
        weights1[6160] <= 16'b1111111111111011;
        weights1[6161] <= 16'b1111111111111111;
        weights1[6162] <= 16'b1111111111111110;
        weights1[6163] <= 16'b0000000000010000;
        weights1[6164] <= 16'b0000000000011000;
        weights1[6165] <= 16'b1111111111111110;
        weights1[6166] <= 16'b1111111111111001;
        weights1[6167] <= 16'b1111111111111110;
        weights1[6168] <= 16'b1111111111111110;
        weights1[6169] <= 16'b0000000000001111;
        weights1[6170] <= 16'b0000000000001011;
        weights1[6171] <= 16'b0000000000001000;
        weights1[6172] <= 16'b0000000000010000;
        weights1[6173] <= 16'b0000000000011011;
        weights1[6174] <= 16'b0000000000011111;
        weights1[6175] <= 16'b0000000000000111;
        weights1[6176] <= 16'b0000000000011001;
        weights1[6177] <= 16'b0000000000010010;
        weights1[6178] <= 16'b0000000000100111;
        weights1[6179] <= 16'b0000000000100110;
        weights1[6180] <= 16'b0000000000011001;
        weights1[6181] <= 16'b1111111111111010;
        weights1[6182] <= 16'b1111111111101110;
        weights1[6183] <= 16'b1111111111011001;
        weights1[6184] <= 16'b1111111111011001;
        weights1[6185] <= 16'b1111111111100010;
        weights1[6186] <= 16'b1111111111110000;
        weights1[6187] <= 16'b1111111111111001;
        weights1[6188] <= 16'b0000000000000011;
        weights1[6189] <= 16'b1111111111111011;
        weights1[6190] <= 16'b1111111111110101;
        weights1[6191] <= 16'b0000000000010101;
        weights1[6192] <= 16'b0000000000001011;
        weights1[6193] <= 16'b0000000000000011;
        weights1[6194] <= 16'b0000000000000100;
        weights1[6195] <= 16'b0000000000001001;
        weights1[6196] <= 16'b0000000000000001;
        weights1[6197] <= 16'b0000000000001110;
        weights1[6198] <= 16'b0000000000000011;
        weights1[6199] <= 16'b0000000000010010;
        weights1[6200] <= 16'b0000000000000001;
        weights1[6201] <= 16'b0000000000000011;
        weights1[6202] <= 16'b0000000000000100;
        weights1[6203] <= 16'b0000000000010010;
        weights1[6204] <= 16'b0000000000000010;
        weights1[6205] <= 16'b0000000000001000;
        weights1[6206] <= 16'b0000000000010010;
        weights1[6207] <= 16'b0000000000100010;
        weights1[6208] <= 16'b0000000000010000;
        weights1[6209] <= 16'b1111111111111101;
        weights1[6210] <= 16'b1111111111110011;
        weights1[6211] <= 16'b1111111111101011;
        weights1[6212] <= 16'b1111111111100110;
        weights1[6213] <= 16'b1111111111110110;
        weights1[6214] <= 16'b1111111111111101;
        weights1[6215] <= 16'b1111111111111101;
        weights1[6216] <= 16'b0000000000000000;
        weights1[6217] <= 16'b0000000000000001;
        weights1[6218] <= 16'b0000000000000010;
        weights1[6219] <= 16'b0000000000000110;
        weights1[6220] <= 16'b0000000000000100;
        weights1[6221] <= 16'b0000000000001000;
        weights1[6222] <= 16'b1111111111110101;
        weights1[6223] <= 16'b0000000000000011;
        weights1[6224] <= 16'b1111111111111100;
        weights1[6225] <= 16'b0000000000000000;
        weights1[6226] <= 16'b0000000000000111;
        weights1[6227] <= 16'b1111111111111100;
        weights1[6228] <= 16'b0000000000001000;
        weights1[6229] <= 16'b0000000000010101;
        weights1[6230] <= 16'b1111111111111100;
        weights1[6231] <= 16'b0000000000011111;
        weights1[6232] <= 16'b0000000000001110;
        weights1[6233] <= 16'b0000000000100110;
        weights1[6234] <= 16'b0000000000010010;
        weights1[6235] <= 16'b0000000000001001;
        weights1[6236] <= 16'b0000000000010011;
        weights1[6237] <= 16'b1111111111111101;
        weights1[6238] <= 16'b0000000000000100;
        weights1[6239] <= 16'b1111111111110110;
        weights1[6240] <= 16'b1111111111111010;
        weights1[6241] <= 16'b1111111111111110;
        weights1[6242] <= 16'b1111111111111110;
        weights1[6243] <= 16'b1111111111111111;
        weights1[6244] <= 16'b0000000000000010;
        weights1[6245] <= 16'b0000000000001011;
        weights1[6246] <= 16'b0000000000001111;
        weights1[6247] <= 16'b0000000000001110;
        weights1[6248] <= 16'b0000000000001011;
        weights1[6249] <= 16'b0000000000001001;
        weights1[6250] <= 16'b0000000000001101;
        weights1[6251] <= 16'b0000000000011100;
        weights1[6252] <= 16'b0000000000011100;
        weights1[6253] <= 16'b0000000000010001;
        weights1[6254] <= 16'b0000000000101001;
        weights1[6255] <= 16'b0000000000101101;
        weights1[6256] <= 16'b0000000000101000;
        weights1[6257] <= 16'b0000000000011010;
        weights1[6258] <= 16'b0000000000100100;
        weights1[6259] <= 16'b0000000000100100;
        weights1[6260] <= 16'b0000000000110001;
        weights1[6261] <= 16'b0000000000011011;
        weights1[6262] <= 16'b0000000000010001;
        weights1[6263] <= 16'b0000000000000110;
        weights1[6264] <= 16'b0000000000010100;
        weights1[6265] <= 16'b0000000000001011;
        weights1[6266] <= 16'b1111111111111101;
        weights1[6267] <= 16'b1111111111111010;
        weights1[6268] <= 16'b0000000000000000;
        weights1[6269] <= 16'b0000000000000000;
        weights1[6270] <= 16'b1111111111111110;
        weights1[6271] <= 16'b0000000000000000;
        weights1[6272] <= 16'b0000000000000000;
        weights1[6273] <= 16'b1111111111111110;
        weights1[6274] <= 16'b1111111111111110;
        weights1[6275] <= 16'b1111111111111110;
        weights1[6276] <= 16'b1111111111111011;
        weights1[6277] <= 16'b1111111111111100;
        weights1[6278] <= 16'b0000000000000001;
        weights1[6279] <= 16'b0000000000000101;
        weights1[6280] <= 16'b0000000000000111;
        weights1[6281] <= 16'b0000000000001001;
        weights1[6282] <= 16'b0000000000010010;
        weights1[6283] <= 16'b0000000000000010;
        weights1[6284] <= 16'b0000000000001010;
        weights1[6285] <= 16'b0000000000010000;
        weights1[6286] <= 16'b0000000000011110;
        weights1[6287] <= 16'b0000000000010011;
        weights1[6288] <= 16'b0000000000001011;
        weights1[6289] <= 16'b0000000000010010;
        weights1[6290] <= 16'b0000000000001010;
        weights1[6291] <= 16'b0000000000001010;
        weights1[6292] <= 16'b0000000000000000;
        weights1[6293] <= 16'b0000000000000000;
        weights1[6294] <= 16'b1111111111111111;
        weights1[6295] <= 16'b0000000000000001;
        weights1[6296] <= 16'b0000000000000001;
        weights1[6297] <= 16'b1111111111111111;
        weights1[6298] <= 16'b0000000000000000;
        weights1[6299] <= 16'b0000000000000011;
        weights1[6300] <= 16'b1111111111111111;
        weights1[6301] <= 16'b1111111111111110;
        weights1[6302] <= 16'b1111111111111100;
        weights1[6303] <= 16'b1111111111111000;
        weights1[6304] <= 16'b1111111111110110;
        weights1[6305] <= 16'b1111111111110100;
        weights1[6306] <= 16'b1111111111111000;
        weights1[6307] <= 16'b1111111111111010;
        weights1[6308] <= 16'b0000000000000101;
        weights1[6309] <= 16'b0000000000000100;
        weights1[6310] <= 16'b0000000000001011;
        weights1[6311] <= 16'b0000000000010110;
        weights1[6312] <= 16'b0000000000100000;
        weights1[6313] <= 16'b0000000000010101;
        weights1[6314] <= 16'b0000000000001011;
        weights1[6315] <= 16'b0000000000001100;
        weights1[6316] <= 16'b0000000000010101;
        weights1[6317] <= 16'b0000000000001110;
        weights1[6318] <= 16'b0000000000010111;
        weights1[6319] <= 16'b0000000000001000;
        weights1[6320] <= 16'b0000000000000110;
        weights1[6321] <= 16'b0000000000001010;
        weights1[6322] <= 16'b0000000000010111;
        weights1[6323] <= 16'b0000000000001101;
        weights1[6324] <= 16'b0000000000001101;
        weights1[6325] <= 16'b0000000000001101;
        weights1[6326] <= 16'b0000000000000111;
        weights1[6327] <= 16'b0000000000000010;
        weights1[6328] <= 16'b1111111111111111;
        weights1[6329] <= 16'b1111111111111100;
        weights1[6330] <= 16'b1111111111111010;
        weights1[6331] <= 16'b1111111111110111;
        weights1[6332] <= 16'b1111111111110001;
        weights1[6333] <= 16'b1111111111101111;
        weights1[6334] <= 16'b1111111111110010;
        weights1[6335] <= 16'b0000000000000010;
        weights1[6336] <= 16'b1111111111111010;
        weights1[6337] <= 16'b0000000000000000;
        weights1[6338] <= 16'b1111111111111111;
        weights1[6339] <= 16'b0000000000001010;
        weights1[6340] <= 16'b0000000000000001;
        weights1[6341] <= 16'b0000000000000001;
        weights1[6342] <= 16'b0000000000000100;
        weights1[6343] <= 16'b1111111111111001;
        weights1[6344] <= 16'b0000000000010000;
        weights1[6345] <= 16'b0000000000001001;
        weights1[6346] <= 16'b0000000000000010;
        weights1[6347] <= 16'b0000000000001110;
        weights1[6348] <= 16'b0000000000000110;
        weights1[6349] <= 16'b0000000000010000;
        weights1[6350] <= 16'b0000000000011010;
        weights1[6351] <= 16'b1111111111111111;
        weights1[6352] <= 16'b0000000000000101;
        weights1[6353] <= 16'b0000000000001110;
        weights1[6354] <= 16'b0000000000001010;
        weights1[6355] <= 16'b0000000000001100;
        weights1[6356] <= 16'b1111111111111111;
        weights1[6357] <= 16'b1111111111111111;
        weights1[6358] <= 16'b1111111111111011;
        weights1[6359] <= 16'b1111111111110001;
        weights1[6360] <= 16'b1111111111101011;
        weights1[6361] <= 16'b1111111111110000;
        weights1[6362] <= 16'b1111111111110111;
        weights1[6363] <= 16'b1111111111111111;
        weights1[6364] <= 16'b0000000000001100;
        weights1[6365] <= 16'b1111111111110011;
        weights1[6366] <= 16'b0000000000001011;
        weights1[6367] <= 16'b1111111111111000;
        weights1[6368] <= 16'b1111111111111111;
        weights1[6369] <= 16'b0000000000001001;
        weights1[6370] <= 16'b1111111111110001;
        weights1[6371] <= 16'b1111111111101010;
        weights1[6372] <= 16'b1111111111111011;
        weights1[6373] <= 16'b1111111111111001;
        weights1[6374] <= 16'b1111111111111101;
        weights1[6375] <= 16'b0000000000000111;
        weights1[6376] <= 16'b0000000000001001;
        weights1[6377] <= 16'b0000000000010001;
        weights1[6378] <= 16'b0000000000010110;
        weights1[6379] <= 16'b0000000000010101;
        weights1[6380] <= 16'b0000000000010111;
        weights1[6381] <= 16'b0000000000001010;
        weights1[6382] <= 16'b0000000000010000;
        weights1[6383] <= 16'b0000000000010000;
        weights1[6384] <= 16'b1111111111111011;
        weights1[6385] <= 16'b1111111111111001;
        weights1[6386] <= 16'b1111111111111000;
        weights1[6387] <= 16'b1111111111110010;
        weights1[6388] <= 16'b1111111111101100;
        weights1[6389] <= 16'b1111111111101001;
        weights1[6390] <= 16'b1111111111110110;
        weights1[6391] <= 16'b0000000000000011;
        weights1[6392] <= 16'b1111111111110010;
        weights1[6393] <= 16'b0000000000010010;
        weights1[6394] <= 16'b0000000000010110;
        weights1[6395] <= 16'b1111111111110101;
        weights1[6396] <= 16'b0000000000001111;
        weights1[6397] <= 16'b0000000000000110;
        weights1[6398] <= 16'b1111111111111000;
        weights1[6399] <= 16'b0000000000010001;
        weights1[6400] <= 16'b0000000000001100;
        weights1[6401] <= 16'b1111111111111010;
        weights1[6402] <= 16'b1111111111101111;
        weights1[6403] <= 16'b1111111111111011;
        weights1[6404] <= 16'b0000000000001101;
        weights1[6405] <= 16'b1111111111111001;
        weights1[6406] <= 16'b1111111111111100;
        weights1[6407] <= 16'b0000000000000111;
        weights1[6408] <= 16'b1111111111111000;
        weights1[6409] <= 16'b0000000000001000;
        weights1[6410] <= 16'b0000000000010000;
        weights1[6411] <= 16'b0000000000001011;
        weights1[6412] <= 16'b1111111111111100;
        weights1[6413] <= 16'b1111111111111000;
        weights1[6414] <= 16'b1111111111111010;
        weights1[6415] <= 16'b1111111111111100;
        weights1[6416] <= 16'b1111111111110111;
        weights1[6417] <= 16'b1111111111100101;
        weights1[6418] <= 16'b1111111111101101;
        weights1[6419] <= 16'b0000000000000101;
        weights1[6420] <= 16'b1111111111101110;
        weights1[6421] <= 16'b0000000000001001;
        weights1[6422] <= 16'b0000000000000110;
        weights1[6423] <= 16'b0000000000000100;
        weights1[6424] <= 16'b0000000000001010;
        weights1[6425] <= 16'b1111111111101011;
        weights1[6426] <= 16'b0000000000001110;
        weights1[6427] <= 16'b1111111111111001;
        weights1[6428] <= 16'b0000000000011101;
        weights1[6429] <= 16'b0000000000001110;
        weights1[6430] <= 16'b0000000000011101;
        weights1[6431] <= 16'b0000000000001001;
        weights1[6432] <= 16'b0000000000010111;
        weights1[6433] <= 16'b0000000000010110;
        weights1[6434] <= 16'b0000000000001010;
        weights1[6435] <= 16'b1111111111110110;
        weights1[6436] <= 16'b0000000000000111;
        weights1[6437] <= 16'b0000000000100001;
        weights1[6438] <= 16'b0000000000001110;
        weights1[6439] <= 16'b0000000000010001;
        weights1[6440] <= 16'b1111111111111001;
        weights1[6441] <= 16'b1111111111110000;
        weights1[6442] <= 16'b1111111111110001;
        weights1[6443] <= 16'b1111111111110110;
        weights1[6444] <= 16'b1111111111111000;
        weights1[6445] <= 16'b1111111111101000;
        weights1[6446] <= 16'b1111111111101010;
        weights1[6447] <= 16'b1111111111100101;
        weights1[6448] <= 16'b1111111111110001;
        weights1[6449] <= 16'b0000000000011001;
        weights1[6450] <= 16'b1111111111101111;
        weights1[6451] <= 16'b1111111111111110;
        weights1[6452] <= 16'b0000000000001110;
        weights1[6453] <= 16'b0000000000000010;
        weights1[6454] <= 16'b1111111111111100;
        weights1[6455] <= 16'b0000000000010000;
        weights1[6456] <= 16'b1111111111111001;
        weights1[6457] <= 16'b1111111111111010;
        weights1[6458] <= 16'b0000000000010111;
        weights1[6459] <= 16'b0000000000001010;
        weights1[6460] <= 16'b0000000000000000;
        weights1[6461] <= 16'b0000000000011000;
        weights1[6462] <= 16'b1111111111110000;
        weights1[6463] <= 16'b0000000000000110;
        weights1[6464] <= 16'b0000000000011111;
        weights1[6465] <= 16'b0000000000011001;
        weights1[6466] <= 16'b0000000000010110;
        weights1[6467] <= 16'b1111111111111111;
        weights1[6468] <= 16'b1111111111110101;
        weights1[6469] <= 16'b1111111111110100;
        weights1[6470] <= 16'b1111111111111111;
        weights1[6471] <= 16'b1111111111111010;
        weights1[6472] <= 16'b0000000000000011;
        weights1[6473] <= 16'b1111111111101101;
        weights1[6474] <= 16'b1111111111100101;
        weights1[6475] <= 16'b1111111111110011;
        weights1[6476] <= 16'b0000000000000000;
        weights1[6477] <= 16'b1111111111111000;
        weights1[6478] <= 16'b0000000000001111;
        weights1[6479] <= 16'b0000000000000110;
        weights1[6480] <= 16'b1111111111111100;
        weights1[6481] <= 16'b0000000000001000;
        weights1[6482] <= 16'b1111111111110001;
        weights1[6483] <= 16'b0000000000000001;
        weights1[6484] <= 16'b0000000000001001;
        weights1[6485] <= 16'b0000000000000110;
        weights1[6486] <= 16'b0000000000000110;
        weights1[6487] <= 16'b1111111111101110;
        weights1[6488] <= 16'b0000000000000011;
        weights1[6489] <= 16'b1111111111101101;
        weights1[6490] <= 16'b0000000000100000;
        weights1[6491] <= 16'b0000000000001110;
        weights1[6492] <= 16'b0000000000000000;
        weights1[6493] <= 16'b0000000000000110;
        weights1[6494] <= 16'b0000000000001100;
        weights1[6495] <= 16'b0000000000000011;
        weights1[6496] <= 16'b1111111111111010;
        weights1[6497] <= 16'b1111111111111011;
        weights1[6498] <= 16'b1111111111111110;
        weights1[6499] <= 16'b1111111111110011;
        weights1[6500] <= 16'b1111111111111111;
        weights1[6501] <= 16'b1111111111100110;
        weights1[6502] <= 16'b0000000000000010;
        weights1[6503] <= 16'b1111111111101000;
        weights1[6504] <= 16'b1111111111101111;
        weights1[6505] <= 16'b1111111111110010;
        weights1[6506] <= 16'b1111111111111010;
        weights1[6507] <= 16'b0000000000001111;
        weights1[6508] <= 16'b0000000000001001;
        weights1[6509] <= 16'b0000000000010011;
        weights1[6510] <= 16'b0000000000001110;
        weights1[6511] <= 16'b0000000000000100;
        weights1[6512] <= 16'b0000000000000111;
        weights1[6513] <= 16'b0000000000000110;
        weights1[6514] <= 16'b1111111111111110;
        weights1[6515] <= 16'b0000000000010001;
        weights1[6516] <= 16'b0000000000010001;
        weights1[6517] <= 16'b0000000000010010;
        weights1[6518] <= 16'b0000000000000110;
        weights1[6519] <= 16'b0000000000001001;
        weights1[6520] <= 16'b0000000000100010;
        weights1[6521] <= 16'b0000000000000000;
        weights1[6522] <= 16'b1111111111111000;
        weights1[6523] <= 16'b1111111111111000;
        weights1[6524] <= 16'b1111111111111101;
        weights1[6525] <= 16'b0000000000000010;
        weights1[6526] <= 16'b0000000000001000;
        weights1[6527] <= 16'b1111111111110110;
        weights1[6528] <= 16'b1111111111110001;
        weights1[6529] <= 16'b0000000000000110;
        weights1[6530] <= 16'b0000000000000010;
        weights1[6531] <= 16'b0000000000001000;
        weights1[6532] <= 16'b0000000000000010;
        weights1[6533] <= 16'b1111111111111001;
        weights1[6534] <= 16'b1111111111110110;
        weights1[6535] <= 16'b1111111111111110;
        weights1[6536] <= 16'b1111111111110111;
        weights1[6537] <= 16'b1111111111101110;
        weights1[6538] <= 16'b1111111111110011;
        weights1[6539] <= 16'b1111111111101111;
        weights1[6540] <= 16'b1111111111011110;
        weights1[6541] <= 16'b0000000000000101;
        weights1[6542] <= 16'b1111111111110000;
        weights1[6543] <= 16'b1111111111110111;
        weights1[6544] <= 16'b1111111111110111;
        weights1[6545] <= 16'b0000000000010000;
        weights1[6546] <= 16'b0000000000100010;
        weights1[6547] <= 16'b0000000000100101;
        weights1[6548] <= 16'b0000000000010011;
        weights1[6549] <= 16'b0000000000000001;
        weights1[6550] <= 16'b1111111111111000;
        weights1[6551] <= 16'b1111111111011010;
        weights1[6552] <= 16'b1111111111110100;
        weights1[6553] <= 16'b0000000000000101;
        weights1[6554] <= 16'b1111111111111100;
        weights1[6555] <= 16'b1111111111101110;
        weights1[6556] <= 16'b0000000000000111;
        weights1[6557] <= 16'b0000000000011011;
        weights1[6558] <= 16'b0000000000001010;
        weights1[6559] <= 16'b1111111111110011;
        weights1[6560] <= 16'b0000000000001101;
        weights1[6561] <= 16'b0000000000010001;
        weights1[6562] <= 16'b1111111111111010;
        weights1[6563] <= 16'b1111111111110011;
        weights1[6564] <= 16'b1111111111111101;
        weights1[6565] <= 16'b1111111111100110;
        weights1[6566] <= 16'b1111111111011011;
        weights1[6567] <= 16'b1111111111011100;
        weights1[6568] <= 16'b1111111111111101;
        weights1[6569] <= 16'b1111111111100011;
        weights1[6570] <= 16'b0000000000000111;
        weights1[6571] <= 16'b1111111111111011;
        weights1[6572] <= 16'b1111111111110001;
        weights1[6573] <= 16'b1111111111111110;
        weights1[6574] <= 16'b0000000000010101;
        weights1[6575] <= 16'b0000000000101100;
        weights1[6576] <= 16'b1111111111110011;
        weights1[6577] <= 16'b1111111111101111;
        weights1[6578] <= 16'b1111111111001100;
        weights1[6579] <= 16'b1111111111000010;
        weights1[6580] <= 16'b1111111111110011;
        weights1[6581] <= 16'b1111111111110111;
        weights1[6582] <= 16'b1111111111111000;
        weights1[6583] <= 16'b1111111111101110;
        weights1[6584] <= 16'b0000000000010111;
        weights1[6585] <= 16'b0000000000100010;
        weights1[6586] <= 16'b0000000000010110;
        weights1[6587] <= 16'b0000000000001100;
        weights1[6588] <= 16'b1111111111110000;
        weights1[6589] <= 16'b1111111111100011;
        weights1[6590] <= 16'b1111111111110010;
        weights1[6591] <= 16'b1111111111110000;
        weights1[6592] <= 16'b1111111111110110;
        weights1[6593] <= 16'b1111111111110010;
        weights1[6594] <= 16'b0000000000000110;
        weights1[6595] <= 16'b1111111111010011;
        weights1[6596] <= 16'b1111111111011001;
        weights1[6597] <= 16'b1111111111100000;
        weights1[6598] <= 16'b1111111111110111;
        weights1[6599] <= 16'b1111111111111101;
        weights1[6600] <= 16'b0000000000000010;
        weights1[6601] <= 16'b0000000000001100;
        weights1[6602] <= 16'b0000000000100010;
        weights1[6603] <= 16'b1111111111110111;
        weights1[6604] <= 16'b1111111111000010;
        weights1[6605] <= 16'b1111111111000101;
        weights1[6606] <= 16'b1111111110110110;
        weights1[6607] <= 16'b1111111110111100;
        weights1[6608] <= 16'b1111111111111100;
        weights1[6609] <= 16'b1111111111110010;
        weights1[6610] <= 16'b1111111111110010;
        weights1[6611] <= 16'b1111111111111101;
        weights1[6612] <= 16'b0000000000010001;
        weights1[6613] <= 16'b0000000000000101;
        weights1[6614] <= 16'b1111111111100001;
        weights1[6615] <= 16'b0000000000000001;
        weights1[6616] <= 16'b1111111111111011;
        weights1[6617] <= 16'b1111111111100001;
        weights1[6618] <= 16'b1111111111100111;
        weights1[6619] <= 16'b1111111111111010;
        weights1[6620] <= 16'b1111111111100101;
        weights1[6621] <= 16'b0000000000001101;
        weights1[6622] <= 16'b0000000000000010;
        weights1[6623] <= 16'b1111111111101000;
        weights1[6624] <= 16'b1111111111100001;
        weights1[6625] <= 16'b1111111111001101;
        weights1[6626] <= 16'b1111111111011101;
        weights1[6627] <= 16'b1111111111100100;
        weights1[6628] <= 16'b1111111111100100;
        weights1[6629] <= 16'b1111111111101001;
        weights1[6630] <= 16'b1111111111000010;
        weights1[6631] <= 16'b1111111110001101;
        weights1[6632] <= 16'b1111111110001000;
        weights1[6633] <= 16'b1111111110010111;
        weights1[6634] <= 16'b1111111110111000;
        weights1[6635] <= 16'b1111111110110101;
        weights1[6636] <= 16'b1111111111110010;
        weights1[6637] <= 16'b1111111111110001;
        weights1[6638] <= 16'b1111111111110001;
        weights1[6639] <= 16'b1111111111110100;
        weights1[6640] <= 16'b1111111111011000;
        weights1[6641] <= 16'b1111111111011010;
        weights1[6642] <= 16'b1111111111011111;
        weights1[6643] <= 16'b1111111111011001;
        weights1[6644] <= 16'b1111111111011001;
        weights1[6645] <= 16'b1111111111111010;
        weights1[6646] <= 16'b1111111111100001;
        weights1[6647] <= 16'b1111111111100110;
        weights1[6648] <= 16'b0000000000011111;
        weights1[6649] <= 16'b0000000000010111;
        weights1[6650] <= 16'b0000000000101111;
        weights1[6651] <= 16'b0000000000000001;
        weights1[6652] <= 16'b1111111111011000;
        weights1[6653] <= 16'b1111111111100101;
        weights1[6654] <= 16'b1111111111011000;
        weights1[6655] <= 16'b1111111111001101;
        weights1[6656] <= 16'b1111111110100010;
        weights1[6657] <= 16'b1111111101110000;
        weights1[6658] <= 16'b1111111101011010;
        weights1[6659] <= 16'b1111111101101010;
        weights1[6660] <= 16'b1111111101111001;
        weights1[6661] <= 16'b1111111110011111;
        weights1[6662] <= 16'b1111111110110000;
        weights1[6663] <= 16'b1111111110110111;
        weights1[6664] <= 16'b1111111111101101;
        weights1[6665] <= 16'b1111111111101101;
        weights1[6666] <= 16'b1111111111100001;
        weights1[6667] <= 16'b1111111111011100;
        weights1[6668] <= 16'b1111111111010100;
        weights1[6669] <= 16'b1111111110111110;
        weights1[6670] <= 16'b1111111111011011;
        weights1[6671] <= 16'b1111111111011000;
        weights1[6672] <= 16'b1111111111010111;
        weights1[6673] <= 16'b1111111111011101;
        weights1[6674] <= 16'b1111111111101111;
        weights1[6675] <= 16'b0000000000010011;
        weights1[6676] <= 16'b0000000000100101;
        weights1[6677] <= 16'b0000000000100100;
        weights1[6678] <= 16'b0000000000001101;
        weights1[6679] <= 16'b0000000000100011;
        weights1[6680] <= 16'b0000000000001000;
        weights1[6681] <= 16'b1111111111111000;
        weights1[6682] <= 16'b1111111111100110;
        weights1[6683] <= 16'b1111111111011100;
        weights1[6684] <= 16'b1111111110110000;
        weights1[6685] <= 16'b1111111110010011;
        weights1[6686] <= 16'b1111111101011001;
        weights1[6687] <= 16'b1111111101100100;
        weights1[6688] <= 16'b1111111101111011;
        weights1[6689] <= 16'b1111111110010101;
        weights1[6690] <= 16'b1111111110100101;
        weights1[6691] <= 16'b1111111110101111;
        weights1[6692] <= 16'b1111111111101111;
        weights1[6693] <= 16'b1111111111101001;
        weights1[6694] <= 16'b1111111111010110;
        weights1[6695] <= 16'b1111111111001100;
        weights1[6696] <= 16'b1111111111000110;
        weights1[6697] <= 16'b1111111111001101;
        weights1[6698] <= 16'b1111111110111101;
        weights1[6699] <= 16'b1111111111110011;
        weights1[6700] <= 16'b1111111111110000;
        weights1[6701] <= 16'b0000000000000000;
        weights1[6702] <= 16'b0000000000000100;
        weights1[6703] <= 16'b0000000000000010;
        weights1[6704] <= 16'b0000000000001111;
        weights1[6705] <= 16'b0000000000101000;
        weights1[6706] <= 16'b0000000000101010;
        weights1[6707] <= 16'b0000000000011100;
        weights1[6708] <= 16'b0000000000011011;
        weights1[6709] <= 16'b0000000000000000;
        weights1[6710] <= 16'b1111111111110110;
        weights1[6711] <= 16'b1111111111110100;
        weights1[6712] <= 16'b1111111111011101;
        weights1[6713] <= 16'b1111111111000010;
        weights1[6714] <= 16'b1111111110111111;
        weights1[6715] <= 16'b1111111110100000;
        weights1[6716] <= 16'b1111111110010100;
        weights1[6717] <= 16'b1111111110010011;
        weights1[6718] <= 16'b1111111110100101;
        weights1[6719] <= 16'b1111111110110000;
        weights1[6720] <= 16'b1111111111101110;
        weights1[6721] <= 16'b1111111111100110;
        weights1[6722] <= 16'b1111111111001110;
        weights1[6723] <= 16'b1111111111000011;
        weights1[6724] <= 16'b1111111111001001;
        weights1[6725] <= 16'b1111111111011011;
        weights1[6726] <= 16'b1111111111110101;
        weights1[6727] <= 16'b0000000000001010;
        weights1[6728] <= 16'b0000000000000011;
        weights1[6729] <= 16'b0000000000010010;
        weights1[6730] <= 16'b0000000000011101;
        weights1[6731] <= 16'b0000000000001010;
        weights1[6732] <= 16'b0000000000001110;
        weights1[6733] <= 16'b1111111111111111;
        weights1[6734] <= 16'b0000000000100100;
        weights1[6735] <= 16'b0000000000101001;
        weights1[6736] <= 16'b1111111111111101;
        weights1[6737] <= 16'b1111111111111100;
        weights1[6738] <= 16'b1111111111100110;
        weights1[6739] <= 16'b0000000000000000;
        weights1[6740] <= 16'b1111111111110010;
        weights1[6741] <= 16'b1111111111110011;
        weights1[6742] <= 16'b1111111111110010;
        weights1[6743] <= 16'b1111111111011110;
        weights1[6744] <= 16'b1111111111001010;
        weights1[6745] <= 16'b1111111110110010;
        weights1[6746] <= 16'b1111111110101101;
        weights1[6747] <= 16'b1111111111000100;
        weights1[6748] <= 16'b1111111111101111;
        weights1[6749] <= 16'b1111111111100101;
        weights1[6750] <= 16'b1111111111010011;
        weights1[6751] <= 16'b1111111111011010;
        weights1[6752] <= 16'b1111111111100101;
        weights1[6753] <= 16'b0000000000000001;
        weights1[6754] <= 16'b0000000000010010;
        weights1[6755] <= 16'b0000000000000110;
        weights1[6756] <= 16'b0000000000001110;
        weights1[6757] <= 16'b0000000000010011;
        weights1[6758] <= 16'b1111111111111101;
        weights1[6759] <= 16'b1111111111110101;
        weights1[6760] <= 16'b0000000000100001;
        weights1[6761] <= 16'b0000000000001010;
        weights1[6762] <= 16'b1111111111111101;
        weights1[6763] <= 16'b1111111111111111;
        weights1[6764] <= 16'b0000000000010011;
        weights1[6765] <= 16'b1111111111111000;
        weights1[6766] <= 16'b0000000000000111;
        weights1[6767] <= 16'b0000000000001011;
        weights1[6768] <= 16'b0000000000011100;
        weights1[6769] <= 16'b0000000000011011;
        weights1[6770] <= 16'b0000000000010111;
        weights1[6771] <= 16'b1111111111110011;
        weights1[6772] <= 16'b1111111111101111;
        weights1[6773] <= 16'b1111111111100000;
        weights1[6774] <= 16'b1111111111001100;
        weights1[6775] <= 16'b1111111111011100;
        weights1[6776] <= 16'b1111111111110010;
        weights1[6777] <= 16'b1111111111100010;
        weights1[6778] <= 16'b1111111111100010;
        weights1[6779] <= 16'b1111111111101111;
        weights1[6780] <= 16'b0000000000001101;
        weights1[6781] <= 16'b0000000000011001;
        weights1[6782] <= 16'b0000000000011101;
        weights1[6783] <= 16'b0000000000010100;
        weights1[6784] <= 16'b1111111111111101;
        weights1[6785] <= 16'b0000000000011110;
        weights1[6786] <= 16'b0000000000000110;
        weights1[6787] <= 16'b0000000000000110;
        weights1[6788] <= 16'b0000000000001111;
        weights1[6789] <= 16'b0000000000001100;
        weights1[6790] <= 16'b1111111111110011;
        weights1[6791] <= 16'b0000000000000110;
        weights1[6792] <= 16'b0000000000010110;
        weights1[6793] <= 16'b0000000000010010;
        weights1[6794] <= 16'b0000000000010001;
        weights1[6795] <= 16'b0000000000100010;
        weights1[6796] <= 16'b0000000000101001;
        weights1[6797] <= 16'b0000000000011000;
        weights1[6798] <= 16'b0000000000110000;
        weights1[6799] <= 16'b0000000000011100;
        weights1[6800] <= 16'b0000000000010010;
        weights1[6801] <= 16'b0000000000000100;
        weights1[6802] <= 16'b1111111111110000;
        weights1[6803] <= 16'b1111111111111011;
        weights1[6804] <= 16'b1111111111111011;
        weights1[6805] <= 16'b1111111111111100;
        weights1[6806] <= 16'b1111111111110111;
        weights1[6807] <= 16'b0000000000000101;
        weights1[6808] <= 16'b0000000000001011;
        weights1[6809] <= 16'b0000000000000011;
        weights1[6810] <= 16'b0000000000001001;
        weights1[6811] <= 16'b0000000000001011;
        weights1[6812] <= 16'b0000000000000001;
        weights1[6813] <= 16'b0000000000000101;
        weights1[6814] <= 16'b0000000000011001;
        weights1[6815] <= 16'b0000000000000000;
        weights1[6816] <= 16'b1111111111111101;
        weights1[6817] <= 16'b0000000000001010;
        weights1[6818] <= 16'b0000000000000001;
        weights1[6819] <= 16'b0000000000010110;
        weights1[6820] <= 16'b0000000000000010;
        weights1[6821] <= 16'b0000000000010110;
        weights1[6822] <= 16'b0000000000001001;
        weights1[6823] <= 16'b0000000000011101;
        weights1[6824] <= 16'b0000000000011101;
        weights1[6825] <= 16'b0000000001000001;
        weights1[6826] <= 16'b0000000001000110;
        weights1[6827] <= 16'b0000000001010101;
        weights1[6828] <= 16'b0000000000100001;
        weights1[6829] <= 16'b0000000000100110;
        weights1[6830] <= 16'b0000000000100011;
        weights1[6831] <= 16'b0000000000010101;
        weights1[6832] <= 16'b0000000000001011;
        weights1[6833] <= 16'b0000000000000111;
        weights1[6834] <= 16'b0000000000001100;
        weights1[6835] <= 16'b0000000000000011;
        weights1[6836] <= 16'b1111111111111101;
        weights1[6837] <= 16'b0000000000110101;
        weights1[6838] <= 16'b0000000000011010;
        weights1[6839] <= 16'b0000000000011101;
        weights1[6840] <= 16'b0000000000001100;
        weights1[6841] <= 16'b0000000000000010;
        weights1[6842] <= 16'b0000000000011010;
        weights1[6843] <= 16'b0000000000001010;
        weights1[6844] <= 16'b1111111111111010;
        weights1[6845] <= 16'b0000000000010011;
        weights1[6846] <= 16'b0000000000000001;
        weights1[6847] <= 16'b0000000000001001;
        weights1[6848] <= 16'b0000000000010011;
        weights1[6849] <= 16'b0000000000011011;
        weights1[6850] <= 16'b0000000000110110;
        weights1[6851] <= 16'b0000000000001110;
        weights1[6852] <= 16'b0000000000111001;
        weights1[6853] <= 16'b0000000000101110;
        weights1[6854] <= 16'b0000000000111000;
        weights1[6855] <= 16'b0000000001100001;
        weights1[6856] <= 16'b0000000000110110;
        weights1[6857] <= 16'b0000000000110111;
        weights1[6858] <= 16'b0000000000110100;
        weights1[6859] <= 16'b0000000000011010;
        weights1[6860] <= 16'b0000000000010001;
        weights1[6861] <= 16'b0000000000010101;
        weights1[6862] <= 16'b0000000000010010;
        weights1[6863] <= 16'b1111111111110110;
        weights1[6864] <= 16'b1111111111110111;
        weights1[6865] <= 16'b0000000000011011;
        weights1[6866] <= 16'b0000000000001010;
        weights1[6867] <= 16'b0000000000001001;
        weights1[6868] <= 16'b0000000000010001;
        weights1[6869] <= 16'b0000000000011000;
        weights1[6870] <= 16'b1111111111111010;
        weights1[6871] <= 16'b0000000000001011;
        weights1[6872] <= 16'b0000000000010100;
        weights1[6873] <= 16'b0000000000100111;
        weights1[6874] <= 16'b0000000000011100;
        weights1[6875] <= 16'b0000000000000111;
        weights1[6876] <= 16'b0000000000001110;
        weights1[6877] <= 16'b0000000000010111;
        weights1[6878] <= 16'b0000000000100110;
        weights1[6879] <= 16'b0000000000101101;
        weights1[6880] <= 16'b0000000000110100;
        weights1[6881] <= 16'b0000000000110011;
        weights1[6882] <= 16'b0000000000111000;
        weights1[6883] <= 16'b0000000001001100;
        weights1[6884] <= 16'b0000000000110111;
        weights1[6885] <= 16'b0000000001000110;
        weights1[6886] <= 16'b0000000000101110;
        weights1[6887] <= 16'b0000000000011100;
        weights1[6888] <= 16'b0000000000001101;
        weights1[6889] <= 16'b0000000000010001;
        weights1[6890] <= 16'b0000000000001010;
        weights1[6891] <= 16'b1111111111111011;
        weights1[6892] <= 16'b0000000000000111;
        weights1[6893] <= 16'b0000000000001101;
        weights1[6894] <= 16'b1111111111110111;
        weights1[6895] <= 16'b0000000000001100;
        weights1[6896] <= 16'b0000000000000010;
        weights1[6897] <= 16'b0000000000010100;
        weights1[6898] <= 16'b0000000000000010;
        weights1[6899] <= 16'b0000000000011111;
        weights1[6900] <= 16'b0000000000000110;
        weights1[6901] <= 16'b1111111111111110;
        weights1[6902] <= 16'b1111111111111101;
        weights1[6903] <= 16'b0000000000011001;
        weights1[6904] <= 16'b1111111111111000;
        weights1[6905] <= 16'b0000000000001110;
        weights1[6906] <= 16'b0000000000010101;
        weights1[6907] <= 16'b0000000000101010;
        weights1[6908] <= 16'b0000000000001111;
        weights1[6909] <= 16'b0000000000100100;
        weights1[6910] <= 16'b0000000000001111;
        weights1[6911] <= 16'b0000000000100010;
        weights1[6912] <= 16'b0000000000101111;
        weights1[6913] <= 16'b0000000000101110;
        weights1[6914] <= 16'b0000000000100010;
        weights1[6915] <= 16'b0000000000010100;
        weights1[6916] <= 16'b0000000000010001;
        weights1[6917] <= 16'b0000000000010110;
        weights1[6918] <= 16'b0000000000000111;
        weights1[6919] <= 16'b0000000000000010;
        weights1[6920] <= 16'b0000000000000111;
        weights1[6921] <= 16'b0000000000010101;
        weights1[6922] <= 16'b0000000000000001;
        weights1[6923] <= 16'b0000000000001100;
        weights1[6924] <= 16'b0000000000001100;
        weights1[6925] <= 16'b0000000000010000;
        weights1[6926] <= 16'b0000000000000110;
        weights1[6927] <= 16'b0000000000010111;
        weights1[6928] <= 16'b0000000000011000;
        weights1[6929] <= 16'b0000000000101011;
        weights1[6930] <= 16'b0000000000001010;
        weights1[6931] <= 16'b0000000000101001;
        weights1[6932] <= 16'b0000000000100000;
        weights1[6933] <= 16'b1111111111111110;
        weights1[6934] <= 16'b0000000000000010;
        weights1[6935] <= 16'b0000000000001001;
        weights1[6936] <= 16'b0000000000100111;
        weights1[6937] <= 16'b1111111111101011;
        weights1[6938] <= 16'b0000000000001100;
        weights1[6939] <= 16'b0000000000010000;
        weights1[6940] <= 16'b0000000000010010;
        weights1[6941] <= 16'b0000000000011010;
        weights1[6942] <= 16'b0000000000010001;
        weights1[6943] <= 16'b0000000000001010;
        weights1[6944] <= 16'b0000000000000110;
        weights1[6945] <= 16'b0000000000000100;
        weights1[6946] <= 16'b0000000000000011;
        weights1[6947] <= 16'b1111111111111100;
        weights1[6948] <= 16'b0000000000000101;
        weights1[6949] <= 16'b0000000000000010;
        weights1[6950] <= 16'b1111111111011011;
        weights1[6951] <= 16'b1111111111100010;
        weights1[6952] <= 16'b1111111111111110;
        weights1[6953] <= 16'b0000000000000010;
        weights1[6954] <= 16'b1111111111101001;
        weights1[6955] <= 16'b0000000000010100;
        weights1[6956] <= 16'b0000000000010010;
        weights1[6957] <= 16'b0000000000001001;
        weights1[6958] <= 16'b1111111111110100;
        weights1[6959] <= 16'b0000000000000101;
        weights1[6960] <= 16'b0000000000010010;
        weights1[6961] <= 16'b1111111111100010;
        weights1[6962] <= 16'b0000000000011010;
        weights1[6963] <= 16'b1111111111111100;
        weights1[6964] <= 16'b1111111111101101;
        weights1[6965] <= 16'b1111111111111000;
        weights1[6966] <= 16'b1111111111100111;
        weights1[6967] <= 16'b1111111111001010;
        weights1[6968] <= 16'b1111111111110010;
        weights1[6969] <= 16'b0000000000000010;
        weights1[6970] <= 16'b1111111111111111;
        weights1[6971] <= 16'b0000000000000000;
        weights1[6972] <= 16'b0000000000000011;
        weights1[6973] <= 16'b0000000000000111;
        weights1[6974] <= 16'b0000000000000001;
        weights1[6975] <= 16'b0000000000000111;
        weights1[6976] <= 16'b0000000000001010;
        weights1[6977] <= 16'b0000000000000100;
        weights1[6978] <= 16'b1111111111110010;
        weights1[6979] <= 16'b1111111111101110;
        weights1[6980] <= 16'b1111111111110101;
        weights1[6981] <= 16'b1111111111101100;
        weights1[6982] <= 16'b1111111111111110;
        weights1[6983] <= 16'b1111111111010011;
        weights1[6984] <= 16'b1111111111010001;
        weights1[6985] <= 16'b1111111111011101;
        weights1[6986] <= 16'b1111111111101111;
        weights1[6987] <= 16'b1111111111111001;
        weights1[6988] <= 16'b1111111111001001;
        weights1[6989] <= 16'b1111111111100110;
        weights1[6990] <= 16'b1111111111010110;
        weights1[6991] <= 16'b1111111111001011;
        weights1[6992] <= 16'b1111111111001001;
        weights1[6993] <= 16'b1111111110111100;
        weights1[6994] <= 16'b1111111110111101;
        weights1[6995] <= 16'b1111111111000111;
        weights1[6996] <= 16'b1111111111100111;
        weights1[6997] <= 16'b1111111111111001;
        weights1[6998] <= 16'b1111111111111011;
        weights1[6999] <= 16'b1111111111111011;
        weights1[7000] <= 16'b0000000000000000;
        weights1[7001] <= 16'b0000000000000000;
        weights1[7002] <= 16'b1111111111111011;
        weights1[7003] <= 16'b1111111111111001;
        weights1[7004] <= 16'b1111111111110101;
        weights1[7005] <= 16'b1111111111110000;
        weights1[7006] <= 16'b1111111111011101;
        weights1[7007] <= 16'b1111111111100010;
        weights1[7008] <= 16'b1111111111100001;
        weights1[7009] <= 16'b1111111111011101;
        weights1[7010] <= 16'b1111111111001110;
        weights1[7011] <= 16'b1111111111010100;
        weights1[7012] <= 16'b1111111111001111;
        weights1[7013] <= 16'b1111111111000110;
        weights1[7014] <= 16'b1111111111001001;
        weights1[7015] <= 16'b1111111110101011;
        weights1[7016] <= 16'b1111111111001110;
        weights1[7017] <= 16'b1111111110111101;
        weights1[7018] <= 16'b1111111110111000;
        weights1[7019] <= 16'b1111111110101101;
        weights1[7020] <= 16'b1111111110110100;
        weights1[7021] <= 16'b1111111111000010;
        weights1[7022] <= 16'b1111111111010101;
        weights1[7023] <= 16'b1111111111011000;
        weights1[7024] <= 16'b1111111111100100;
        weights1[7025] <= 16'b1111111111110100;
        weights1[7026] <= 16'b1111111111111010;
        weights1[7027] <= 16'b1111111111111100;
        weights1[7028] <= 16'b1111111111111110;
        weights1[7029] <= 16'b0000000000000000;
        weights1[7030] <= 16'b1111111111111111;
        weights1[7031] <= 16'b1111111111111000;
        weights1[7032] <= 16'b1111111111110011;
        weights1[7033] <= 16'b1111111111101111;
        weights1[7034] <= 16'b1111111111100101;
        weights1[7035] <= 16'b1111111111001110;
        weights1[7036] <= 16'b1111111111001100;
        weights1[7037] <= 16'b1111111111001101;
        weights1[7038] <= 16'b1111111110111000;
        weights1[7039] <= 16'b1111111111000111;
        weights1[7040] <= 16'b1111111111000011;
        weights1[7041] <= 16'b1111111110110110;
        weights1[7042] <= 16'b1111111110101110;
        weights1[7043] <= 16'b1111111110110101;
        weights1[7044] <= 16'b1111111111000001;
        weights1[7045] <= 16'b1111111111000001;
        weights1[7046] <= 16'b1111111111001101;
        weights1[7047] <= 16'b1111111111010010;
        weights1[7048] <= 16'b1111111111010110;
        weights1[7049] <= 16'b1111111111010110;
        weights1[7050] <= 16'b1111111111101000;
        weights1[7051] <= 16'b1111111111101101;
        weights1[7052] <= 16'b1111111111101110;
        weights1[7053] <= 16'b1111111111111010;
        weights1[7054] <= 16'b1111111111111101;
        weights1[7055] <= 16'b1111111111111110;
        weights1[7056] <= 16'b0000000000000000;
        weights1[7057] <= 16'b0000000000000000;
        weights1[7058] <= 16'b1111111111111111;
        weights1[7059] <= 16'b1111111111111111;
        weights1[7060] <= 16'b1111111111111111;
        weights1[7061] <= 16'b1111111111111101;
        weights1[7062] <= 16'b1111111111111100;
        weights1[7063] <= 16'b1111111111111100;
        weights1[7064] <= 16'b1111111111110101;
        weights1[7065] <= 16'b1111111111110101;
        weights1[7066] <= 16'b1111111111110111;
        weights1[7067] <= 16'b1111111111110111;
        weights1[7068] <= 16'b1111111111110010;
        weights1[7069] <= 16'b1111111111110100;
        weights1[7070] <= 16'b1111111111101110;
        weights1[7071] <= 16'b1111111111101100;
        weights1[7072] <= 16'b1111111111101001;
        weights1[7073] <= 16'b1111111111101011;
        weights1[7074] <= 16'b1111111111101101;
        weights1[7075] <= 16'b1111111111101111;
        weights1[7076] <= 16'b1111111111101110;
        weights1[7077] <= 16'b1111111111101010;
        weights1[7078] <= 16'b1111111111110010;
        weights1[7079] <= 16'b1111111111110110;
        weights1[7080] <= 16'b1111111111110110;
        weights1[7081] <= 16'b1111111111111000;
        weights1[7082] <= 16'b1111111111111111;
        weights1[7083] <= 16'b0000000000000000;
        weights1[7084] <= 16'b1111111111111110;
        weights1[7085] <= 16'b1111111111111111;
        weights1[7086] <= 16'b1111111111111110;
        weights1[7087] <= 16'b1111111111111010;
        weights1[7088] <= 16'b1111111111111011;
        weights1[7089] <= 16'b1111111111111010;
        weights1[7090] <= 16'b1111111111111000;
        weights1[7091] <= 16'b0000000000000000;
        weights1[7092] <= 16'b1111111111110101;
        weights1[7093] <= 16'b1111111111111000;
        weights1[7094] <= 16'b1111111111110111;
        weights1[7095] <= 16'b1111111111110110;
        weights1[7096] <= 16'b0000000000000001;
        weights1[7097] <= 16'b1111111111101000;
        weights1[7098] <= 16'b1111111111011111;
        weights1[7099] <= 16'b1111111111110001;
        weights1[7100] <= 16'b1111111111110000;
        weights1[7101] <= 16'b1111111111110010;
        weights1[7102] <= 16'b1111111111110000;
        weights1[7103] <= 16'b1111111111110001;
        weights1[7104] <= 16'b1111111111110001;
        weights1[7105] <= 16'b1111111111110100;
        weights1[7106] <= 16'b1111111111100110;
        weights1[7107] <= 16'b1111111111101000;
        weights1[7108] <= 16'b1111111111101111;
        weights1[7109] <= 16'b1111111111111010;
        weights1[7110] <= 16'b1111111111110111;
        weights1[7111] <= 16'b1111111111111110;
        weights1[7112] <= 16'b1111111111111100;
        weights1[7113] <= 16'b1111111111111010;
        weights1[7114] <= 16'b1111111111111100;
        weights1[7115] <= 16'b1111111111110111;
        weights1[7116] <= 16'b1111111111110110;
        weights1[7117] <= 16'b1111111111111001;
        weights1[7118] <= 16'b0000000000000000;
        weights1[7119] <= 16'b0000000000000100;
        weights1[7120] <= 16'b0000000000000000;
        weights1[7121] <= 16'b0000000000000000;
        weights1[7122] <= 16'b1111111111111001;
        weights1[7123] <= 16'b1111111111110100;
        weights1[7124] <= 16'b1111111111110101;
        weights1[7125] <= 16'b1111111111100011;
        weights1[7126] <= 16'b1111111111111011;
        weights1[7127] <= 16'b1111111111101111;
        weights1[7128] <= 16'b1111111111111000;
        weights1[7129] <= 16'b1111111111100110;
        weights1[7130] <= 16'b1111111111110001;
        weights1[7131] <= 16'b1111111111110100;
        weights1[7132] <= 16'b1111111111100001;
        weights1[7133] <= 16'b1111111111110001;
        weights1[7134] <= 16'b1111111111110111;
        weights1[7135] <= 16'b1111111111101110;
        weights1[7136] <= 16'b1111111111110101;
        weights1[7137] <= 16'b1111111111111001;
        weights1[7138] <= 16'b1111111111110011;
        weights1[7139] <= 16'b1111111111110101;
        weights1[7140] <= 16'b1111111111111100;
        weights1[7141] <= 16'b1111111111111110;
        weights1[7142] <= 16'b1111111111111001;
        weights1[7143] <= 16'b1111111111110100;
        weights1[7144] <= 16'b1111111111110110;
        weights1[7145] <= 16'b1111111111110101;
        weights1[7146] <= 16'b1111111111110110;
        weights1[7147] <= 16'b1111111111111011;
        weights1[7148] <= 16'b1111111111110110;
        weights1[7149] <= 16'b1111111111111010;
        weights1[7150] <= 16'b1111111111110011;
        weights1[7151] <= 16'b1111111111111100;
        weights1[7152] <= 16'b1111111111111010;
        weights1[7153] <= 16'b0000000000000000;
        weights1[7154] <= 16'b1111111111110100;
        weights1[7155] <= 16'b1111111111111111;
        weights1[7156] <= 16'b0000000000001001;
        weights1[7157] <= 16'b1111111111111010;
        weights1[7158] <= 16'b1111111111101110;
        weights1[7159] <= 16'b0000000000000001;
        weights1[7160] <= 16'b1111111111110111;
        weights1[7161] <= 16'b1111111111110011;
        weights1[7162] <= 16'b1111111111111100;
        weights1[7163] <= 16'b1111111111110100;
        weights1[7164] <= 16'b1111111111110100;
        weights1[7165] <= 16'b1111111111111001;
        weights1[7166] <= 16'b1111111111110100;
        weights1[7167] <= 16'b1111111111111011;
        weights1[7168] <= 16'b1111111111111101;
        weights1[7169] <= 16'b1111111111111110;
        weights1[7170] <= 16'b1111111111110101;
        weights1[7171] <= 16'b1111111111110110;
        weights1[7172] <= 16'b1111111111110011;
        weights1[7173] <= 16'b1111111111110100;
        weights1[7174] <= 16'b1111111111100110;
        weights1[7175] <= 16'b1111111111100101;
        weights1[7176] <= 16'b1111111111110110;
        weights1[7177] <= 16'b1111111111110011;
        weights1[7178] <= 16'b1111111111101111;
        weights1[7179] <= 16'b1111111111111111;
        weights1[7180] <= 16'b1111111111111011;
        weights1[7181] <= 16'b1111111111101010;
        weights1[7182] <= 16'b1111111111111001;
        weights1[7183] <= 16'b1111111111110111;
        weights1[7184] <= 16'b1111111111011001;
        weights1[7185] <= 16'b0000000000000110;
        weights1[7186] <= 16'b1111111111101110;
        weights1[7187] <= 16'b1111111111101100;
        weights1[7188] <= 16'b0000000000000111;
        weights1[7189] <= 16'b1111111111110110;
        weights1[7190] <= 16'b0000000000001011;
        weights1[7191] <= 16'b1111111111110000;
        weights1[7192] <= 16'b0000000000010101;
        weights1[7193] <= 16'b0000000000000000;
        weights1[7194] <= 16'b1111111111110111;
        weights1[7195] <= 16'b1111111111111001;
        weights1[7196] <= 16'b1111111111111111;
        weights1[7197] <= 16'b1111111111111100;
        weights1[7198] <= 16'b0000000000000011;
        weights1[7199] <= 16'b1111111111111001;
        weights1[7200] <= 16'b1111111111110001;
        weights1[7201] <= 16'b1111111111110000;
        weights1[7202] <= 16'b0000000000000010;
        weights1[7203] <= 16'b1111111111101111;
        weights1[7204] <= 16'b1111111111110101;
        weights1[7205] <= 16'b1111111111111111;
        weights1[7206] <= 16'b1111111111111111;
        weights1[7207] <= 16'b1111111111101110;
        weights1[7208] <= 16'b1111111111110000;
        weights1[7209] <= 16'b0000000000000001;
        weights1[7210] <= 16'b1111111111111000;
        weights1[7211] <= 16'b1111111111100010;
        weights1[7212] <= 16'b0000000000000101;
        weights1[7213] <= 16'b1111111111110010;
        weights1[7214] <= 16'b1111111111111101;
        weights1[7215] <= 16'b0000000000000010;
        weights1[7216] <= 16'b1111111111101111;
        weights1[7217] <= 16'b1111111111100010;
        weights1[7218] <= 16'b0000000000001000;
        weights1[7219] <= 16'b0000000000011001;
        weights1[7220] <= 16'b0000000000000101;
        weights1[7221] <= 16'b1111111111101111;
        weights1[7222] <= 16'b1111111111111000;
        weights1[7223] <= 16'b1111111111110101;
        weights1[7224] <= 16'b1111111111111111;
        weights1[7225] <= 16'b0000000000000010;
        weights1[7226] <= 16'b1111111111111111;
        weights1[7227] <= 16'b1111111111110000;
        weights1[7228] <= 16'b1111111111110101;
        weights1[7229] <= 16'b0000000000000101;
        weights1[7230] <= 16'b1111111111011011;
        weights1[7231] <= 16'b1111111111110110;
        weights1[7232] <= 16'b1111111111011011;
        weights1[7233] <= 16'b1111111111011010;
        weights1[7234] <= 16'b1111111111111010;
        weights1[7235] <= 16'b1111111111100101;
        weights1[7236] <= 16'b1111111111110110;
        weights1[7237] <= 16'b1111111111110011;
        weights1[7238] <= 16'b1111111111111100;
        weights1[7239] <= 16'b1111111111101100;
        weights1[7240] <= 16'b1111111111111110;
        weights1[7241] <= 16'b1111111111111110;
        weights1[7242] <= 16'b1111111111111001;
        weights1[7243] <= 16'b1111111111111001;
        weights1[7244] <= 16'b0000000000000111;
        weights1[7245] <= 16'b0000000000000100;
        weights1[7246] <= 16'b1111111111010100;
        weights1[7247] <= 16'b1111111111101001;
        weights1[7248] <= 16'b0000000000001011;
        weights1[7249] <= 16'b1111111111110111;
        weights1[7250] <= 16'b1111111111110110;
        weights1[7251] <= 16'b1111111111110110;
        weights1[7252] <= 16'b0000000000000100;
        weights1[7253] <= 16'b0000000000000010;
        weights1[7254] <= 16'b0000000000000101;
        weights1[7255] <= 16'b1111111111110111;
        weights1[7256] <= 16'b1111111111110111;
        weights1[7257] <= 16'b1111111111100000;
        weights1[7258] <= 16'b1111111111100010;
        weights1[7259] <= 16'b1111111111100001;
        weights1[7260] <= 16'b1111111111111100;
        weights1[7261] <= 16'b1111111111101110;
        weights1[7262] <= 16'b1111111111100011;
        weights1[7263] <= 16'b1111111111100011;
        weights1[7264] <= 16'b1111111111011101;
        weights1[7265] <= 16'b1111111111110001;
        weights1[7266] <= 16'b1111111111101101;
        weights1[7267] <= 16'b0000000000000001;
        weights1[7268] <= 16'b1111111111101110;
        weights1[7269] <= 16'b0000000000001000;
        weights1[7270] <= 16'b1111111111101100;
        weights1[7271] <= 16'b1111111111101110;
        weights1[7272] <= 16'b1111111111011100;
        weights1[7273] <= 16'b1111111111100001;
        weights1[7274] <= 16'b1111111111111100;
        weights1[7275] <= 16'b1111111111011001;
        weights1[7276] <= 16'b1111111111101011;
        weights1[7277] <= 16'b1111111111101000;
        weights1[7278] <= 16'b1111111111110001;
        weights1[7279] <= 16'b1111111111100110;
        weights1[7280] <= 16'b0000000000000010;
        weights1[7281] <= 16'b0000000000000100;
        weights1[7282] <= 16'b0000000000001011;
        weights1[7283] <= 16'b1111111111111101;
        weights1[7284] <= 16'b1111111111110111;
        weights1[7285] <= 16'b1111111111010100;
        weights1[7286] <= 16'b1111111111011010;
        weights1[7287] <= 16'b1111111111110000;
        weights1[7288] <= 16'b1111111111011011;
        weights1[7289] <= 16'b1111111111001100;
        weights1[7290] <= 16'b1111111111100101;
        weights1[7291] <= 16'b1111111111011000;
        weights1[7292] <= 16'b1111111111111001;
        weights1[7293] <= 16'b1111111111011011;
        weights1[7294] <= 16'b1111111111100111;
        weights1[7295] <= 16'b1111111111100000;
        weights1[7296] <= 16'b1111111111110001;
        weights1[7297] <= 16'b1111111111100001;
        weights1[7298] <= 16'b1111111111110000;
        weights1[7299] <= 16'b1111111111100001;
        weights1[7300] <= 16'b0000000000000101;
        weights1[7301] <= 16'b1111111111110001;
        weights1[7302] <= 16'b1111111111111100;
        weights1[7303] <= 16'b1111111111101000;
        weights1[7304] <= 16'b1111111111001111;
        weights1[7305] <= 16'b1111111111011000;
        weights1[7306] <= 16'b1111111111110100;
        weights1[7307] <= 16'b1111111111100000;
        weights1[7308] <= 16'b0000000000000001;
        weights1[7309] <= 16'b0000000000000010;
        weights1[7310] <= 16'b0000000000001000;
        weights1[7311] <= 16'b0000000000000011;
        weights1[7312] <= 16'b1111111111110111;
        weights1[7313] <= 16'b1111111111100001;
        weights1[7314] <= 16'b1111111111100110;
        weights1[7315] <= 16'b1111111111101000;
        weights1[7316] <= 16'b1111111111010100;
        weights1[7317] <= 16'b1111111111110010;
        weights1[7318] <= 16'b1111111111100010;
        weights1[7319] <= 16'b1111111111100011;
        weights1[7320] <= 16'b1111111111100011;
        weights1[7321] <= 16'b1111111111101010;
        weights1[7322] <= 16'b1111111111101011;
        weights1[7323] <= 16'b1111111111011000;
        weights1[7324] <= 16'b1111111111101101;
        weights1[7325] <= 16'b1111111111011000;
        weights1[7326] <= 16'b1111111111101000;
        weights1[7327] <= 16'b1111111111100000;
        weights1[7328] <= 16'b1111111111010100;
        weights1[7329] <= 16'b1111111111011011;
        weights1[7330] <= 16'b1111111111100001;
        weights1[7331] <= 16'b1111111111011010;
        weights1[7332] <= 16'b1111111111100100;
        weights1[7333] <= 16'b1111111111100000;
        weights1[7334] <= 16'b1111111111011110;
        weights1[7335] <= 16'b1111111111011011;
        weights1[7336] <= 16'b0000000000000011;
        weights1[7337] <= 16'b1111111111111101;
        weights1[7338] <= 16'b1111111111111011;
        weights1[7339] <= 16'b1111111111101111;
        weights1[7340] <= 16'b1111111111011111;
        weights1[7341] <= 16'b1111111111101000;
        weights1[7342] <= 16'b1111111111111001;
        weights1[7343] <= 16'b1111111111110000;
        weights1[7344] <= 16'b1111111111010010;
        weights1[7345] <= 16'b1111111111100001;
        weights1[7346] <= 16'b1111111111101001;
        weights1[7347] <= 16'b1111111111011001;
        weights1[7348] <= 16'b1111111111100010;
        weights1[7349] <= 16'b1111111111100100;
        weights1[7350] <= 16'b1111111111011110;
        weights1[7351] <= 16'b1111111111011000;
        weights1[7352] <= 16'b1111111111010111;
        weights1[7353] <= 16'b1111111111100010;
        weights1[7354] <= 16'b1111111111011011;
        weights1[7355] <= 16'b1111111111011000;
        weights1[7356] <= 16'b1111111111100001;
        weights1[7357] <= 16'b1111111111011011;
        weights1[7358] <= 16'b1111111111011010;
        weights1[7359] <= 16'b1111111111011110;
        weights1[7360] <= 16'b1111111111001101;
        weights1[7361] <= 16'b1111111111100001;
        weights1[7362] <= 16'b1111111111011001;
        weights1[7363] <= 16'b1111111111011011;
        weights1[7364] <= 16'b1111111111111111;
        weights1[7365] <= 16'b1111111111111100;
        weights1[7366] <= 16'b0000000000000100;
        weights1[7367] <= 16'b1111111111110110;
        weights1[7368] <= 16'b1111111111110111;
        weights1[7369] <= 16'b1111111111110001;
        weights1[7370] <= 16'b1111111111111100;
        weights1[7371] <= 16'b1111111111111001;
        weights1[7372] <= 16'b1111111111110100;
        weights1[7373] <= 16'b1111111111111001;
        weights1[7374] <= 16'b1111111111110011;
        weights1[7375] <= 16'b1111111111010010;
        weights1[7376] <= 16'b1111111111100111;
        weights1[7377] <= 16'b1111111111011100;
        weights1[7378] <= 16'b1111111111010111;
        weights1[7379] <= 16'b1111111111101000;
        weights1[7380] <= 16'b1111111111100110;
        weights1[7381] <= 16'b1111111111011101;
        weights1[7382] <= 16'b1111111111100010;
        weights1[7383] <= 16'b1111111111111000;
        weights1[7384] <= 16'b1111111111011100;
        weights1[7385] <= 16'b1111111111100111;
        weights1[7386] <= 16'b1111111111010011;
        weights1[7387] <= 16'b1111111111010101;
        weights1[7388] <= 16'b1111111111000110;
        weights1[7389] <= 16'b1111111111011000;
        weights1[7390] <= 16'b1111111111011001;
        weights1[7391] <= 16'b1111111111100110;
        weights1[7392] <= 16'b0000000000000000;
        weights1[7393] <= 16'b0000000000000011;
        weights1[7394] <= 16'b1111111111111110;
        weights1[7395] <= 16'b0000000000001110;
        weights1[7396] <= 16'b0000000000000000;
        weights1[7397] <= 16'b0000000000000111;
        weights1[7398] <= 16'b1111111111110100;
        weights1[7399] <= 16'b1111111111110000;
        weights1[7400] <= 16'b0000000000000000;
        weights1[7401] <= 16'b1111111111011100;
        weights1[7402] <= 16'b1111111111101010;
        weights1[7403] <= 16'b1111111111010100;
        weights1[7404] <= 16'b1111111111110011;
        weights1[7405] <= 16'b1111111111011010;
        weights1[7406] <= 16'b1111111111110000;
        weights1[7407] <= 16'b1111111111110011;
        weights1[7408] <= 16'b1111111111010110;
        weights1[7409] <= 16'b1111111111100101;
        weights1[7410] <= 16'b1111111111100101;
        weights1[7411] <= 16'b1111111111100010;
        weights1[7412] <= 16'b1111111111001100;
        weights1[7413] <= 16'b1111111111101010;
        weights1[7414] <= 16'b1111111111011111;
        weights1[7415] <= 16'b1111111111010111;
        weights1[7416] <= 16'b1111111111000001;
        weights1[7417] <= 16'b1111111111011111;
        weights1[7418] <= 16'b1111111111101001;
        weights1[7419] <= 16'b1111111111100101;
        weights1[7420] <= 16'b1111111111111101;
        weights1[7421] <= 16'b0000000000001110;
        weights1[7422] <= 16'b0000000000000101;
        weights1[7423] <= 16'b0000000000110010;
        weights1[7424] <= 16'b0000000000010100;
        weights1[7425] <= 16'b0000000000000000;
        weights1[7426] <= 16'b0000000000100110;
        weights1[7427] <= 16'b1111111111101101;
        weights1[7428] <= 16'b1111111111111000;
        weights1[7429] <= 16'b1111111111111010;
        weights1[7430] <= 16'b0000000000001011;
        weights1[7431] <= 16'b1111111111101110;
        weights1[7432] <= 16'b1111111111011100;
        weights1[7433] <= 16'b1111111111101010;
        weights1[7434] <= 16'b1111111111110101;
        weights1[7435] <= 16'b1111111111010111;
        weights1[7436] <= 16'b1111111111100101;
        weights1[7437] <= 16'b1111111111111011;
        weights1[7438] <= 16'b1111111111100101;
        weights1[7439] <= 16'b1111111110111101;
        weights1[7440] <= 16'b1111111111100000;
        weights1[7441] <= 16'b1111111111100111;
        weights1[7442] <= 16'b1111111111101000;
        weights1[7443] <= 16'b1111111111101011;
        weights1[7444] <= 16'b1111111111101110;
        weights1[7445] <= 16'b1111111111100010;
        weights1[7446] <= 16'b1111111111110010;
        weights1[7447] <= 16'b1111111111101111;
        weights1[7448] <= 16'b1111111111111111;
        weights1[7449] <= 16'b0000000000010101;
        weights1[7450] <= 16'b0000000000110000;
        weights1[7451] <= 16'b0000000000110111;
        weights1[7452] <= 16'b0000000000111010;
        weights1[7453] <= 16'b0000000000010100;
        weights1[7454] <= 16'b0000000000011011;
        weights1[7455] <= 16'b0000000000011111;
        weights1[7456] <= 16'b1111111111110111;
        weights1[7457] <= 16'b0000000000000100;
        weights1[7458] <= 16'b1111111111001101;
        weights1[7459] <= 16'b1111111111100000;
        weights1[7460] <= 16'b1111111111101100;
        weights1[7461] <= 16'b1111111111100101;
        weights1[7462] <= 16'b1111111111100011;
        weights1[7463] <= 16'b1111111111100100;
        weights1[7464] <= 16'b1111111111110100;
        weights1[7465] <= 16'b1111111111111111;
        weights1[7466] <= 16'b1111111111110001;
        weights1[7467] <= 16'b1111111111101110;
        weights1[7468] <= 16'b0000000000001001;
        weights1[7469] <= 16'b0000000000001000;
        weights1[7470] <= 16'b1111111111111010;
        weights1[7471] <= 16'b0000000000001000;
        weights1[7472] <= 16'b0000000000001001;
        weights1[7473] <= 16'b0000000000011000;
        weights1[7474] <= 16'b0000000000000000;
        weights1[7475] <= 16'b1111111111111111;
        weights1[7476] <= 16'b0000000000010100;
        weights1[7477] <= 16'b0000000000011011;
        weights1[7478] <= 16'b0000000000111011;
        weights1[7479] <= 16'b0000000000110011;
        weights1[7480] <= 16'b0000000001000010;
        weights1[7481] <= 16'b0000000000101010;
        weights1[7482] <= 16'b0000000000110100;
        weights1[7483] <= 16'b0000000000100110;
        weights1[7484] <= 16'b0000000000100101;
        weights1[7485] <= 16'b0000000000100001;
        weights1[7486] <= 16'b0000000000001111;
        weights1[7487] <= 16'b1111111111101001;
        weights1[7488] <= 16'b1111111111111110;
        weights1[7489] <= 16'b0000000000000001;
        weights1[7490] <= 16'b1111111111110010;
        weights1[7491] <= 16'b1111111111101101;
        weights1[7492] <= 16'b1111111111101111;
        weights1[7493] <= 16'b0000000000000110;
        weights1[7494] <= 16'b1111111111111011;
        weights1[7495] <= 16'b0000000000011011;
        weights1[7496] <= 16'b0000000000010111;
        weights1[7497] <= 16'b0000000000001110;
        weights1[7498] <= 16'b0000000000001010;
        weights1[7499] <= 16'b1111111111101000;
        weights1[7500] <= 16'b0000000000010001;
        weights1[7501] <= 16'b0000000000100111;
        weights1[7502] <= 16'b0000000000100001;
        weights1[7503] <= 16'b0000000000011000;
        weights1[7504] <= 16'b0000000000011010;
        weights1[7505] <= 16'b0000000000011110;
        weights1[7506] <= 16'b0000000000101000;
        weights1[7507] <= 16'b0000000000110001;
        weights1[7508] <= 16'b0000000000111001;
        weights1[7509] <= 16'b0000000001001010;
        weights1[7510] <= 16'b0000000000110110;
        weights1[7511] <= 16'b0000000001000110;
        weights1[7512] <= 16'b0000000001000100;
        weights1[7513] <= 16'b0000000001000010;
        weights1[7514] <= 16'b0000000001001101;
        weights1[7515] <= 16'b0000000000100100;
        weights1[7516] <= 16'b0000000000101010;
        weights1[7517] <= 16'b0000000000100110;
        weights1[7518] <= 16'b0000000000011011;
        weights1[7519] <= 16'b0000000000010111;
        weights1[7520] <= 16'b0000000000001110;
        weights1[7521] <= 16'b0000000000011010;
        weights1[7522] <= 16'b0000000000010010;
        weights1[7523] <= 16'b0000000000010001;
        weights1[7524] <= 16'b0000000000101001;
        weights1[7525] <= 16'b0000000000110001;
        weights1[7526] <= 16'b0000000000100001;
        weights1[7527] <= 16'b0000000000010010;
        weights1[7528] <= 16'b0000000000101001;
        weights1[7529] <= 16'b0000000000111100;
        weights1[7530] <= 16'b0000000000101111;
        weights1[7531] <= 16'b0000000000011100;
        weights1[7532] <= 16'b0000000000011000;
        weights1[7533] <= 16'b0000000000100011;
        weights1[7534] <= 16'b0000000000101101;
        weights1[7535] <= 16'b0000000000011011;
        weights1[7536] <= 16'b0000000000011110;
        weights1[7537] <= 16'b0000000000101001;
        weights1[7538] <= 16'b0000000000100110;
        weights1[7539] <= 16'b0000000000110000;
        weights1[7540] <= 16'b0000000001010100;
        weights1[7541] <= 16'b0000000000111100;
        weights1[7542] <= 16'b0000000000110110;
        weights1[7543] <= 16'b0000000000111101;
        weights1[7544] <= 16'b0000000000101101;
        weights1[7545] <= 16'b0000000001000001;
        weights1[7546] <= 16'b0000000000101111;
        weights1[7547] <= 16'b0000000000100110;
        weights1[7548] <= 16'b0000000000110110;
        weights1[7549] <= 16'b0000000000100101;
        weights1[7550] <= 16'b0000000000101111;
        weights1[7551] <= 16'b0000000000101001;
        weights1[7552] <= 16'b0000000000111011;
        weights1[7553] <= 16'b0000000001000000;
        weights1[7554] <= 16'b0000000001010001;
        weights1[7555] <= 16'b0000000000101010;
        weights1[7556] <= 16'b0000000000110111;
        weights1[7557] <= 16'b0000000001010000;
        weights1[7558] <= 16'b0000000000101110;
        weights1[7559] <= 16'b0000000000101110;
        weights1[7560] <= 16'b0000000000001001;
        weights1[7561] <= 16'b0000000000010101;
        weights1[7562] <= 16'b0000000000011101;
        weights1[7563] <= 16'b0000000000011011;
        weights1[7564] <= 16'b0000000000100110;
        weights1[7565] <= 16'b0000000000100011;
        weights1[7566] <= 16'b0000000000101010;
        weights1[7567] <= 16'b0000000000110010;
        weights1[7568] <= 16'b0000000000101000;
        weights1[7569] <= 16'b0000000000100110;
        weights1[7570] <= 16'b0000000001000111;
        weights1[7571] <= 16'b0000000000101000;
        weights1[7572] <= 16'b0000000001001111;
        weights1[7573] <= 16'b0000000000110100;
        weights1[7574] <= 16'b0000000001010000;
        weights1[7575] <= 16'b0000000000101011;
        weights1[7576] <= 16'b0000000000111010;
        weights1[7577] <= 16'b0000000000110101;
        weights1[7578] <= 16'b0000000000101001;
        weights1[7579] <= 16'b0000000000110100;
        weights1[7580] <= 16'b0000000000111010;
        weights1[7581] <= 16'b0000000000111010;
        weights1[7582] <= 16'b0000000000111000;
        weights1[7583] <= 16'b0000000000100111;
        weights1[7584] <= 16'b0000000001010010;
        weights1[7585] <= 16'b0000000001000001;
        weights1[7586] <= 16'b0000000000110100;
        weights1[7587] <= 16'b0000000000101010;
        weights1[7588] <= 16'b0000000000001001;
        weights1[7589] <= 16'b0000000000001011;
        weights1[7590] <= 16'b0000000000001010;
        weights1[7591] <= 16'b0000000000001101;
        weights1[7592] <= 16'b0000000000010010;
        weights1[7593] <= 16'b0000000000001010;
        weights1[7594] <= 16'b0000000000011001;
        weights1[7595] <= 16'b0000000000100000;
        weights1[7596] <= 16'b0000000000110000;
        weights1[7597] <= 16'b0000000000110110;
        weights1[7598] <= 16'b0000000000101101;
        weights1[7599] <= 16'b0000000000101110;
        weights1[7600] <= 16'b0000000000110110;
        weights1[7601] <= 16'b0000000000111011;
        weights1[7602] <= 16'b0000000000110011;
        weights1[7603] <= 16'b0000000000110101;
        weights1[7604] <= 16'b0000000000101010;
        weights1[7605] <= 16'b0000000000110100;
        weights1[7606] <= 16'b0000000000111000;
        weights1[7607] <= 16'b0000000000111010;
        weights1[7608] <= 16'b0000000000101110;
        weights1[7609] <= 16'b0000000001000110;
        weights1[7610] <= 16'b0000000000111110;
        weights1[7611] <= 16'b0000000000111000;
        weights1[7612] <= 16'b0000000000101100;
        weights1[7613] <= 16'b0000000000100101;
        weights1[7614] <= 16'b0000000000101110;
        weights1[7615] <= 16'b0000000000100100;
        weights1[7616] <= 16'b0000000000001000;
        weights1[7617] <= 16'b0000000000000010;
        weights1[7618] <= 16'b1111111111111111;
        weights1[7619] <= 16'b0000000000000101;
        weights1[7620] <= 16'b0000000000010001;
        weights1[7621] <= 16'b0000000000001100;
        weights1[7622] <= 16'b1111111111110100;
        weights1[7623] <= 16'b0000000000011001;
        weights1[7624] <= 16'b0000000000000110;
        weights1[7625] <= 16'b0000000000000100;
        weights1[7626] <= 16'b0000000000010100;
        weights1[7627] <= 16'b0000000000101011;
        weights1[7628] <= 16'b0000000000011010;
        weights1[7629] <= 16'b0000000000001101;
        weights1[7630] <= 16'b0000000000011101;
        weights1[7631] <= 16'b0000000000110101;
        weights1[7632] <= 16'b0000000000100111;
        weights1[7633] <= 16'b0000000000101110;
        weights1[7634] <= 16'b0000000001000111;
        weights1[7635] <= 16'b0000000000110101;
        weights1[7636] <= 16'b0000000000110100;
        weights1[7637] <= 16'b1111111111111001;
        weights1[7638] <= 16'b0000000000101100;
        weights1[7639] <= 16'b0000000000011000;
        weights1[7640] <= 16'b0000000000010010;
        weights1[7641] <= 16'b0000000000010001;
        weights1[7642] <= 16'b0000000000100011;
        weights1[7643] <= 16'b0000000000100000;
        weights1[7644] <= 16'b0000000000000000;
        weights1[7645] <= 16'b1111111111111011;
        weights1[7646] <= 16'b1111111111110110;
        weights1[7647] <= 16'b1111111111110101;
        weights1[7648] <= 16'b0000000000001001;
        weights1[7649] <= 16'b0000000000010100;
        weights1[7650] <= 16'b0000000000010101;
        weights1[7651] <= 16'b0000000000000000;
        weights1[7652] <= 16'b1111111111110110;
        weights1[7653] <= 16'b0000000000001010;
        weights1[7654] <= 16'b0000000000000111;
        weights1[7655] <= 16'b1111111111111010;
        weights1[7656] <= 16'b0000000000001011;
        weights1[7657] <= 16'b0000000000011001;
        weights1[7658] <= 16'b0000000000011101;
        weights1[7659] <= 16'b1111111111111000;
        weights1[7660] <= 16'b0000000000100000;
        weights1[7661] <= 16'b0000000000010001;
        weights1[7662] <= 16'b0000000000001000;
        weights1[7663] <= 16'b0000000000000100;
        weights1[7664] <= 16'b0000000000011110;
        weights1[7665] <= 16'b0000000000011110;
        weights1[7666] <= 16'b0000000000100101;
        weights1[7667] <= 16'b0000000000010111;
        weights1[7668] <= 16'b0000000000010000;
        weights1[7669] <= 16'b0000000000001110;
        weights1[7670] <= 16'b0000000000010100;
        weights1[7671] <= 16'b0000000000001010;
        weights1[7672] <= 16'b0000000000000000;
        weights1[7673] <= 16'b1111111111110100;
        weights1[7674] <= 16'b1111111111100111;
        weights1[7675] <= 16'b1111111111111110;
        weights1[7676] <= 16'b1111111111111110;
        weights1[7677] <= 16'b0000000000001011;
        weights1[7678] <= 16'b1111111111110110;
        weights1[7679] <= 16'b0000000000001100;
        weights1[7680] <= 16'b1111111111101111;
        weights1[7681] <= 16'b0000000000001101;
        weights1[7682] <= 16'b1111111111111011;
        weights1[7683] <= 16'b0000000000010001;
        weights1[7684] <= 16'b1111111111111111;
        weights1[7685] <= 16'b0000000000000000;
        weights1[7686] <= 16'b1111111111110000;
        weights1[7687] <= 16'b1111111111111010;
        weights1[7688] <= 16'b1111111111110101;
        weights1[7689] <= 16'b0000000000000111;
        weights1[7690] <= 16'b0000000000001001;
        weights1[7691] <= 16'b0000000000001100;
        weights1[7692] <= 16'b0000000000010100;
        weights1[7693] <= 16'b0000000000010001;
        weights1[7694] <= 16'b0000000000001101;
        weights1[7695] <= 16'b0000000000000010;
        weights1[7696] <= 16'b0000000000010001;
        weights1[7697] <= 16'b0000000000001100;
        weights1[7698] <= 16'b1111111111111110;
        weights1[7699] <= 16'b0000000000000110;
        weights1[7700] <= 16'b1111111111111010;
        weights1[7701] <= 16'b1111111111101100;
        weights1[7702] <= 16'b1111111111100000;
        weights1[7703] <= 16'b1111111111110001;
        weights1[7704] <= 16'b1111111111101011;
        weights1[7705] <= 16'b1111111111101001;
        weights1[7706] <= 16'b1111111111100111;
        weights1[7707] <= 16'b1111111111110110;
        weights1[7708] <= 16'b1111111111101001;
        weights1[7709] <= 16'b1111111111110011;
        weights1[7710] <= 16'b1111111111110100;
        weights1[7711] <= 16'b1111111111100110;
        weights1[7712] <= 16'b1111111111100010;
        weights1[7713] <= 16'b1111111111011110;
        weights1[7714] <= 16'b1111111111101100;
        weights1[7715] <= 16'b0000000000011101;
        weights1[7716] <= 16'b1111111111011010;
        weights1[7717] <= 16'b1111111111101101;
        weights1[7718] <= 16'b0000000000001001;
        weights1[7719] <= 16'b0000000000000001;
        weights1[7720] <= 16'b1111111111111110;
        weights1[7721] <= 16'b1111111111110101;
        weights1[7722] <= 16'b1111111111111111;
        weights1[7723] <= 16'b1111111111110110;
        weights1[7724] <= 16'b1111111111111111;
        weights1[7725] <= 16'b1111111111111011;
        weights1[7726] <= 16'b1111111111111101;
        weights1[7727] <= 16'b1111111111111110;
        weights1[7728] <= 16'b1111111111111100;
        weights1[7729] <= 16'b1111111111111011;
        weights1[7730] <= 16'b1111111111101010;
        weights1[7731] <= 16'b1111111111011111;
        weights1[7732] <= 16'b1111111111001111;
        weights1[7733] <= 16'b1111111111001111;
        weights1[7734] <= 16'b1111111111010011;
        weights1[7735] <= 16'b1111111111011000;
        weights1[7736] <= 16'b1111111111010000;
        weights1[7737] <= 16'b1111111111111101;
        weights1[7738] <= 16'b1111111111101011;
        weights1[7739] <= 16'b1111111111111110;
        weights1[7740] <= 16'b1111111111111001;
        weights1[7741] <= 16'b0000000000001000;
        weights1[7742] <= 16'b1111111111100001;
        weights1[7743] <= 16'b0000000000000111;
        weights1[7744] <= 16'b1111111111111010;
        weights1[7745] <= 16'b0000000000001001;
        weights1[7746] <= 16'b1111111111110011;
        weights1[7747] <= 16'b1111111111011111;
        weights1[7748] <= 16'b1111111111110000;
        weights1[7749] <= 16'b1111111111110101;
        weights1[7750] <= 16'b1111111111110010;
        weights1[7751] <= 16'b1111111111101101;
        weights1[7752] <= 16'b1111111111111001;
        weights1[7753] <= 16'b0000000000000110;
        weights1[7754] <= 16'b0000000000000111;
        weights1[7755] <= 16'b0000000000000010;
        weights1[7756] <= 16'b1111111111111100;
        weights1[7757] <= 16'b0000000000000011;
        weights1[7758] <= 16'b1111111111111001;
        weights1[7759] <= 16'b1111111111100001;
        weights1[7760] <= 16'b1111111111010000;
        weights1[7761] <= 16'b1111111111010110;
        weights1[7762] <= 16'b1111111111001101;
        weights1[7763] <= 16'b1111111111001110;
        weights1[7764] <= 16'b1111111111000101;
        weights1[7765] <= 16'b1111111111001011;
        weights1[7766] <= 16'b1111111111001011;
        weights1[7767] <= 16'b1111111111010110;
        weights1[7768] <= 16'b1111111111011111;
        weights1[7769] <= 16'b1111111111011000;
        weights1[7770] <= 16'b1111111111011000;
        weights1[7771] <= 16'b1111111111011101;
        weights1[7772] <= 16'b1111111111011010;
        weights1[7773] <= 16'b1111111111010111;
        weights1[7774] <= 16'b1111111111100101;
        weights1[7775] <= 16'b1111111111100100;
        weights1[7776] <= 16'b1111111111011000;
        weights1[7777] <= 16'b1111111111101000;
        weights1[7778] <= 16'b1111111111011110;
        weights1[7779] <= 16'b1111111111100011;
        weights1[7780] <= 16'b1111111111111000;
        weights1[7781] <= 16'b1111111111111111;
        weights1[7782] <= 16'b1111111111111110;
        weights1[7783] <= 16'b0000000000000000;
        weights1[7784] <= 16'b1111111111111110;
        weights1[7785] <= 16'b0000000000000000;
        weights1[7786] <= 16'b1111111111111011;
        weights1[7787] <= 16'b1111111111101110;
        weights1[7788] <= 16'b1111111111101110;
        weights1[7789] <= 16'b1111111111101011;
        weights1[7790] <= 16'b1111111111110100;
        weights1[7791] <= 16'b1111111111101100;
        weights1[7792] <= 16'b1111111111100011;
        weights1[7793] <= 16'b1111111111011100;
        weights1[7794] <= 16'b1111111111001000;
        weights1[7795] <= 16'b1111111111011101;
        weights1[7796] <= 16'b1111111111100111;
        weights1[7797] <= 16'b1111111111011011;
        weights1[7798] <= 16'b1111111111010011;
        weights1[7799] <= 16'b1111111111001011;
        weights1[7800] <= 16'b1111111111010111;
        weights1[7801] <= 16'b1111111111100011;
        weights1[7802] <= 16'b1111111111100010;
        weights1[7803] <= 16'b1111111111110001;
        weights1[7804] <= 16'b1111111111100011;
        weights1[7805] <= 16'b1111111111011111;
        weights1[7806] <= 16'b1111111111011111;
        weights1[7807] <= 16'b1111111111101110;
        weights1[7808] <= 16'b1111111111111100;
        weights1[7809] <= 16'b0000000000000010;
        weights1[7810] <= 16'b1111111111111110;
        weights1[7811] <= 16'b0000000000000000;
        weights1[7812] <= 16'b0000000000000010;
        weights1[7813] <= 16'b0000000000000011;
        weights1[7814] <= 16'b0000000000000011;
        weights1[7815] <= 16'b1111111111111110;
        weights1[7816] <= 16'b1111111111111010;
        weights1[7817] <= 16'b1111111111111111;
        weights1[7818] <= 16'b1111111111111100;
        weights1[7819] <= 16'b1111111111110110;
        weights1[7820] <= 16'b1111111111100001;
        weights1[7821] <= 16'b1111111111011111;
        weights1[7822] <= 16'b1111111111011111;
        weights1[7823] <= 16'b1111111111101110;
        weights1[7824] <= 16'b1111111111011110;
        weights1[7825] <= 16'b1111111111100101;
        weights1[7826] <= 16'b1111111111100000;
        weights1[7827] <= 16'b1111111111110001;
        weights1[7828] <= 16'b1111111111011111;
        weights1[7829] <= 16'b1111111111101001;
        weights1[7830] <= 16'b1111111111100000;
        weights1[7831] <= 16'b1111111111011011;
        weights1[7832] <= 16'b1111111111011000;
        weights1[7833] <= 16'b1111111111100011;
        weights1[7834] <= 16'b1111111111100100;
        weights1[7835] <= 16'b1111111111110001;
        weights1[7836] <= 16'b1111111111110011;
        weights1[7837] <= 16'b1111111111111101;
        weights1[7838] <= 16'b0000000000000001;
        weights1[7839] <= 16'b0000000000000010;
        weights1[7840] <= 16'b0000000000000000;
        weights1[7841] <= 16'b0000000000000000;
        weights1[7842] <= 16'b0000000000000000;
        weights1[7843] <= 16'b0000000000000000;
        weights1[7844] <= 16'b1111111111111110;
        weights1[7845] <= 16'b1111111111111111;
        weights1[7846] <= 16'b1111111111111111;
        weights1[7847] <= 16'b0000000000000001;
        weights1[7848] <= 16'b0000000000001011;
        weights1[7849] <= 16'b0000000000001011;
        weights1[7850] <= 16'b0000000000010101;
        weights1[7851] <= 16'b0000000000010001;
        weights1[7852] <= 16'b0000000000011111;
        weights1[7853] <= 16'b0000000000100110;
        weights1[7854] <= 16'b0000000000101010;
        weights1[7855] <= 16'b0000000000011010;
        weights1[7856] <= 16'b0000000000100001;
        weights1[7857] <= 16'b0000000000010001;
        weights1[7858] <= 16'b0000000000000011;
        weights1[7859] <= 16'b0000000000011111;
        weights1[7860] <= 16'b0000000000010100;
        weights1[7861] <= 16'b0000000000000110;
        weights1[7862] <= 16'b0000000000001111;
        weights1[7863] <= 16'b0000000000011011;
        weights1[7864] <= 16'b0000000000001101;
        weights1[7865] <= 16'b0000000000000101;
        weights1[7866] <= 16'b0000000000000010;
        weights1[7867] <= 16'b0000000000000000;
        weights1[7868] <= 16'b0000000000000000;
        weights1[7869] <= 16'b0000000000000000;
        weights1[7870] <= 16'b1111111111111111;
        weights1[7871] <= 16'b1111111111111011;
        weights1[7872] <= 16'b1111111111111010;
        weights1[7873] <= 16'b1111111111111111;
        weights1[7874] <= 16'b0000000000001001;
        weights1[7875] <= 16'b0000000000000100;
        weights1[7876] <= 16'b1111111111111010;
        weights1[7877] <= 16'b0000000000000011;
        weights1[7878] <= 16'b0000000000001000;
        weights1[7879] <= 16'b0000000000100001;
        weights1[7880] <= 16'b0000000000100010;
        weights1[7881] <= 16'b0000000000011010;
        weights1[7882] <= 16'b0000000000101100;
        weights1[7883] <= 16'b0000000000011010;
        weights1[7884] <= 16'b0000000000010010;
        weights1[7885] <= 16'b0000000000010100;
        weights1[7886] <= 16'b0000000000011101;
        weights1[7887] <= 16'b0000000000001000;
        weights1[7888] <= 16'b0000000000011110;
        weights1[7889] <= 16'b0000000000010000;
        weights1[7890] <= 16'b0000000000011100;
        weights1[7891] <= 16'b0000000000000111;
        weights1[7892] <= 16'b0000000000000010;
        weights1[7893] <= 16'b0000000000001110;
        weights1[7894] <= 16'b0000000000001010;
        weights1[7895] <= 16'b0000000000000011;
        weights1[7896] <= 16'b0000000000000000;
        weights1[7897] <= 16'b0000000000000001;
        weights1[7898] <= 16'b1111111111111110;
        weights1[7899] <= 16'b1111111111111100;
        weights1[7900] <= 16'b1111111111111001;
        weights1[7901] <= 16'b1111111111111101;
        weights1[7902] <= 16'b0000000000001010;
        weights1[7903] <= 16'b0000000000000100;
        weights1[7904] <= 16'b1111111111111101;
        weights1[7905] <= 16'b0000000000000001;
        weights1[7906] <= 16'b0000000000010011;
        weights1[7907] <= 16'b0000000000010100;
        weights1[7908] <= 16'b0000000000011100;
        weights1[7909] <= 16'b0000000000100101;
        weights1[7910] <= 16'b0000000000100010;
        weights1[7911] <= 16'b0000000000011010;
        weights1[7912] <= 16'b0000000000011100;
        weights1[7913] <= 16'b0000000000001100;
        weights1[7914] <= 16'b1111111111111111;
        weights1[7915] <= 16'b0000000000001100;
        weights1[7916] <= 16'b0000000000010000;
        weights1[7917] <= 16'b0000000000001101;
        weights1[7918] <= 16'b0000000000000111;
        weights1[7919] <= 16'b0000000000000101;
        weights1[7920] <= 16'b1111111111111110;
        weights1[7921] <= 16'b0000000000010000;
        weights1[7922] <= 16'b0000000000001000;
        weights1[7923] <= 16'b0000000000010101;
        weights1[7924] <= 16'b0000000000000001;
        weights1[7925] <= 16'b1111111111111111;
        weights1[7926] <= 16'b1111111111111100;
        weights1[7927] <= 16'b1111111111110101;
        weights1[7928] <= 16'b1111111111110110;
        weights1[7929] <= 16'b1111111111111100;
        weights1[7930] <= 16'b0000000000000101;
        weights1[7931] <= 16'b0000000000000010;
        weights1[7932] <= 16'b1111111111111010;
        weights1[7933] <= 16'b0000000000000011;
        weights1[7934] <= 16'b0000000000000010;
        weights1[7935] <= 16'b1111111111111001;
        weights1[7936] <= 16'b0000000000011011;
        weights1[7937] <= 16'b0000000000010110;
        weights1[7938] <= 16'b0000000000010110;
        weights1[7939] <= 16'b0000000000010101;
        weights1[7940] <= 16'b0000000000010011;
        weights1[7941] <= 16'b0000000000010011;
        weights1[7942] <= 16'b0000000000011010;
        weights1[7943] <= 16'b0000000000010001;
        weights1[7944] <= 16'b0000000000010111;
        weights1[7945] <= 16'b1111111111111001;
        weights1[7946] <= 16'b0000000000000010;
        weights1[7947] <= 16'b0000000000001000;
        weights1[7948] <= 16'b0000000000001110;
        weights1[7949] <= 16'b0000000000011000;
        weights1[7950] <= 16'b0000000000011011;
        weights1[7951] <= 16'b0000000000011100;
        weights1[7952] <= 16'b0000000000000000;
        weights1[7953] <= 16'b1111111111111101;
        weights1[7954] <= 16'b1111111111110111;
        weights1[7955] <= 16'b1111111111110000;
        weights1[7956] <= 16'b1111111111101100;
        weights1[7957] <= 16'b1111111111110000;
        weights1[7958] <= 16'b1111111111110000;
        weights1[7959] <= 16'b1111111111101100;
        weights1[7960] <= 16'b1111111111110000;
        weights1[7961] <= 16'b1111111111110110;
        weights1[7962] <= 16'b1111111111110001;
        weights1[7963] <= 16'b1111111111110000;
        weights1[7964] <= 16'b0000000000000001;
        weights1[7965] <= 16'b0000000000000011;
        weights1[7966] <= 16'b0000000000010100;
        weights1[7967] <= 16'b0000000000010110;
        weights1[7968] <= 16'b0000000000001011;
        weights1[7969] <= 16'b0000000000011001;
        weights1[7970] <= 16'b0000000000011000;
        weights1[7971] <= 16'b0000000000010000;
        weights1[7972] <= 16'b0000000000001111;
        weights1[7973] <= 16'b0000000000010101;
        weights1[7974] <= 16'b0000000000000111;
        weights1[7975] <= 16'b0000000000010010;
        weights1[7976] <= 16'b0000000000010011;
        weights1[7977] <= 16'b0000000000100010;
        weights1[7978] <= 16'b0000000000100100;
        weights1[7979] <= 16'b0000000000011000;
        weights1[7980] <= 16'b0000000000000000;
        weights1[7981] <= 16'b1111111111111101;
        weights1[7982] <= 16'b1111111111110001;
        weights1[7983] <= 16'b1111111111101011;
        weights1[7984] <= 16'b1111111111101110;
        weights1[7985] <= 16'b1111111111110000;
        weights1[7986] <= 16'b1111111111100000;
        weights1[7987] <= 16'b1111111111011001;
        weights1[7988] <= 16'b1111111111100010;
        weights1[7989] <= 16'b1111111111110011;
        weights1[7990] <= 16'b1111111111110100;
        weights1[7991] <= 16'b0000000000001011;
        weights1[7992] <= 16'b0000000000000000;
        weights1[7993] <= 16'b1111111111101000;
        weights1[7994] <= 16'b0000000000011101;
        weights1[7995] <= 16'b0000000000100111;
        weights1[7996] <= 16'b0000000000000001;
        weights1[7997] <= 16'b0000000000011001;
        weights1[7998] <= 16'b0000000000001111;
        weights1[7999] <= 16'b0000000000010010;
        weights1[8000] <= 16'b0000000000010011;
        weights1[8001] <= 16'b0000000000001010;
        weights1[8002] <= 16'b0000000000010011;
        weights1[8003] <= 16'b0000000000010110;
        weights1[8004] <= 16'b0000000000000110;
        weights1[8005] <= 16'b0000000000011011;
        weights1[8006] <= 16'b0000000000011100;
        weights1[8007] <= 16'b0000000000100000;
        weights1[8008] <= 16'b0000000000000000;
        weights1[8009] <= 16'b1111111111111011;
        weights1[8010] <= 16'b1111111111101010;
        weights1[8011] <= 16'b1111111111101000;
        weights1[8012] <= 16'b1111111111100100;
        weights1[8013] <= 16'b1111111111011101;
        weights1[8014] <= 16'b1111111111011010;
        weights1[8015] <= 16'b1111111111110100;
        weights1[8016] <= 16'b1111111111101101;
        weights1[8017] <= 16'b1111111111111000;
        weights1[8018] <= 16'b1111111111110011;
        weights1[8019] <= 16'b1111111111111011;
        weights1[8020] <= 16'b0000000000000110;
        weights1[8021] <= 16'b0000000000001001;
        weights1[8022] <= 16'b0000000000010010;
        weights1[8023] <= 16'b0000000000010101;
        weights1[8024] <= 16'b0000000000000100;
        weights1[8025] <= 16'b0000000000010000;
        weights1[8026] <= 16'b1111111111111010;
        weights1[8027] <= 16'b1111111111110100;
        weights1[8028] <= 16'b0000000000010001;
        weights1[8029] <= 16'b0000000000000101;
        weights1[8030] <= 16'b0000000000001000;
        weights1[8031] <= 16'b0000000000001011;
        weights1[8032] <= 16'b0000000000001010;
        weights1[8033] <= 16'b0000000000001100;
        weights1[8034] <= 16'b0000000000001101;
        weights1[8035] <= 16'b0000000000010101;
        weights1[8036] <= 16'b1111111111111100;
        weights1[8037] <= 16'b1111111111110010;
        weights1[8038] <= 16'b1111111111101000;
        weights1[8039] <= 16'b1111111111100010;
        weights1[8040] <= 16'b1111111111011101;
        weights1[8041] <= 16'b1111111111011000;
        weights1[8042] <= 16'b1111111111101010;
        weights1[8043] <= 16'b1111111111101010;
        weights1[8044] <= 16'b1111111111011101;
        weights1[8045] <= 16'b1111111111101000;
        weights1[8046] <= 16'b1111111111110011;
        weights1[8047] <= 16'b1111111111101110;
        weights1[8048] <= 16'b0000000000000110;
        weights1[8049] <= 16'b0000000000000111;
        weights1[8050] <= 16'b0000000000001001;
        weights1[8051] <= 16'b0000000000011001;
        weights1[8052] <= 16'b0000000000000101;
        weights1[8053] <= 16'b0000000000010000;
        weights1[8054] <= 16'b0000000000001111;
        weights1[8055] <= 16'b0000000000011110;
        weights1[8056] <= 16'b0000000000000111;
        weights1[8057] <= 16'b0000000000000110;
        weights1[8058] <= 16'b1111111111111011;
        weights1[8059] <= 16'b0000000000000110;
        weights1[8060] <= 16'b0000000000000111;
        weights1[8061] <= 16'b0000000000001000;
        weights1[8062] <= 16'b0000000000000100;
        weights1[8063] <= 16'b0000000000010111;
        weights1[8064] <= 16'b1111111111111110;
        weights1[8065] <= 16'b1111111111101101;
        weights1[8066] <= 16'b1111111111100110;
        weights1[8067] <= 16'b1111111111010010;
        weights1[8068] <= 16'b1111111111010010;
        weights1[8069] <= 16'b1111111111001011;
        weights1[8070] <= 16'b1111111111010101;
        weights1[8071] <= 16'b1111111111101111;
        weights1[8072] <= 16'b1111111111011011;
        weights1[8073] <= 16'b1111111111110001;
        weights1[8074] <= 16'b0000000000010001;
        weights1[8075] <= 16'b0000000000010000;
        weights1[8076] <= 16'b0000000000001001;
        weights1[8077] <= 16'b0000000000100000;
        weights1[8078] <= 16'b0000000000101001;
        weights1[8079] <= 16'b0000000000101100;
        weights1[8080] <= 16'b0000000000100101;
        weights1[8081] <= 16'b0000000000101100;
        weights1[8082] <= 16'b0000000000011010;
        weights1[8083] <= 16'b0000000000001100;
        weights1[8084] <= 16'b0000000000000110;
        weights1[8085] <= 16'b0000000000000111;
        weights1[8086] <= 16'b1111111111111101;
        weights1[8087] <= 16'b0000000000000101;
        weights1[8088] <= 16'b0000000000001001;
        weights1[8089] <= 16'b0000000000001110;
        weights1[8090] <= 16'b0000000000001010;
        weights1[8091] <= 16'b0000000000010000;
        weights1[8092] <= 16'b1111111111111001;
        weights1[8093] <= 16'b1111111111101110;
        weights1[8094] <= 16'b1111111111100010;
        weights1[8095] <= 16'b1111111111100000;
        weights1[8096] <= 16'b1111111111001101;
        weights1[8097] <= 16'b1111111111000001;
        weights1[8098] <= 16'b1111111110111101;
        weights1[8099] <= 16'b1111111110111101;
        weights1[8100] <= 16'b1111111111010111;
        weights1[8101] <= 16'b1111111111100111;
        weights1[8102] <= 16'b1111111111110111;
        weights1[8103] <= 16'b1111111111110111;
        weights1[8104] <= 16'b0000000000010001;
        weights1[8105] <= 16'b0000000000000111;
        weights1[8106] <= 16'b0000000000111100;
        weights1[8107] <= 16'b0000000001000110;
        weights1[8108] <= 16'b0000000001010000;
        weights1[8109] <= 16'b0000000000110001;
        weights1[8110] <= 16'b0000000000101101;
        weights1[8111] <= 16'b0000000000100001;
        weights1[8112] <= 16'b0000000000010110;
        weights1[8113] <= 16'b0000000000001101;
        weights1[8114] <= 16'b0000000000001111;
        weights1[8115] <= 16'b0000000000001101;
        weights1[8116] <= 16'b1111111111111101;
        weights1[8117] <= 16'b1111111111111111;
        weights1[8118] <= 16'b0000000000001101;
        weights1[8119] <= 16'b0000000000010001;
        weights1[8120] <= 16'b1111111111111010;
        weights1[8121] <= 16'b1111111111101000;
        weights1[8122] <= 16'b1111111111011110;
        weights1[8123] <= 16'b1111111111100100;
        weights1[8124] <= 16'b1111111111010001;
        weights1[8125] <= 16'b1111111111000001;
        weights1[8126] <= 16'b1111111110101011;
        weights1[8127] <= 16'b1111111110111000;
        weights1[8128] <= 16'b1111111110101110;
        weights1[8129] <= 16'b1111111110110101;
        weights1[8130] <= 16'b1111111111001011;
        weights1[8131] <= 16'b1111111111010111;
        weights1[8132] <= 16'b1111111111110101;
        weights1[8133] <= 16'b0000000000001111;
        weights1[8134] <= 16'b0000000000001110;
        weights1[8135] <= 16'b0000000000010110;
        weights1[8136] <= 16'b0000000001000000;
        weights1[8137] <= 16'b0000000000101110;
        weights1[8138] <= 16'b0000000000010111;
        weights1[8139] <= 16'b0000000000100101;
        weights1[8140] <= 16'b0000000000011100;
        weights1[8141] <= 16'b0000000000011001;
        weights1[8142] <= 16'b1111111111111100;
        weights1[8143] <= 16'b0000000000010111;
        weights1[8144] <= 16'b0000000000000011;
        weights1[8145] <= 16'b0000000000010001;
        weights1[8146] <= 16'b0000000000010101;
        weights1[8147] <= 16'b0000000000011010;
        weights1[8148] <= 16'b1111111111111101;
        weights1[8149] <= 16'b1111111111101111;
        weights1[8150] <= 16'b1111111111101101;
        weights1[8151] <= 16'b1111111111110011;
        weights1[8152] <= 16'b1111111111001011;
        weights1[8153] <= 16'b1111111111010011;
        weights1[8154] <= 16'b1111111111000110;
        weights1[8155] <= 16'b1111111110101101;
        weights1[8156] <= 16'b1111111110001110;
        weights1[8157] <= 16'b1111111110001000;
        weights1[8158] <= 16'b1111111110100110;
        weights1[8159] <= 16'b1111111111000111;
        weights1[8160] <= 16'b1111111111100000;
        weights1[8161] <= 16'b1111111111100101;
        weights1[8162] <= 16'b0000000000000111;
        weights1[8163] <= 16'b0000000000101011;
        weights1[8164] <= 16'b0000000000101111;
        weights1[8165] <= 16'b0000000000100010;
        weights1[8166] <= 16'b0000000000010000;
        weights1[8167] <= 16'b0000000000001010;
        weights1[8168] <= 16'b0000000000001110;
        weights1[8169] <= 16'b0000000000001110;
        weights1[8170] <= 16'b0000000000010110;
        weights1[8171] <= 16'b0000000000011100;
        weights1[8172] <= 16'b0000000000001010;
        weights1[8173] <= 16'b1111111111111001;
        weights1[8174] <= 16'b0000000000010000;
        weights1[8175] <= 16'b0000000000010111;
        weights1[8176] <= 16'b1111111111111010;
        weights1[8177] <= 16'b1111111111110101;
        weights1[8178] <= 16'b1111111111111010;
        weights1[8179] <= 16'b0000000000000001;
        weights1[8180] <= 16'b1111111111110011;
        weights1[8181] <= 16'b1111111111100100;
        weights1[8182] <= 16'b1111111111011111;
        weights1[8183] <= 16'b1111111110111111;
        weights1[8184] <= 16'b1111111110011011;
        weights1[8185] <= 16'b1111111110000001;
        weights1[8186] <= 16'b1111111110000110;
        weights1[8187] <= 16'b1111111101111110;
        weights1[8188] <= 16'b1111111110100001;
        weights1[8189] <= 16'b1111111111000111;
        weights1[8190] <= 16'b1111111111100111;
        weights1[8191] <= 16'b0000000000011001;
        weights1[8192] <= 16'b0000000000111101;
        weights1[8193] <= 16'b0000000000010000;
        weights1[8194] <= 16'b0000000000010001;
        weights1[8195] <= 16'b0000000000010011;
        weights1[8196] <= 16'b0000000000001101;
        weights1[8197] <= 16'b0000000000000011;
        weights1[8198] <= 16'b0000000000001010;
        weights1[8199] <= 16'b1111111111111111;
        weights1[8200] <= 16'b1111111111111000;
        weights1[8201] <= 16'b1111111111111011;
        weights1[8202] <= 16'b0000000000000101;
        weights1[8203] <= 16'b0000000000000000;
        weights1[8204] <= 16'b0000000000000100;
        weights1[8205] <= 16'b1111111111111111;
        weights1[8206] <= 16'b1111111111111011;
        weights1[8207] <= 16'b0000000000001001;
        weights1[8208] <= 16'b0000000000001000;
        weights1[8209] <= 16'b0000000000001011;
        weights1[8210] <= 16'b0000000000000000;
        weights1[8211] <= 16'b0000000000000000;
        weights1[8212] <= 16'b1111111111011111;
        weights1[8213] <= 16'b1111111110110001;
        weights1[8214] <= 16'b1111111110011000;
        weights1[8215] <= 16'b1111111110010000;
        weights1[8216] <= 16'b1111111101110011;
        weights1[8217] <= 16'b1111111110010000;
        weights1[8218] <= 16'b1111111110110001;
        weights1[8219] <= 16'b0000000000011100;
        weights1[8220] <= 16'b0000000000111101;
        weights1[8221] <= 16'b0000000000110100;
        weights1[8222] <= 16'b0000000000001001;
        weights1[8223] <= 16'b0000000000000111;
        weights1[8224] <= 16'b0000000000100000;
        weights1[8225] <= 16'b1111111111111000;
        weights1[8226] <= 16'b1111111111111110;
        weights1[8227] <= 16'b1111111111110111;
        weights1[8228] <= 16'b1111111111111101;
        weights1[8229] <= 16'b1111111111110111;
        weights1[8230] <= 16'b1111111111110010;
        weights1[8231] <= 16'b1111111111110000;
        weights1[8232] <= 16'b0000000000001001;
        weights1[8233] <= 16'b0000000000000011;
        weights1[8234] <= 16'b0000000000001010;
        weights1[8235] <= 16'b0000000000010010;
        weights1[8236] <= 16'b0000000000011011;
        weights1[8237] <= 16'b0000000000010110;
        weights1[8238] <= 16'b0000000000011000;
        weights1[8239] <= 16'b0000000000101010;
        weights1[8240] <= 16'b0000000000001101;
        weights1[8241] <= 16'b0000000000001000;
        weights1[8242] <= 16'b1111111111100100;
        weights1[8243] <= 16'b1111111110111011;
        weights1[8244] <= 16'b1111111110001110;
        weights1[8245] <= 16'b1111111110000110;
        weights1[8246] <= 16'b1111111110001111;
        weights1[8247] <= 16'b1111111111010001;
        weights1[8248] <= 16'b0000000000100011;
        weights1[8249] <= 16'b0000000000010000;
        weights1[8250] <= 16'b0000000000011100;
        weights1[8251] <= 16'b0000000000001110;
        weights1[8252] <= 16'b0000000000000110;
        weights1[8253] <= 16'b0000000000000101;
        weights1[8254] <= 16'b0000000000001000;
        weights1[8255] <= 16'b0000000000000111;
        weights1[8256] <= 16'b0000000000000011;
        weights1[8257] <= 16'b1111111111111001;
        weights1[8258] <= 16'b1111111111101101;
        weights1[8259] <= 16'b1111111111100001;
        weights1[8260] <= 16'b0000000000000101;
        weights1[8261] <= 16'b0000000000000111;
        weights1[8262] <= 16'b0000000000001110;
        weights1[8263] <= 16'b0000000000001001;
        weights1[8264] <= 16'b0000000000101000;
        weights1[8265] <= 16'b0000000000100011;
        weights1[8266] <= 16'b0000000000101101;
        weights1[8267] <= 16'b0000000000111101;
        weights1[8268] <= 16'b0000000000110110;
        weights1[8269] <= 16'b0000000000111000;
        weights1[8270] <= 16'b0000000000010001;
        weights1[8271] <= 16'b1111111111111001;
        weights1[8272] <= 16'b1111111111011011;
        weights1[8273] <= 16'b1111111110010100;
        weights1[8274] <= 16'b1111111110000100;
        weights1[8275] <= 16'b1111111110111111;
        weights1[8276] <= 16'b0000000000000000;
        weights1[8277] <= 16'b0000000000010110;
        weights1[8278] <= 16'b0000000000011100;
        weights1[8279] <= 16'b0000000000000001;
        weights1[8280] <= 16'b0000000000000010;
        weights1[8281] <= 16'b0000000000100001;
        weights1[8282] <= 16'b0000000000010101;
        weights1[8283] <= 16'b1111111111110101;
        weights1[8284] <= 16'b1111111111110101;
        weights1[8285] <= 16'b0000000000000010;
        weights1[8286] <= 16'b1111111111100111;
        weights1[8287] <= 16'b1111111111101010;
        weights1[8288] <= 16'b1111111111111111;
        weights1[8289] <= 16'b1111111111111111;
        weights1[8290] <= 16'b0000000000001011;
        weights1[8291] <= 16'b0000000000000011;
        weights1[8292] <= 16'b0000000000100111;
        weights1[8293] <= 16'b1111111111110000;
        weights1[8294] <= 16'b0000000000001100;
        weights1[8295] <= 16'b1111111111110100;
        weights1[8296] <= 16'b0000000000001011;
        weights1[8297] <= 16'b0000000000011111;
        weights1[8298] <= 16'b0000000000001100;
        weights1[8299] <= 16'b0000000000001011;
        weights1[8300] <= 16'b1111111111111011;
        weights1[8301] <= 16'b1111111111000100;
        weights1[8302] <= 16'b1111111110011000;
        weights1[8303] <= 16'b1111111110110001;
        weights1[8304] <= 16'b1111111111011111;
        weights1[8305] <= 16'b0000000000011010;
        weights1[8306] <= 16'b0000000000001110;
        weights1[8307] <= 16'b1111111111111101;
        weights1[8308] <= 16'b0000000000010010;
        weights1[8309] <= 16'b1111111111111101;
        weights1[8310] <= 16'b0000000000011000;
        weights1[8311] <= 16'b0000000000001101;
        weights1[8312] <= 16'b1111111111111000;
        weights1[8313] <= 16'b1111111111111111;
        weights1[8314] <= 16'b1111111111101111;
        weights1[8315] <= 16'b1111111111100100;
        weights1[8316] <= 16'b1111111111111001;
        weights1[8317] <= 16'b1111111111101101;
        weights1[8318] <= 16'b1111111111101100;
        weights1[8319] <= 16'b1111111111100111;
        weights1[8320] <= 16'b0000000000001011;
        weights1[8321] <= 16'b0000000000000100;
        weights1[8322] <= 16'b1111111111100110;
        weights1[8323] <= 16'b1111111111111110;
        weights1[8324] <= 16'b0000000000000001;
        weights1[8325] <= 16'b0000000000000000;
        weights1[8326] <= 16'b1111111111111000;
        weights1[8327] <= 16'b0000000000010000;
        weights1[8328] <= 16'b1111111111111111;
        weights1[8329] <= 16'b1111111111100000;
        weights1[8330] <= 16'b1111111110110100;
        weights1[8331] <= 16'b1111111110111101;
        weights1[8332] <= 16'b1111111111011110;
        weights1[8333] <= 16'b0000000000000011;
        weights1[8334] <= 16'b0000000000001010;
        weights1[8335] <= 16'b0000000000010000;
        weights1[8336] <= 16'b0000000000001100;
        weights1[8337] <= 16'b0000000000000101;
        weights1[8338] <= 16'b0000000000000000;
        weights1[8339] <= 16'b0000000000000100;
        weights1[8340] <= 16'b0000000000010000;
        weights1[8341] <= 16'b1111111111110111;
        weights1[8342] <= 16'b1111111111100111;
        weights1[8343] <= 16'b1111111111101000;
        weights1[8344] <= 16'b1111111111111000;
        weights1[8345] <= 16'b1111111111110001;
        weights1[8346] <= 16'b1111111111100100;
        weights1[8347] <= 16'b1111111111011111;
        weights1[8348] <= 16'b1111111111110011;
        weights1[8349] <= 16'b1111111111010110;
        weights1[8350] <= 16'b1111111111100110;
        weights1[8351] <= 16'b1111111111111010;
        weights1[8352] <= 16'b1111111111101111;
        weights1[8353] <= 16'b1111111111111101;
        weights1[8354] <= 16'b1111111111101000;
        weights1[8355] <= 16'b1111111111111011;
        weights1[8356] <= 16'b0000000000001001;
        weights1[8357] <= 16'b1111111111110010;
        weights1[8358] <= 16'b1111111111100000;
        weights1[8359] <= 16'b1111111111001110;
        weights1[8360] <= 16'b1111111111010110;
        weights1[8361] <= 16'b0000000000000100;
        weights1[8362] <= 16'b0000000000000101;
        weights1[8363] <= 16'b0000000000001111;
        weights1[8364] <= 16'b0000000000010011;
        weights1[8365] <= 16'b0000000000010011;
        weights1[8366] <= 16'b0000000000001111;
        weights1[8367] <= 16'b0000000000011100;
        weights1[8368] <= 16'b0000000000010001;
        weights1[8369] <= 16'b1111111111110011;
        weights1[8370] <= 16'b1111111111101100;
        weights1[8371] <= 16'b1111111111011101;
        weights1[8372] <= 16'b1111111111111010;
        weights1[8373] <= 16'b1111111111110111;
        weights1[8374] <= 16'b1111111111101101;
        weights1[8375] <= 16'b1111111111101000;
        weights1[8376] <= 16'b1111111111100110;
        weights1[8377] <= 16'b1111111111011100;
        weights1[8378] <= 16'b1111111111110101;
        weights1[8379] <= 16'b1111111111111110;
        weights1[8380] <= 16'b1111111111110001;
        weights1[8381] <= 16'b0000000000000001;
        weights1[8382] <= 16'b1111111111110001;
        weights1[8383] <= 16'b1111111111110100;
        weights1[8384] <= 16'b1111111111110110;
        weights1[8385] <= 16'b1111111111110100;
        weights1[8386] <= 16'b1111111111110100;
        weights1[8387] <= 16'b1111111111101111;
        weights1[8388] <= 16'b1111111111110111;
        weights1[8389] <= 16'b1111111111101100;
        weights1[8390] <= 16'b1111111111110101;
        weights1[8391] <= 16'b0000000000001110;
        weights1[8392] <= 16'b0000000000010100;
        weights1[8393] <= 16'b0000000000010110;
        weights1[8394] <= 16'b0000000000011000;
        weights1[8395] <= 16'b0000000000010000;
        weights1[8396] <= 16'b0000000000000101;
        weights1[8397] <= 16'b1111111111101100;
        weights1[8398] <= 16'b1111111111011101;
        weights1[8399] <= 16'b1111111111010110;
        weights1[8400] <= 16'b1111111111111100;
        weights1[8401] <= 16'b1111111111111000;
        weights1[8402] <= 16'b1111111111110010;
        weights1[8403] <= 16'b1111111111100000;
        weights1[8404] <= 16'b1111111111001110;
        weights1[8405] <= 16'b1111111111111011;
        weights1[8406] <= 16'b1111111111110011;
        weights1[8407] <= 16'b1111111111111000;
        weights1[8408] <= 16'b1111111111101011;
        weights1[8409] <= 16'b1111111111110110;
        weights1[8410] <= 16'b1111111111111011;
        weights1[8411] <= 16'b1111111111101110;
        weights1[8412] <= 16'b1111111111111111;
        weights1[8413] <= 16'b1111111111101100;
        weights1[8414] <= 16'b1111111111101101;
        weights1[8415] <= 16'b1111111111011010;
        weights1[8416] <= 16'b1111111111011111;
        weights1[8417] <= 16'b1111111111011111;
        weights1[8418] <= 16'b1111111111111001;
        weights1[8419] <= 16'b0000000000001001;
        weights1[8420] <= 16'b0000000000011001;
        weights1[8421] <= 16'b1111111111111010;
        weights1[8422] <= 16'b0000000000001111;
        weights1[8423] <= 16'b0000000000000100;
        weights1[8424] <= 16'b1111111111110101;
        weights1[8425] <= 16'b1111111111101101;
        weights1[8426] <= 16'b1111111111100001;
        weights1[8427] <= 16'b1111111111100001;
        weights1[8428] <= 16'b1111111111111100;
        weights1[8429] <= 16'b1111111111110101;
        weights1[8430] <= 16'b1111111111110000;
        weights1[8431] <= 16'b1111111111100100;
        weights1[8432] <= 16'b1111111111101100;
        weights1[8433] <= 16'b1111111111111110;
        weights1[8434] <= 16'b1111111111111010;
        weights1[8435] <= 16'b1111111111101010;
        weights1[8436] <= 16'b1111111111101110;
        weights1[8437] <= 16'b1111111111111000;
        weights1[8438] <= 16'b1111111111110111;
        weights1[8439] <= 16'b0000000000010000;
        weights1[8440] <= 16'b1111111111110001;
        weights1[8441] <= 16'b1111111111100111;
        weights1[8442] <= 16'b1111111111100100;
        weights1[8443] <= 16'b1111111111010101;
        weights1[8444] <= 16'b1111111111100101;
        weights1[8445] <= 16'b1111111111101010;
        weights1[8446] <= 16'b1111111111101110;
        weights1[8447] <= 16'b0000000000000011;
        weights1[8448] <= 16'b0000000000000100;
        weights1[8449] <= 16'b0000000000010000;
        weights1[8450] <= 16'b0000000000001110;
        weights1[8451] <= 16'b0000000000011011;
        weights1[8452] <= 16'b1111111111101100;
        weights1[8453] <= 16'b1111111111111111;
        weights1[8454] <= 16'b1111111111100101;
        weights1[8455] <= 16'b1111111111101011;
        weights1[8456] <= 16'b1111111111111101;
        weights1[8457] <= 16'b1111111111111010;
        weights1[8458] <= 16'b1111111111110011;
        weights1[8459] <= 16'b1111111111110111;
        weights1[8460] <= 16'b0000000000000100;
        weights1[8461] <= 16'b1111111111110001;
        weights1[8462] <= 16'b1111111111111100;
        weights1[8463] <= 16'b1111111111110100;
        weights1[8464] <= 16'b1111111111001010;
        weights1[8465] <= 16'b0000000000000001;
        weights1[8466] <= 16'b1111111111110000;
        weights1[8467] <= 16'b0000000000000011;
        weights1[8468] <= 16'b1111111111110001;
        weights1[8469] <= 16'b1111111111101111;
        weights1[8470] <= 16'b0000000000000000;
        weights1[8471] <= 16'b1111111111111111;
        weights1[8472] <= 16'b1111111111101001;
        weights1[8473] <= 16'b1111111111101111;
        weights1[8474] <= 16'b1111111111100001;
        weights1[8475] <= 16'b1111111111111010;
        weights1[8476] <= 16'b0000000000000001;
        weights1[8477] <= 16'b0000000000010011;
        weights1[8478] <= 16'b0000000000010101;
        weights1[8479] <= 16'b0000000000001001;
        weights1[8480] <= 16'b1111111111110111;
        weights1[8481] <= 16'b1111111111101011;
        weights1[8482] <= 16'b1111111111101010;
        weights1[8483] <= 16'b1111111111110100;
        weights1[8484] <= 16'b0000000000000000;
        weights1[8485] <= 16'b1111111111111011;
        weights1[8486] <= 16'b1111111111111110;
        weights1[8487] <= 16'b0000000000000001;
        weights1[8488] <= 16'b0000000000001101;
        weights1[8489] <= 16'b1111111111111110;
        weights1[8490] <= 16'b1111111111110000;
        weights1[8491] <= 16'b1111111111111011;
        weights1[8492] <= 16'b1111111111110011;
        weights1[8493] <= 16'b0000000000000110;
        weights1[8494] <= 16'b1111111111101101;
        weights1[8495] <= 16'b1111111111110000;
        weights1[8496] <= 16'b1111111111110111;
        weights1[8497] <= 16'b1111111111011101;
        weights1[8498] <= 16'b1111111111101100;
        weights1[8499] <= 16'b1111111111011101;
        weights1[8500] <= 16'b1111111111101111;
        weights1[8501] <= 16'b0000000000001101;
        weights1[8502] <= 16'b1111111111111110;
        weights1[8503] <= 16'b0000000000000001;
        weights1[8504] <= 16'b0000000000000010;
        weights1[8505] <= 16'b0000000000001001;
        weights1[8506] <= 16'b0000000000011010;
        weights1[8507] <= 16'b1111111111110010;
        weights1[8508] <= 16'b1111111111110100;
        weights1[8509] <= 16'b1111111111100101;
        weights1[8510] <= 16'b1111111111100101;
        weights1[8511] <= 16'b1111111111110010;
        weights1[8512] <= 16'b0000000000000000;
        weights1[8513] <= 16'b1111111111111101;
        weights1[8514] <= 16'b1111111111111011;
        weights1[8515] <= 16'b1111111111111100;
        weights1[8516] <= 16'b1111111111111110;
        weights1[8517] <= 16'b1111111111110101;
        weights1[8518] <= 16'b1111111111100111;
        weights1[8519] <= 16'b1111111111101011;
        weights1[8520] <= 16'b1111111111100010;
        weights1[8521] <= 16'b1111111111011101;
        weights1[8522] <= 16'b1111111111100101;
        weights1[8523] <= 16'b1111111111110100;
        weights1[8524] <= 16'b1111111111101100;
        weights1[8525] <= 16'b1111111111100000;
        weights1[8526] <= 16'b0000000000000001;
        weights1[8527] <= 16'b1111111111100110;
        weights1[8528] <= 16'b0000000000000011;
        weights1[8529] <= 16'b0000000000000111;
        weights1[8530] <= 16'b0000000000001001;
        weights1[8531] <= 16'b0000000000000011;
        weights1[8532] <= 16'b0000000000010000;
        weights1[8533] <= 16'b0000000000000000;
        weights1[8534] <= 16'b0000000000011000;
        weights1[8535] <= 16'b1111111111111101;
        weights1[8536] <= 16'b1111111111110001;
        weights1[8537] <= 16'b1111111111100010;
        weights1[8538] <= 16'b1111111111101100;
        weights1[8539] <= 16'b1111111111110111;
        weights1[8540] <= 16'b0000000000000000;
        weights1[8541] <= 16'b1111111111111111;
        weights1[8542] <= 16'b1111111111111011;
        weights1[8543] <= 16'b1111111111111001;
        weights1[8544] <= 16'b1111111111111100;
        weights1[8545] <= 16'b1111111111111100;
        weights1[8546] <= 16'b1111111111101110;
        weights1[8547] <= 16'b1111111111101001;
        weights1[8548] <= 16'b1111111111101100;
        weights1[8549] <= 16'b1111111111101000;
        weights1[8550] <= 16'b1111111111110001;
        weights1[8551] <= 16'b1111111111111110;
        weights1[8552] <= 16'b1111111111110101;
        weights1[8553] <= 16'b1111111111101100;
        weights1[8554] <= 16'b1111111111111100;
        weights1[8555] <= 16'b1111111111111000;
        weights1[8556] <= 16'b1111111111111011;
        weights1[8557] <= 16'b1111111111111001;
        weights1[8558] <= 16'b1111111111110110;
        weights1[8559] <= 16'b1111111111110110;
        weights1[8560] <= 16'b0000000000000011;
        weights1[8561] <= 16'b0000000000001100;
        weights1[8562] <= 16'b0000000000000110;
        weights1[8563] <= 16'b1111111111101110;
        weights1[8564] <= 16'b1111111111110001;
        weights1[8565] <= 16'b1111111111101010;
        weights1[8566] <= 16'b1111111111101111;
        weights1[8567] <= 16'b1111111111111110;
        weights1[8568] <= 16'b0000000000000000;
        weights1[8569] <= 16'b0000000000000000;
        weights1[8570] <= 16'b1111111111111100;
        weights1[8571] <= 16'b1111111111111011;
        weights1[8572] <= 16'b1111111111111010;
        weights1[8573] <= 16'b1111111111110001;
        weights1[8574] <= 16'b1111111111110110;
        weights1[8575] <= 16'b1111111111110110;
        weights1[8576] <= 16'b1111111111110101;
        weights1[8577] <= 16'b1111111111101111;
        weights1[8578] <= 16'b1111111111110011;
        weights1[8579] <= 16'b1111111111110000;
        weights1[8580] <= 16'b1111111111101011;
        weights1[8581] <= 16'b1111111111111010;
        weights1[8582] <= 16'b1111111111110100;
        weights1[8583] <= 16'b1111111111101001;
        weights1[8584] <= 16'b1111111111110110;
        weights1[8585] <= 16'b1111111111110001;
        weights1[8586] <= 16'b1111111111111000;
        weights1[8587] <= 16'b1111111111101101;
        weights1[8588] <= 16'b1111111111111110;
        weights1[8589] <= 16'b0000000000001010;
        weights1[8590] <= 16'b0000000000000000;
        weights1[8591] <= 16'b1111111111101100;
        weights1[8592] <= 16'b1111111111110000;
        weights1[8593] <= 16'b1111111111110110;
        weights1[8594] <= 16'b1111111111111010;
        weights1[8595] <= 16'b1111111111111111;
        weights1[8596] <= 16'b0000000000000000;
        weights1[8597] <= 16'b1111111111111110;
        weights1[8598] <= 16'b1111111111111110;
        weights1[8599] <= 16'b1111111111111100;
        weights1[8600] <= 16'b1111111111111010;
        weights1[8601] <= 16'b1111111111111001;
        weights1[8602] <= 16'b1111111111110101;
        weights1[8603] <= 16'b1111111111111000;
        weights1[8604] <= 16'b1111111111110110;
        weights1[8605] <= 16'b1111111111110111;
        weights1[8606] <= 16'b1111111111111010;
        weights1[8607] <= 16'b1111111111101100;
        weights1[8608] <= 16'b1111111111110101;
        weights1[8609] <= 16'b1111111111101111;
        weights1[8610] <= 16'b1111111111100010;
        weights1[8611] <= 16'b1111111111111100;
        weights1[8612] <= 16'b1111111111110000;
        weights1[8613] <= 16'b1111111111110110;
        weights1[8614] <= 16'b0000000000001011;
        weights1[8615] <= 16'b0000000000010010;
        weights1[8616] <= 16'b0000000000000111;
        weights1[8617] <= 16'b0000000000001111;
        weights1[8618] <= 16'b0000000000000000;
        weights1[8619] <= 16'b1111111111111111;
        weights1[8620] <= 16'b1111111111111100;
        weights1[8621] <= 16'b1111111111111101;
        weights1[8622] <= 16'b1111111111111101;
        weights1[8623] <= 16'b1111111111111111;
        weights1[8624] <= 16'b0000000000000000;
        weights1[8625] <= 16'b0000000000000000;
        weights1[8626] <= 16'b0000000000000000;
        weights1[8627] <= 16'b1111111111111110;
        weights1[8628] <= 16'b0000000000000010;
        weights1[8629] <= 16'b0000000000000011;
        weights1[8630] <= 16'b1111111111111110;
        weights1[8631] <= 16'b1111111111111101;
        weights1[8632] <= 16'b1111111111111010;
        weights1[8633] <= 16'b1111111111110101;
        weights1[8634] <= 16'b1111111111110000;
        weights1[8635] <= 16'b1111111111101011;
        weights1[8636] <= 16'b0000000000000011;
        weights1[8637] <= 16'b1111111111110100;
        weights1[8638] <= 16'b1111111111101111;
        weights1[8639] <= 16'b1111111111111011;
        weights1[8640] <= 16'b1111111111110111;
        weights1[8641] <= 16'b0000000000001000;
        weights1[8642] <= 16'b0000000000000001;
        weights1[8643] <= 16'b0000000000000011;
        weights1[8644] <= 16'b0000000000000101;
        weights1[8645] <= 16'b1111111111111111;
        weights1[8646] <= 16'b1111111111110110;
        weights1[8647] <= 16'b1111111111101101;
        weights1[8648] <= 16'b1111111111101110;
        weights1[8649] <= 16'b1111111111110100;
        weights1[8650] <= 16'b1111111111111001;
        weights1[8651] <= 16'b1111111111111100;
        weights1[8652] <= 16'b0000000000000000;
        weights1[8653] <= 16'b0000000000000001;
        weights1[8654] <= 16'b0000000000000100;
        weights1[8655] <= 16'b0000000000000100;
        weights1[8656] <= 16'b0000000000000111;
        weights1[8657] <= 16'b0000000000000100;
        weights1[8658] <= 16'b1111111111111010;
        weights1[8659] <= 16'b1111111111111101;
        weights1[8660] <= 16'b0000000000000110;
        weights1[8661] <= 16'b1111111111111011;
        weights1[8662] <= 16'b0000000000000110;
        weights1[8663] <= 16'b1111111111111111;
        weights1[8664] <= 16'b1111111111110110;
        weights1[8665] <= 16'b1111111111111011;
        weights1[8666] <= 16'b0000000000000010;
        weights1[8667] <= 16'b1111111111110111;
        weights1[8668] <= 16'b1111111111111010;
        weights1[8669] <= 16'b1111111111110111;
        weights1[8670] <= 16'b0000000000001100;
        weights1[8671] <= 16'b1111111111111110;
        weights1[8672] <= 16'b1111111111111001;
        weights1[8673] <= 16'b0000000000000011;
        weights1[8674] <= 16'b1111111111111000;
        weights1[8675] <= 16'b1111111111111011;
        weights1[8676] <= 16'b1111111111101100;
        weights1[8677] <= 16'b1111111111110111;
        weights1[8678] <= 16'b1111111111110111;
        weights1[8679] <= 16'b1111111111111110;
        weights1[8680] <= 16'b0000000000000001;
        weights1[8681] <= 16'b0000000000000100;
        weights1[8682] <= 16'b0000000000000111;
        weights1[8683] <= 16'b0000000000000110;
        weights1[8684] <= 16'b0000000000000111;
        weights1[8685] <= 16'b0000000000000010;
        weights1[8686] <= 16'b0000000000001000;
        weights1[8687] <= 16'b1111111111110000;
        weights1[8688] <= 16'b1111111111111101;
        weights1[8689] <= 16'b1111111111110111;
        weights1[8690] <= 16'b1111111111111101;
        weights1[8691] <= 16'b0000000000000001;
        weights1[8692] <= 16'b0000000000000000;
        weights1[8693] <= 16'b0000000000000110;
        weights1[8694] <= 16'b0000000000010010;
        weights1[8695] <= 16'b1111111111111000;
        weights1[8696] <= 16'b1111111111111010;
        weights1[8697] <= 16'b1111111111101110;
        weights1[8698] <= 16'b1111111111101110;
        weights1[8699] <= 16'b1111111111101100;
        weights1[8700] <= 16'b1111111111111111;
        weights1[8701] <= 16'b1111111111111001;
        weights1[8702] <= 16'b1111111111110110;
        weights1[8703] <= 16'b1111111111111101;
        weights1[8704] <= 16'b1111111111111011;
        weights1[8705] <= 16'b0000000000000000;
        weights1[8706] <= 16'b0000000000001000;
        weights1[8707] <= 16'b1111111111111111;
        weights1[8708] <= 16'b0000000000000100;
        weights1[8709] <= 16'b0000000000000111;
        weights1[8710] <= 16'b0000000000000001;
        weights1[8711] <= 16'b1111111111111001;
        weights1[8712] <= 16'b0000000000000001;
        weights1[8713] <= 16'b0000000000000000;
        weights1[8714] <= 16'b0000000000001000;
        weights1[8715] <= 16'b1111111111111100;
        weights1[8716] <= 16'b0000000000001000;
        weights1[8717] <= 16'b0000000000010000;
        weights1[8718] <= 16'b0000000000001101;
        weights1[8719] <= 16'b0000000000010000;
        weights1[8720] <= 16'b1111111111111100;
        weights1[8721] <= 16'b1111111111100010;
        weights1[8722] <= 16'b1111111111101100;
        weights1[8723] <= 16'b1111111111101011;
        weights1[8724] <= 16'b0000000000000011;
        weights1[8725] <= 16'b0000000000100000;
        weights1[8726] <= 16'b1111111111111100;
        weights1[8727] <= 16'b1111111111111111;
        weights1[8728] <= 16'b1111111111111010;
        weights1[8729] <= 16'b0000000000000000;
        weights1[8730] <= 16'b0000000000000001;
        weights1[8731] <= 16'b1111111111110100;
        weights1[8732] <= 16'b1111111111111110;
        weights1[8733] <= 16'b1111111111110111;
        weights1[8734] <= 16'b0000000000000000;
        weights1[8735] <= 16'b1111111111111100;
        weights1[8736] <= 16'b0000000000000110;
        weights1[8737] <= 16'b0000000000001010;
        weights1[8738] <= 16'b1111111111111100;
        weights1[8739] <= 16'b1111111111110100;
        weights1[8740] <= 16'b0000000000000010;
        weights1[8741] <= 16'b0000000000011000;
        weights1[8742] <= 16'b0000000000010010;
        weights1[8743] <= 16'b0000000000001011;
        weights1[8744] <= 16'b0000000000001000;
        weights1[8745] <= 16'b1111111111110101;
        weights1[8746] <= 16'b1111111111110111;
        weights1[8747] <= 16'b0000000000000001;
        weights1[8748] <= 16'b0000000000000011;
        weights1[8749] <= 16'b1111111111111011;
        weights1[8750] <= 16'b0000000000010001;
        weights1[8751] <= 16'b0000000000011010;
        weights1[8752] <= 16'b1111111111111101;
        weights1[8753] <= 16'b1111111111111001;
        weights1[8754] <= 16'b0000000000010111;
        weights1[8755] <= 16'b1111111111110011;
        weights1[8756] <= 16'b0000000000011101;
        weights1[8757] <= 16'b1111111111110000;
        weights1[8758] <= 16'b0000000000001111;
        weights1[8759] <= 16'b0000000000001010;
        weights1[8760] <= 16'b1111111111101011;
        weights1[8761] <= 16'b1111111111111001;
        weights1[8762] <= 16'b1111111111111111;
        weights1[8763] <= 16'b1111111111111011;
        weights1[8764] <= 16'b0000000000000011;
        weights1[8765] <= 16'b0000000000000110;
        weights1[8766] <= 16'b1111111111111101;
        weights1[8767] <= 16'b1111111111111011;
        weights1[8768] <= 16'b0000000000010010;
        weights1[8769] <= 16'b1111111111111011;
        weights1[8770] <= 16'b0000000000001111;
        weights1[8771] <= 16'b0000000000001100;
        weights1[8772] <= 16'b1111111111111110;
        weights1[8773] <= 16'b1111111111110111;
        weights1[8774] <= 16'b0000000000001100;
        weights1[8775] <= 16'b0000000000001110;
        weights1[8776] <= 16'b0000000000000110;
        weights1[8777] <= 16'b1111111111111110;
        weights1[8778] <= 16'b1111111111110001;
        weights1[8779] <= 16'b1111111111111010;
        weights1[8780] <= 16'b0000000000000000;
        weights1[8781] <= 16'b0000000000000000;
        weights1[8782] <= 16'b1111111111111101;
        weights1[8783] <= 16'b0000000000010100;
        weights1[8784] <= 16'b0000000000001110;
        weights1[8785] <= 16'b0000000000000010;
        weights1[8786] <= 16'b1111111111111001;
        weights1[8787] <= 16'b0000000000001001;
        weights1[8788] <= 16'b1111111111111110;
        weights1[8789] <= 16'b1111111111111110;
        weights1[8790] <= 16'b1111111111111010;
        weights1[8791] <= 16'b1111111111110110;
        weights1[8792] <= 16'b0000000000000001;
        weights1[8793] <= 16'b0000000000000101;
        weights1[8794] <= 16'b0000000000001001;
        weights1[8795] <= 16'b0000000000000110;
        weights1[8796] <= 16'b0000000000010010;
        weights1[8797] <= 16'b0000000000000000;
        weights1[8798] <= 16'b0000000000010101;
        weights1[8799] <= 16'b0000000000000001;
        weights1[8800] <= 16'b1111111111110001;
        weights1[8801] <= 16'b0000000000010011;
        weights1[8802] <= 16'b0000000000011101;
        weights1[8803] <= 16'b0000000000000111;
        weights1[8804] <= 16'b0000000000001010;
        weights1[8805] <= 16'b1111111111111011;
        weights1[8806] <= 16'b0000000000010111;
        weights1[8807] <= 16'b1111111111111101;
        weights1[8808] <= 16'b0000000000000110;
        weights1[8809] <= 16'b1111111111111010;
        weights1[8810] <= 16'b0000000000000001;
        weights1[8811] <= 16'b0000000000000000;
        weights1[8812] <= 16'b1111111111110010;
        weights1[8813] <= 16'b1111111111110110;
        weights1[8814] <= 16'b1111111111111001;
        weights1[8815] <= 16'b1111111111110110;
        weights1[8816] <= 16'b0000000000000100;
        weights1[8817] <= 16'b1111111111110111;
        weights1[8818] <= 16'b1111111111111111;
        weights1[8819] <= 16'b1111111111101110;
        weights1[8820] <= 16'b0000000000000110;
        weights1[8821] <= 16'b0000000000000000;
        weights1[8822] <= 16'b0000000000010010;
        weights1[8823] <= 16'b0000000000001100;
        weights1[8824] <= 16'b1111111111110110;
        weights1[8825] <= 16'b1111111111111101;
        weights1[8826] <= 16'b0000000000011001;
        weights1[8827] <= 16'b0000000000001101;
        weights1[8828] <= 16'b0000000000011110;
        weights1[8829] <= 16'b0000000000011111;
        weights1[8830] <= 16'b0000000000010100;
        weights1[8831] <= 16'b1111111111111100;
        weights1[8832] <= 16'b0000000000000111;
        weights1[8833] <= 16'b0000000000010111;
        weights1[8834] <= 16'b0000000000000101;
        weights1[8835] <= 16'b0000000000001111;
        weights1[8836] <= 16'b0000000000001111;
        weights1[8837] <= 16'b0000000000001110;
        weights1[8838] <= 16'b0000000000000000;
        weights1[8839] <= 16'b0000000000000100;
        weights1[8840] <= 16'b0000000000010011;
        weights1[8841] <= 16'b1111111111111101;
        weights1[8842] <= 16'b0000000000001010;
        weights1[8843] <= 16'b1111111111111011;
        weights1[8844] <= 16'b1111111111111100;
        weights1[8845] <= 16'b1111111111110111;
        weights1[8846] <= 16'b1111111111111010;
        weights1[8847] <= 16'b1111111111110011;
        weights1[8848] <= 16'b0000000000001100;
        weights1[8849] <= 16'b0000000000001001;
        weights1[8850] <= 16'b0000000000010101;
        weights1[8851] <= 16'b0000000000001111;
        weights1[8852] <= 16'b0000000000100100;
        weights1[8853] <= 16'b0000000000000011;
        weights1[8854] <= 16'b0000000000000111;
        weights1[8855] <= 16'b0000000000011100;
        weights1[8856] <= 16'b0000000000101010;
        weights1[8857] <= 16'b0000000000001110;
        weights1[8858] <= 16'b1111111111110110;
        weights1[8859] <= 16'b0000000000101110;
        weights1[8860] <= 16'b0000000000001010;
        weights1[8861] <= 16'b0000000000000000;
        weights1[8862] <= 16'b0000000000100100;
        weights1[8863] <= 16'b0000000000001101;
        weights1[8864] <= 16'b0000000000010001;
        weights1[8865] <= 16'b1111111111111110;
        weights1[8866] <= 16'b1111111111110010;
        weights1[8867] <= 16'b0000000000000100;
        weights1[8868] <= 16'b0000000000000101;
        weights1[8869] <= 16'b1111111111110111;
        weights1[8870] <= 16'b0000000000000101;
        weights1[8871] <= 16'b0000000000000111;
        weights1[8872] <= 16'b0000000000000100;
        weights1[8873] <= 16'b0000000000000111;
        weights1[8874] <= 16'b0000000000000100;
        weights1[8875] <= 16'b1111111111110001;
        weights1[8876] <= 16'b0000000000001011;
        weights1[8877] <= 16'b0000000000001100;
        weights1[8878] <= 16'b0000000000011001;
        weights1[8879] <= 16'b0000000000100100;
        weights1[8880] <= 16'b0000000000110000;
        weights1[8881] <= 16'b0000000000101011;
        weights1[8882] <= 16'b0000000000100011;
        weights1[8883] <= 16'b0000000000010111;
        weights1[8884] <= 16'b0000000000101000;
        weights1[8885] <= 16'b0000000000101101;
        weights1[8886] <= 16'b0000000000101011;
        weights1[8887] <= 16'b0000000000110111;
        weights1[8888] <= 16'b0000000000101110;
        weights1[8889] <= 16'b0000000000101011;
        weights1[8890] <= 16'b0000000000010100;
        weights1[8891] <= 16'b0000000000000111;
        weights1[8892] <= 16'b0000000000001101;
        weights1[8893] <= 16'b0000000000001100;
        weights1[8894] <= 16'b0000000000001110;
        weights1[8895] <= 16'b0000000000000111;
        weights1[8896] <= 16'b0000000000001100;
        weights1[8897] <= 16'b0000000000000111;
        weights1[8898] <= 16'b1111111111111100;
        weights1[8899] <= 16'b1111111111110000;
        weights1[8900] <= 16'b0000000000001001;
        weights1[8901] <= 16'b1111111111101101;
        weights1[8902] <= 16'b1111111111111110;
        weights1[8903] <= 16'b1111111111100111;
        weights1[8904] <= 16'b0000000000001100;
        weights1[8905] <= 16'b0000000000010111;
        weights1[8906] <= 16'b0000000000100110;
        weights1[8907] <= 16'b0000000000101011;
        weights1[8908] <= 16'b0000000000110001;
        weights1[8909] <= 16'b0000000001001111;
        weights1[8910] <= 16'b0000000000100100;
        weights1[8911] <= 16'b0000000000111110;
        weights1[8912] <= 16'b0000000001001101;
        weights1[8913] <= 16'b0000000001010100;
        weights1[8914] <= 16'b0000000000110110;
        weights1[8915] <= 16'b0000000000101110;
        weights1[8916] <= 16'b0000000000011110;
        weights1[8917] <= 16'b0000000000010011;
        weights1[8918] <= 16'b0000000000000010;
        weights1[8919] <= 16'b0000000000001000;
        weights1[8920] <= 16'b0000000000001110;
        weights1[8921] <= 16'b1111111111111111;
        weights1[8922] <= 16'b0000000000000010;
        weights1[8923] <= 16'b0000000000000001;
        weights1[8924] <= 16'b1111111111111010;
        weights1[8925] <= 16'b1111111111110001;
        weights1[8926] <= 16'b1111111111111010;
        weights1[8927] <= 16'b1111111111100110;
        weights1[8928] <= 16'b0000000000000000;
        weights1[8929] <= 16'b1111111111110010;
        weights1[8930] <= 16'b1111111111111011;
        weights1[8931] <= 16'b1111111111110100;
        weights1[8932] <= 16'b1111111111111101;
        weights1[8933] <= 16'b1111111111111101;
        weights1[8934] <= 16'b0000000000010100;
        weights1[8935] <= 16'b0000000000010001;
        weights1[8936] <= 16'b0000000000010000;
        weights1[8937] <= 16'b0000000000100110;
        weights1[8938] <= 16'b0000000000100100;
        weights1[8939] <= 16'b0000000000110001;
        weights1[8940] <= 16'b0000000000010000;
        weights1[8941] <= 16'b0000000000000010;
        weights1[8942] <= 16'b1111111111011011;
        weights1[8943] <= 16'b1111111111100111;
        weights1[8944] <= 16'b1111111111011111;
        weights1[8945] <= 16'b1111111111010110;
        weights1[8946] <= 16'b1111111111100010;
        weights1[8947] <= 16'b1111111111100010;
        weights1[8948] <= 16'b1111111111101000;
        weights1[8949] <= 16'b1111111111110101;
        weights1[8950] <= 16'b1111111111101101;
        weights1[8951] <= 16'b0000000000000101;
        weights1[8952] <= 16'b1111111111111001;
        weights1[8953] <= 16'b1111111111111001;
        weights1[8954] <= 16'b1111111111110010;
        weights1[8955] <= 16'b0000000000000001;
        weights1[8956] <= 16'b1111111111110001;
        weights1[8957] <= 16'b1111111111110011;
        weights1[8958] <= 16'b1111111111111000;
        weights1[8959] <= 16'b1111111111111111;
        weights1[8960] <= 16'b1111111111101101;
        weights1[8961] <= 16'b1111111111101000;
        weights1[8962] <= 16'b1111111111100101;
        weights1[8963] <= 16'b1111111111110100;
        weights1[8964] <= 16'b1111111111101011;
        weights1[8965] <= 16'b1111111111100101;
        weights1[8966] <= 16'b1111111111011010;
        weights1[8967] <= 16'b1111111110101111;
        weights1[8968] <= 16'b1111111110011001;
        weights1[8969] <= 16'b1111111101011001;
        weights1[8970] <= 16'b1111111101101001;
        weights1[8971] <= 16'b1111111101000110;
        weights1[8972] <= 16'b1111111101100011;
        weights1[8973] <= 16'b1111111110011101;
        weights1[8974] <= 16'b1111111110100011;
        weights1[8975] <= 16'b1111111111010010;
        weights1[8976] <= 16'b1111111111100010;
        weights1[8977] <= 16'b1111111111011100;
        weights1[8978] <= 16'b1111111111100001;
        weights1[8979] <= 16'b1111111111101111;
        weights1[8980] <= 16'b1111111111110110;
        weights1[8981] <= 16'b1111111111111110;
        weights1[8982] <= 16'b1111111111110000;
        weights1[8983] <= 16'b1111111111101111;
        weights1[8984] <= 16'b1111111111111000;
        weights1[8985] <= 16'b1111111111111101;
        weights1[8986] <= 16'b1111111111111010;
        weights1[8987] <= 16'b0000000000001011;
        weights1[8988] <= 16'b1111111111010100;
        weights1[8989] <= 16'b1111111110111000;
        weights1[8990] <= 16'b1111111110111000;
        weights1[8991] <= 16'b1111111110011101;
        weights1[8992] <= 16'b1111111110010000;
        weights1[8993] <= 16'b1111111110000010;
        weights1[8994] <= 16'b1111111101100011;
        weights1[8995] <= 16'b1111111011110011;
        weights1[8996] <= 16'b1111111010111001;
        weights1[8997] <= 16'b1111111011011110;
        weights1[8998] <= 16'b1111111100110100;
        weights1[8999] <= 16'b1111111110011011;
        weights1[9000] <= 16'b1111111111001100;
        weights1[9001] <= 16'b1111111111100010;
        weights1[9002] <= 16'b1111111111100010;
        weights1[9003] <= 16'b1111111111011001;
        weights1[9004] <= 16'b1111111111101111;
        weights1[9005] <= 16'b1111111111110100;
        weights1[9006] <= 16'b1111111111110101;
        weights1[9007] <= 16'b1111111111101000;
        weights1[9008] <= 16'b1111111111110001;
        weights1[9009] <= 16'b0000000000000100;
        weights1[9010] <= 16'b1111111111111011;
        weights1[9011] <= 16'b0000000000000111;
        weights1[9012] <= 16'b0000000000001111;
        weights1[9013] <= 16'b1111111111111001;
        weights1[9014] <= 16'b0000000000001011;
        weights1[9015] <= 16'b0000000000001011;
        weights1[9016] <= 16'b1111111110111100;
        weights1[9017] <= 16'b1111111110010110;
        weights1[9018] <= 16'b1111111110010000;
        weights1[9019] <= 16'b1111111101101100;
        weights1[9020] <= 16'b1111111101001011;
        weights1[9021] <= 16'b1111111100011111;
        weights1[9022] <= 16'b1111111100010010;
        weights1[9023] <= 16'b1111111100001000;
        weights1[9024] <= 16'b1111111101110111;
        weights1[9025] <= 16'b1111111111110010;
        weights1[9026] <= 16'b0000000000001111;
        weights1[9027] <= 16'b0000000000001011;
        weights1[9028] <= 16'b0000000000010001;
        weights1[9029] <= 16'b1111111111111001;
        weights1[9030] <= 16'b1111111111111111;
        weights1[9031] <= 16'b0000000000000010;
        weights1[9032] <= 16'b0000000000000110;
        weights1[9033] <= 16'b0000000000000000;
        weights1[9034] <= 16'b0000000000001001;
        weights1[9035] <= 16'b0000000000001011;
        weights1[9036] <= 16'b0000000000000100;
        weights1[9037] <= 16'b0000000000010011;
        weights1[9038] <= 16'b0000000000001111;
        weights1[9039] <= 16'b0000000000001011;
        weights1[9040] <= 16'b0000000000010010;
        weights1[9041] <= 16'b0000000000000101;
        weights1[9042] <= 16'b0000000000010110;
        weights1[9043] <= 16'b0000000000001101;
        weights1[9044] <= 16'b1111111110111011;
        weights1[9045] <= 16'b1111111110010010;
        weights1[9046] <= 16'b1111111110010001;
        weights1[9047] <= 16'b1111111101100001;
        weights1[9048] <= 16'b1111111101000111;
        weights1[9049] <= 16'b1111111101100011;
        weights1[9050] <= 16'b1111111110001011;
        weights1[9051] <= 16'b1111111111101110;
        weights1[9052] <= 16'b0000000000110000;
        weights1[9053] <= 16'b0000000000110100;
        weights1[9054] <= 16'b0000000001000011;
        weights1[9055] <= 16'b0000000000101011;
        weights1[9056] <= 16'b0000000000010110;
        weights1[9057] <= 16'b0000000000011110;
        weights1[9058] <= 16'b0000000000001101;
        weights1[9059] <= 16'b0000000000001001;
        weights1[9060] <= 16'b0000000000000010;
        weights1[9061] <= 16'b0000000000000011;
        weights1[9062] <= 16'b0000000000000000;
        weights1[9063] <= 16'b0000000000001101;
        weights1[9064] <= 16'b0000000000000110;
        weights1[9065] <= 16'b0000000000000000;
        weights1[9066] <= 16'b1111111111111011;
        weights1[9067] <= 16'b0000000000001110;
        weights1[9068] <= 16'b1111111111111111;
        weights1[9069] <= 16'b0000000000000101;
        weights1[9070] <= 16'b1111111111111110;
        weights1[9071] <= 16'b1111111111111110;
        weights1[9072] <= 16'b1111111111000011;
        weights1[9073] <= 16'b1111111110101100;
        weights1[9074] <= 16'b1111111110101111;
        weights1[9075] <= 16'b1111111110011101;
        weights1[9076] <= 16'b1111111110101011;
        weights1[9077] <= 16'b1111111111100000;
        weights1[9078] <= 16'b0000000000010101;
        weights1[9079] <= 16'b0000000001000100;
        weights1[9080] <= 16'b0000000000110111;
        weights1[9081] <= 16'b0000000000011010;
        weights1[9082] <= 16'b0000000000010110;
        weights1[9083] <= 16'b0000000000000101;
        weights1[9084] <= 16'b0000000000000011;
        weights1[9085] <= 16'b0000000000001001;
        weights1[9086] <= 16'b0000000000010000;
        weights1[9087] <= 16'b1111111111111101;
        weights1[9088] <= 16'b0000000000000011;
        weights1[9089] <= 16'b0000000000000110;
        weights1[9090] <= 16'b0000000000010001;
        weights1[9091] <= 16'b1111111111111010;
        weights1[9092] <= 16'b1111111111111101;
        weights1[9093] <= 16'b0000000000001100;
        weights1[9094] <= 16'b0000000000000110;
        weights1[9095] <= 16'b0000000000010101;
        weights1[9096] <= 16'b0000000000000000;
        weights1[9097] <= 16'b0000000000001010;
        weights1[9098] <= 16'b1111111111111111;
        weights1[9099] <= 16'b1111111111111111;
        weights1[9100] <= 16'b1111111111010000;
        weights1[9101] <= 16'b1111111111000110;
        weights1[9102] <= 16'b1111111111001100;
        weights1[9103] <= 16'b1111111111101010;
        weights1[9104] <= 16'b0000000000010010;
        weights1[9105] <= 16'b0000000000111010;
        weights1[9106] <= 16'b0000000001000110;
        weights1[9107] <= 16'b0000000000001000;
        weights1[9108] <= 16'b0000000000011010;
        weights1[9109] <= 16'b0000000000001111;
        weights1[9110] <= 16'b1111111111111001;
        weights1[9111] <= 16'b1111111111111011;
        weights1[9112] <= 16'b0000000000001001;
        weights1[9113] <= 16'b0000000000000010;
        weights1[9114] <= 16'b0000000000000010;
        weights1[9115] <= 16'b0000000000001010;
        weights1[9116] <= 16'b0000000000000111;
        weights1[9117] <= 16'b0000000000000110;
        weights1[9118] <= 16'b1111111111110111;
        weights1[9119] <= 16'b0000000000000111;
        weights1[9120] <= 16'b0000000000001111;
        weights1[9121] <= 16'b0000000000010011;
        weights1[9122] <= 16'b1111111111111010;
        weights1[9123] <= 16'b0000000000000101;
        weights1[9124] <= 16'b1111111111110000;
        weights1[9125] <= 16'b1111111111101111;
        weights1[9126] <= 16'b1111111111111010;
        weights1[9127] <= 16'b1111111111111101;
        weights1[9128] <= 16'b1111111111100011;
        weights1[9129] <= 16'b1111111111100000;
        weights1[9130] <= 16'b1111111111110011;
        weights1[9131] <= 16'b0000000000010001;
        weights1[9132] <= 16'b0000000000101001;
        weights1[9133] <= 16'b0000000000111010;
        weights1[9134] <= 16'b0000000000001101;
        weights1[9135] <= 16'b1111111111110101;
        weights1[9136] <= 16'b1111111111101100;
        weights1[9137] <= 16'b1111111111110001;
        weights1[9138] <= 16'b0000000000010011;
        weights1[9139] <= 16'b1111111111111001;
        weights1[9140] <= 16'b0000000000010000;
        weights1[9141] <= 16'b1111111111111110;
        weights1[9142] <= 16'b0000000000000001;
        weights1[9143] <= 16'b1111111111111001;
        weights1[9144] <= 16'b1111111111110001;
        weights1[9145] <= 16'b0000000000000110;
        weights1[9146] <= 16'b0000000000000100;
        weights1[9147] <= 16'b0000000000000101;
        weights1[9148] <= 16'b1111111111110100;
        weights1[9149] <= 16'b1111111111110001;
        weights1[9150] <= 16'b1111111111110000;
        weights1[9151] <= 16'b1111111111101001;
        weights1[9152] <= 16'b0000000000010011;
        weights1[9153] <= 16'b1111111111111110;
        weights1[9154] <= 16'b1111111111110110;
        weights1[9155] <= 16'b0000000000000011;
        weights1[9156] <= 16'b1111111111111100;
        weights1[9157] <= 16'b0000000000000100;
        weights1[9158] <= 16'b0000000000001011;
        weights1[9159] <= 16'b0000000000010110;
        weights1[9160] <= 16'b0000000000001100;
        weights1[9161] <= 16'b1111111111110110;
        weights1[9162] <= 16'b1111111111110000;
        weights1[9163] <= 16'b0000000000011001;
        weights1[9164] <= 16'b0000000000001100;
        weights1[9165] <= 16'b0000000000010001;
        weights1[9166] <= 16'b1111111111111111;
        weights1[9167] <= 16'b0000000000001010;
        weights1[9168] <= 16'b0000000000000011;
        weights1[9169] <= 16'b1111111111111111;
        weights1[9170] <= 16'b0000000000000001;
        weights1[9171] <= 16'b1111111111111010;
        weights1[9172] <= 16'b1111111111111111;
        weights1[9173] <= 16'b1111111111111100;
        weights1[9174] <= 16'b1111111111101000;
        weights1[9175] <= 16'b1111111111111011;
        weights1[9176] <= 16'b0000000000001000;
        weights1[9177] <= 16'b1111111111110010;
        weights1[9178] <= 16'b0000000000010111;
        weights1[9179] <= 16'b1111111111111011;
        weights1[9180] <= 16'b1111111111101011;
        weights1[9181] <= 16'b1111111111111011;
        weights1[9182] <= 16'b1111111111110011;
        weights1[9183] <= 16'b0000000000001001;
        weights1[9184] <= 16'b0000000000010101;
        weights1[9185] <= 16'b0000000000011101;
        weights1[9186] <= 16'b1111111111111111;
        weights1[9187] <= 16'b0000000000001010;
        weights1[9188] <= 16'b0000000000001100;
        weights1[9189] <= 16'b1111111111111010;
        weights1[9190] <= 16'b0000000000001110;
        weights1[9191] <= 16'b0000000000001100;
        weights1[9192] <= 16'b0000000000001010;
        weights1[9193] <= 16'b0000000000001110;
        weights1[9194] <= 16'b1111111111101010;
        weights1[9195] <= 16'b1111111111111110;
        weights1[9196] <= 16'b1111111111111110;
        weights1[9197] <= 16'b0000000000001001;
        weights1[9198] <= 16'b1111111111101101;
        weights1[9199] <= 16'b0000000000000100;
        weights1[9200] <= 16'b0000000000000000;
        weights1[9201] <= 16'b1111111111110101;
        weights1[9202] <= 16'b0000000000000100;
        weights1[9203] <= 16'b1111111111110001;
        weights1[9204] <= 16'b0000000000000001;
        weights1[9205] <= 16'b1111111111111000;
        weights1[9206] <= 16'b0000000000000100;
        weights1[9207] <= 16'b1111111111110001;
        weights1[9208] <= 16'b0000000000010000;
        weights1[9209] <= 16'b1111111111110001;
        weights1[9210] <= 16'b1111111111101101;
        weights1[9211] <= 16'b1111111111111100;
        weights1[9212] <= 16'b0000000000010010;
        weights1[9213] <= 16'b0000000000010001;
        weights1[9214] <= 16'b0000000000000001;
        weights1[9215] <= 16'b0000000000001100;
        weights1[9216] <= 16'b1111111111110111;
        weights1[9217] <= 16'b0000000000010010;
        weights1[9218] <= 16'b1111111111111100;
        weights1[9219] <= 16'b0000000000000100;
        weights1[9220] <= 16'b1111111111111000;
        weights1[9221] <= 16'b0000000000001001;
        weights1[9222] <= 16'b0000000000001001;
        weights1[9223] <= 16'b0000000000000000;
        weights1[9224] <= 16'b0000000000001010;
        weights1[9225] <= 16'b1111111111101001;
        weights1[9226] <= 16'b0000000000001011;
        weights1[9227] <= 16'b0000000000000100;
        weights1[9228] <= 16'b1111111111110110;
        weights1[9229] <= 16'b1111111111111100;
        weights1[9230] <= 16'b0000000000001000;
        weights1[9231] <= 16'b1111111111111001;
        weights1[9232] <= 16'b1111111111111100;
        weights1[9233] <= 16'b0000000000001101;
        weights1[9234] <= 16'b0000000000000111;
        weights1[9235] <= 16'b0000000000010001;
        weights1[9236] <= 16'b1111111111111101;
        weights1[9237] <= 16'b1111111111111100;
        weights1[9238] <= 16'b1111111111111001;
        weights1[9239] <= 16'b0000000000001000;
        weights1[9240] <= 16'b0000000000000101;
        weights1[9241] <= 16'b0000000000001110;
        weights1[9242] <= 16'b0000000000000110;
        weights1[9243] <= 16'b0000000000010011;
        weights1[9244] <= 16'b0000000000000111;
        weights1[9245] <= 16'b1111111111111100;
        weights1[9246] <= 16'b1111111111111010;
        weights1[9247] <= 16'b1111111111111100;
        weights1[9248] <= 16'b0000000000001010;
        weights1[9249] <= 16'b1111111111111100;
        weights1[9250] <= 16'b0000000000000111;
        weights1[9251] <= 16'b1111111111111110;
        weights1[9252] <= 16'b1111111111111111;
        weights1[9253] <= 16'b0000000000000100;
        weights1[9254] <= 16'b0000000000000001;
        weights1[9255] <= 16'b0000000000000001;
        weights1[9256] <= 16'b0000000000011100;
        weights1[9257] <= 16'b0000000000000001;
        weights1[9258] <= 16'b1111111111110110;
        weights1[9259] <= 16'b1111111111110111;
        weights1[9260] <= 16'b0000000000010101;
        weights1[9261] <= 16'b1111111111110110;
        weights1[9262] <= 16'b1111111111110110;
        weights1[9263] <= 16'b0000000000000001;
        weights1[9264] <= 16'b0000000000000100;
        weights1[9265] <= 16'b1111111111111100;
        weights1[9266] <= 16'b0000000000000000;
        weights1[9267] <= 16'b0000000000000110;
        weights1[9268] <= 16'b1111111111111110;
        weights1[9269] <= 16'b0000000000001011;
        weights1[9270] <= 16'b0000000000001000;
        weights1[9271] <= 16'b1111111111110111;
        weights1[9272] <= 16'b1111111111110110;
        weights1[9273] <= 16'b0000000000000110;
        weights1[9274] <= 16'b0000000000000011;
        weights1[9275] <= 16'b0000000000000000;
        weights1[9276] <= 16'b1111111111111101;
        weights1[9277] <= 16'b0000000000000110;
        weights1[9278] <= 16'b1111111111111101;
        weights1[9279] <= 16'b0000000000001101;
        weights1[9280] <= 16'b1111111111110110;
        weights1[9281] <= 16'b1111111111111101;
        weights1[9282] <= 16'b0000000000001010;
        weights1[9283] <= 16'b1111111111110001;
        weights1[9284] <= 16'b1111111111110111;
        weights1[9285] <= 16'b0000000000000110;
        weights1[9286] <= 16'b0000000000011101;
        weights1[9287] <= 16'b1111111111111100;
        weights1[9288] <= 16'b1111111111110001;
        weights1[9289] <= 16'b1111111111110010;
        weights1[9290] <= 16'b1111111111101011;
        weights1[9291] <= 16'b0000000000001000;
        weights1[9292] <= 16'b0000000000010101;
        weights1[9293] <= 16'b1111111111111101;
        weights1[9294] <= 16'b1111111111111110;
        weights1[9295] <= 16'b0000000000001010;
        weights1[9296] <= 16'b0000000000001011;
        weights1[9297] <= 16'b0000000000000010;
        weights1[9298] <= 16'b0000000000001010;
        weights1[9299] <= 16'b1111111111111111;
        weights1[9300] <= 16'b0000000000000100;
        weights1[9301] <= 16'b0000000000000100;
        weights1[9302] <= 16'b0000000000001110;
        weights1[9303] <= 16'b1111111111111000;
        weights1[9304] <= 16'b0000000000000010;
        weights1[9305] <= 16'b0000000000001010;
        weights1[9306] <= 16'b1111111111110010;
        weights1[9307] <= 16'b1111111111111001;
        weights1[9308] <= 16'b1111111111110010;
        weights1[9309] <= 16'b0000000000000010;
        weights1[9310] <= 16'b1111111111111100;
        weights1[9311] <= 16'b0000000000010001;
        weights1[9312] <= 16'b1111111111111110;
        weights1[9313] <= 16'b0000000000000100;
        weights1[9314] <= 16'b0000000000000011;
        weights1[9315] <= 16'b0000000000010000;
        weights1[9316] <= 16'b0000000000001000;
        weights1[9317] <= 16'b0000000000001000;
        weights1[9318] <= 16'b0000000000000000;
        weights1[9319] <= 16'b1111111111101110;
        weights1[9320] <= 16'b0000000000001101;
        weights1[9321] <= 16'b0000000000000100;
        weights1[9322] <= 16'b0000000000000110;
        weights1[9323] <= 16'b0000000000001000;
        weights1[9324] <= 16'b0000000000000110;
        weights1[9325] <= 16'b1111111111111111;
        weights1[9326] <= 16'b1111111111111110;
        weights1[9327] <= 16'b1111111111111011;
        weights1[9328] <= 16'b1111111111110111;
        weights1[9329] <= 16'b1111111111111010;
        weights1[9330] <= 16'b0000000000000100;
        weights1[9331] <= 16'b0000000000001000;
        weights1[9332] <= 16'b0000000000000111;
        weights1[9333] <= 16'b0000000000001100;
        weights1[9334] <= 16'b0000000000010011;
        weights1[9335] <= 16'b1111111111110111;
        weights1[9336] <= 16'b0000000000001100;
        weights1[9337] <= 16'b0000000000001010;
        weights1[9338] <= 16'b1111111111110111;
        weights1[9339] <= 16'b0000000000000000;
        weights1[9340] <= 16'b0000000000000101;
        weights1[9341] <= 16'b1111111111110110;
        weights1[9342] <= 16'b1111111111111101;
        weights1[9343] <= 16'b0000000000001010;
        weights1[9344] <= 16'b1111111111111100;
        weights1[9345] <= 16'b0000000000001001;
        weights1[9346] <= 16'b0000000000000110;
        weights1[9347] <= 16'b0000000000000110;
        weights1[9348] <= 16'b1111111111111010;
        weights1[9349] <= 16'b0000000000001011;
        weights1[9350] <= 16'b0000000000001010;
        weights1[9351] <= 16'b0000000000000110;
        weights1[9352] <= 16'b0000000000000001;
        weights1[9353] <= 16'b0000000000000010;
        weights1[9354] <= 16'b0000000000000000;
        weights1[9355] <= 16'b0000000000000011;
        weights1[9356] <= 16'b0000000000001011;
        weights1[9357] <= 16'b1111111111110011;
        weights1[9358] <= 16'b0000000000000100;
        weights1[9359] <= 16'b0000000000000001;
        weights1[9360] <= 16'b1111111111101111;
        weights1[9361] <= 16'b1111111111111011;
        weights1[9362] <= 16'b0000000000000010;
        weights1[9363] <= 16'b1111111111111100;
        weights1[9364] <= 16'b1111111111111101;
        weights1[9365] <= 16'b1111111111111111;
        weights1[9366] <= 16'b1111111111111111;
        weights1[9367] <= 16'b0000000000000010;
        weights1[9368] <= 16'b1111111111111110;
        weights1[9369] <= 16'b0000000000001001;
        weights1[9370] <= 16'b1111111111111001;
        weights1[9371] <= 16'b0000000000000011;
        weights1[9372] <= 16'b0000000000000100;
        weights1[9373] <= 16'b0000000000001100;
        weights1[9374] <= 16'b0000000000000011;
        weights1[9375] <= 16'b0000000000001000;
        weights1[9376] <= 16'b0000000000001000;
        weights1[9377] <= 16'b0000000000010001;
        weights1[9378] <= 16'b0000000000001001;
        weights1[9379] <= 16'b0000000000000011;
        weights1[9380] <= 16'b0000000000000110;
        weights1[9381] <= 16'b0000000000001000;
        weights1[9382] <= 16'b0000000000001101;
        weights1[9383] <= 16'b0000000000001100;
        weights1[9384] <= 16'b0000000000001010;
        weights1[9385] <= 16'b1111111111111110;
        weights1[9386] <= 16'b0000000000000100;
        weights1[9387] <= 16'b0000000000001100;
        weights1[9388] <= 16'b0000000000000101;
        weights1[9389] <= 16'b0000000000001001;
        weights1[9390] <= 16'b0000000000000010;
        weights1[9391] <= 16'b1111111111111011;
        weights1[9392] <= 16'b0000000000001010;
        weights1[9393] <= 16'b1111111111111100;
        weights1[9394] <= 16'b0000000000000001;
        weights1[9395] <= 16'b0000000000000011;
        weights1[9396] <= 16'b1111111111111100;
        weights1[9397] <= 16'b0000000000000010;
        weights1[9398] <= 16'b0000000000000101;
        weights1[9399] <= 16'b0000000000001001;
        weights1[9400] <= 16'b0000000000001110;
        weights1[9401] <= 16'b0000000000000101;
        weights1[9402] <= 16'b0000000000000111;
        weights1[9403] <= 16'b0000000000001101;
        weights1[9404] <= 16'b0000000000000111;
        weights1[9405] <= 16'b0000000000001000;
        weights1[9406] <= 16'b0000000000000110;
        weights1[9407] <= 16'b0000000000000100;
        weights1[9408] <= 16'b0000000000000000;
        weights1[9409] <= 16'b0000000000000010;
        weights1[9410] <= 16'b0000000000000011;
        weights1[9411] <= 16'b0000000000001000;
        weights1[9412] <= 16'b0000000000000011;
        weights1[9413] <= 16'b0000000000001100;
        weights1[9414] <= 16'b0000000000001111;
        weights1[9415] <= 16'b0000000000001001;
        weights1[9416] <= 16'b0000000000010101;
        weights1[9417] <= 16'b0000000000100001;
        weights1[9418] <= 16'b0000000000011111;
        weights1[9419] <= 16'b0000000000001110;
        weights1[9420] <= 16'b0000000000100001;
        weights1[9421] <= 16'b0000000000010111;
        weights1[9422] <= 16'b0000000000001101;
        weights1[9423] <= 16'b0000000000010100;
        weights1[9424] <= 16'b0000000000010101;
        weights1[9425] <= 16'b0000000000010000;
        weights1[9426] <= 16'b0000000000001011;
        weights1[9427] <= 16'b0000000000010001;
        weights1[9428] <= 16'b0000000000010011;
        weights1[9429] <= 16'b0000000000010000;
        weights1[9430] <= 16'b0000000000001000;
        weights1[9431] <= 16'b0000000000010100;
        weights1[9432] <= 16'b0000000000001001;
        weights1[9433] <= 16'b0000000000001011;
        weights1[9434] <= 16'b0000000000000110;
        weights1[9435] <= 16'b0000000000000101;
        weights1[9436] <= 16'b0000000000000001;
        weights1[9437] <= 16'b0000000000000101;
        weights1[9438] <= 16'b0000000000000111;
        weights1[9439] <= 16'b0000000000000110;
        weights1[9440] <= 16'b0000000000001000;
        weights1[9441] <= 16'b0000000000001110;
        weights1[9442] <= 16'b0000000000011101;
        weights1[9443] <= 16'b0000000000010001;
        weights1[9444] <= 16'b0000000000011000;
        weights1[9445] <= 16'b0000000000010110;
        weights1[9446] <= 16'b0000000000000111;
        weights1[9447] <= 16'b1111111111110010;
        weights1[9448] <= 16'b0000000000000111;
        weights1[9449] <= 16'b1111111111111110;
        weights1[9450] <= 16'b0000000000000011;
        weights1[9451] <= 16'b0000000000001010;
        weights1[9452] <= 16'b0000000000010001;
        weights1[9453] <= 16'b0000000000010011;
        weights1[9454] <= 16'b0000000000010110;
        weights1[9455] <= 16'b0000000000010010;
        weights1[9456] <= 16'b0000000000011010;
        weights1[9457] <= 16'b0000000000000100;
        weights1[9458] <= 16'b0000000000000101;
        weights1[9459] <= 16'b0000000000011011;
        weights1[9460] <= 16'b0000000000001011;
        weights1[9461] <= 16'b0000000000000111;
        weights1[9462] <= 16'b0000000000001011;
        weights1[9463] <= 16'b1111111111111010;
        weights1[9464] <= 16'b0000000000000111;
        weights1[9465] <= 16'b0000000000000111;
        weights1[9466] <= 16'b0000000000001010;
        weights1[9467] <= 16'b0000000000001001;
        weights1[9468] <= 16'b0000000000011011;
        weights1[9469] <= 16'b0000000000011111;
        weights1[9470] <= 16'b0000000000011111;
        weights1[9471] <= 16'b0000000000001011;
        weights1[9472] <= 16'b0000000000000111;
        weights1[9473] <= 16'b0000000000000011;
        weights1[9474] <= 16'b1111111111101101;
        weights1[9475] <= 16'b0000000000000011;
        weights1[9476] <= 16'b0000000000000110;
        weights1[9477] <= 16'b1111111111111110;
        weights1[9478] <= 16'b0000000000001000;
        weights1[9479] <= 16'b0000000000000111;
        weights1[9480] <= 16'b1111111111111001;
        weights1[9481] <= 16'b1111111111110010;
        weights1[9482] <= 16'b0000000000001110;
        weights1[9483] <= 16'b0000000000001100;
        weights1[9484] <= 16'b0000000000010001;
        weights1[9485] <= 16'b0000000000001111;
        weights1[9486] <= 16'b0000000000000010;
        weights1[9487] <= 16'b1111111111110100;
        weights1[9488] <= 16'b0000000000001010;
        weights1[9489] <= 16'b0000000000001010;
        weights1[9490] <= 16'b0000000000001001;
        weights1[9491] <= 16'b0000000000000110;
        weights1[9492] <= 16'b0000000000000010;
        weights1[9493] <= 16'b0000000000001101;
        weights1[9494] <= 16'b0000000000001011;
        weights1[9495] <= 16'b0000000000001111;
        weights1[9496] <= 16'b0000000000100000;
        weights1[9497] <= 16'b0000000000100000;
        weights1[9498] <= 16'b1111111111111111;
        weights1[9499] <= 16'b0000000000010011;
        weights1[9500] <= 16'b1111111111111100;
        weights1[9501] <= 16'b0000000000000011;
        weights1[9502] <= 16'b0000000000001010;
        weights1[9503] <= 16'b0000000000000110;
        weights1[9504] <= 16'b0000000000000001;
        weights1[9505] <= 16'b0000000000000111;
        weights1[9506] <= 16'b0000000000001010;
        weights1[9507] <= 16'b1111111111101011;
        weights1[9508] <= 16'b1111111111111101;
        weights1[9509] <= 16'b0000000000000110;
        weights1[9510] <= 16'b1111111111111100;
        weights1[9511] <= 16'b1111111111111111;
        weights1[9512] <= 16'b0000000000000011;
        weights1[9513] <= 16'b1111111111111100;
        weights1[9514] <= 16'b0000000000010000;
        weights1[9515] <= 16'b1111111111111001;
        weights1[9516] <= 16'b0000000000000110;
        weights1[9517] <= 16'b0000000000001011;
        weights1[9518] <= 16'b0000000000010101;
        weights1[9519] <= 16'b0000000000001110;
        weights1[9520] <= 16'b0000000000001000;
        weights1[9521] <= 16'b0000000000001101;
        weights1[9522] <= 16'b0000000000001110;
        weights1[9523] <= 16'b0000000000000111;
        weights1[9524] <= 16'b0000000000001101;
        weights1[9525] <= 16'b0000000000001100;
        weights1[9526] <= 16'b0000000000000011;
        weights1[9527] <= 16'b0000000000000000;
        weights1[9528] <= 16'b0000000000000110;
        weights1[9529] <= 16'b1111111111111110;
        weights1[9530] <= 16'b1111111111101011;
        weights1[9531] <= 16'b1111111111011110;
        weights1[9532] <= 16'b1111111111111101;
        weights1[9533] <= 16'b0000000000000101;
        weights1[9534] <= 16'b1111111111111110;
        weights1[9535] <= 16'b1111111111110010;
        weights1[9536] <= 16'b0000000000000000;
        weights1[9537] <= 16'b1111111111101101;
        weights1[9538] <= 16'b1111111111110110;
        weights1[9539] <= 16'b1111111111110111;
        weights1[9540] <= 16'b0000000000000011;
        weights1[9541] <= 16'b1111111111111010;
        weights1[9542] <= 16'b0000000000001010;
        weights1[9543] <= 16'b1111111111111010;
        weights1[9544] <= 16'b0000000000000001;
        weights1[9545] <= 16'b0000000000010110;
        weights1[9546] <= 16'b0000000000010001;
        weights1[9547] <= 16'b0000000000000101;
        weights1[9548] <= 16'b0000000000000010;
        weights1[9549] <= 16'b0000000000000010;
        weights1[9550] <= 16'b0000000000001000;
        weights1[9551] <= 16'b1111111111101100;
        weights1[9552] <= 16'b1111111111111011;
        weights1[9553] <= 16'b1111111111110100;
        weights1[9554] <= 16'b1111111111110100;
        weights1[9555] <= 16'b1111111111111011;
        weights1[9556] <= 16'b1111111111110111;
        weights1[9557] <= 16'b1111111111101101;
        weights1[9558] <= 16'b1111111111111000;
        weights1[9559] <= 16'b1111111111110100;
        weights1[9560] <= 16'b1111111111101100;
        weights1[9561] <= 16'b1111111111101100;
        weights1[9562] <= 16'b0000000000000001;
        weights1[9563] <= 16'b1111111111100000;
        weights1[9564] <= 16'b1111111111100111;
        weights1[9565] <= 16'b1111111111101101;
        weights1[9566] <= 16'b0000000000001001;
        weights1[9567] <= 16'b0000000000000010;
        weights1[9568] <= 16'b1111111111111000;
        weights1[9569] <= 16'b0000000000000111;
        weights1[9570] <= 16'b0000000000000000;
        weights1[9571] <= 16'b1111111111110000;
        weights1[9572] <= 16'b1111111111111101;
        weights1[9573] <= 16'b1111111111111110;
        weights1[9574] <= 16'b0000000000001100;
        weights1[9575] <= 16'b1111111111111101;
        weights1[9576] <= 16'b0000000000000100;
        weights1[9577] <= 16'b1111111111111100;
        weights1[9578] <= 16'b0000000000000001;
        weights1[9579] <= 16'b1111111111110000;
        weights1[9580] <= 16'b0000000000010010;
        weights1[9581] <= 16'b0000000000000101;
        weights1[9582] <= 16'b0000000000011111;
        weights1[9583] <= 16'b1111111111011111;
        weights1[9584] <= 16'b0000000000001011;
        weights1[9585] <= 16'b0000000000000110;
        weights1[9586] <= 16'b1111111111111111;
        weights1[9587] <= 16'b0000000000101000;
        weights1[9588] <= 16'b0000000000001011;
        weights1[9589] <= 16'b1111111111101100;
        weights1[9590] <= 16'b0000000000001001;
        weights1[9591] <= 16'b0000000000001000;
        weights1[9592] <= 16'b1111111111111010;
        weights1[9593] <= 16'b0000000000000110;
        weights1[9594] <= 16'b0000000000000010;
        weights1[9595] <= 16'b1111111111110010;
        weights1[9596] <= 16'b1111111111111111;
        weights1[9597] <= 16'b1111111111111110;
        weights1[9598] <= 16'b0000000000000010;
        weights1[9599] <= 16'b1111111111110111;
        weights1[9600] <= 16'b1111111111110101;
        weights1[9601] <= 16'b1111111111101011;
        weights1[9602] <= 16'b0000000000000010;
        weights1[9603] <= 16'b0000000000001001;
        weights1[9604] <= 16'b0000000000000010;
        weights1[9605] <= 16'b1111111111110101;
        weights1[9606] <= 16'b0000000000000001;
        weights1[9607] <= 16'b0000000000000100;
        weights1[9608] <= 16'b1111111111111010;
        weights1[9609] <= 16'b0000000000001010;
        weights1[9610] <= 16'b0000000000000111;
        weights1[9611] <= 16'b0000000000000010;
        weights1[9612] <= 16'b0000000000000110;
        weights1[9613] <= 16'b0000000000000111;
        weights1[9614] <= 16'b0000000000001000;
        weights1[9615] <= 16'b1111111111110000;
        weights1[9616] <= 16'b0000000000000101;
        weights1[9617] <= 16'b0000000000001110;
        weights1[9618] <= 16'b0000000000001001;
        weights1[9619] <= 16'b0000000000000010;
        weights1[9620] <= 16'b1111111111110100;
        weights1[9621] <= 16'b1111111111111001;
        weights1[9622] <= 16'b1111111111110111;
        weights1[9623] <= 16'b0000000000001111;
        weights1[9624] <= 16'b1111111111110111;
        weights1[9625] <= 16'b1111111111110111;
        weights1[9626] <= 16'b1111111111110001;
        weights1[9627] <= 16'b1111111111111111;
        weights1[9628] <= 16'b0000000000001001;
        weights1[9629] <= 16'b1111111111110111;
        weights1[9630] <= 16'b0000000000010000;
        weights1[9631] <= 16'b0000000000001111;
        weights1[9632] <= 16'b0000000000000010;
        weights1[9633] <= 16'b1111111111110110;
        weights1[9634] <= 16'b0000000000000010;
        weights1[9635] <= 16'b0000000000000100;
        weights1[9636] <= 16'b0000000000000001;
        weights1[9637] <= 16'b1111111111101111;
        weights1[9638] <= 16'b0000000000001001;
        weights1[9639] <= 16'b1111111111110111;
        weights1[9640] <= 16'b1111111111111011;
        weights1[9641] <= 16'b1111111111111011;
        weights1[9642] <= 16'b0000000000001101;
        weights1[9643] <= 16'b1111111111101111;
        weights1[9644] <= 16'b0000000000010000;
        weights1[9645] <= 16'b0000000000001000;
        weights1[9646] <= 16'b1111111111111100;
        weights1[9647] <= 16'b0000000000000101;
        weights1[9648] <= 16'b0000000000010100;
        weights1[9649] <= 16'b1111111111111100;
        weights1[9650] <= 16'b1111111111111100;
        weights1[9651] <= 16'b1111111111111110;
        weights1[9652] <= 16'b0000000000010110;
        weights1[9653] <= 16'b0000000000000000;
        weights1[9654] <= 16'b0000000000000100;
        weights1[9655] <= 16'b1111111111111111;
        weights1[9656] <= 16'b1111111111110111;
        weights1[9657] <= 16'b1111111111110100;
        weights1[9658] <= 16'b0000000000000001;
        weights1[9659] <= 16'b0000000000011000;
        weights1[9660] <= 16'b0000000000000100;
        weights1[9661] <= 16'b0000000000000000;
        weights1[9662] <= 16'b1111111111111010;
        weights1[9663] <= 16'b1111111111110101;
        weights1[9664] <= 16'b1111111111101000;
        weights1[9665] <= 16'b1111111111101010;
        weights1[9666] <= 16'b1111111111111110;
        weights1[9667] <= 16'b0000000000010000;
        weights1[9668] <= 16'b0000000000001001;
        weights1[9669] <= 16'b0000000000000010;
        weights1[9670] <= 16'b0000000000000000;
        weights1[9671] <= 16'b0000000000001011;
        weights1[9672] <= 16'b1111111111111111;
        weights1[9673] <= 16'b1111111111110011;
        weights1[9674] <= 16'b0000000000001111;
        weights1[9675] <= 16'b1111111111110100;
        weights1[9676] <= 16'b1111111111111101;
        weights1[9677] <= 16'b0000000000000000;
        weights1[9678] <= 16'b0000000000001000;
        weights1[9679] <= 16'b0000000000000101;
        weights1[9680] <= 16'b1111111111101110;
        weights1[9681] <= 16'b0000000000000001;
        weights1[9682] <= 16'b1111111111110111;
        weights1[9683] <= 16'b0000000000000010;
        weights1[9684] <= 16'b1111111111110001;
        weights1[9685] <= 16'b1111111111110100;
        weights1[9686] <= 16'b0000000000000001;
        weights1[9687] <= 16'b0000000000001000;
        weights1[9688] <= 16'b0000000000001000;
        weights1[9689] <= 16'b0000000000000111;
        weights1[9690] <= 16'b1111111111111100;
        weights1[9691] <= 16'b0000000000000111;
        weights1[9692] <= 16'b1111111111101001;
        weights1[9693] <= 16'b1111111111111000;
        weights1[9694] <= 16'b1111111111110110;
        weights1[9695] <= 16'b1111111111111001;
        weights1[9696] <= 16'b0000000000000010;
        weights1[9697] <= 16'b0000000000001101;
        weights1[9698] <= 16'b0000000000001101;
        weights1[9699] <= 16'b0000000000010001;
        weights1[9700] <= 16'b0000000000001100;
        weights1[9701] <= 16'b0000000000010110;
        weights1[9702] <= 16'b0000000000000000;
        weights1[9703] <= 16'b0000000000000111;
        weights1[9704] <= 16'b0000000000000011;
        weights1[9705] <= 16'b0000000000001100;
        weights1[9706] <= 16'b1111111111111111;
        weights1[9707] <= 16'b0000000000000011;
        weights1[9708] <= 16'b0000000000001110;
        weights1[9709] <= 16'b1111111111110110;
        weights1[9710] <= 16'b0000000000001010;
        weights1[9711] <= 16'b1111111111111000;
        weights1[9712] <= 16'b1111111111111101;
        weights1[9713] <= 16'b1111111111111100;
        weights1[9714] <= 16'b0000000000001001;
        weights1[9715] <= 16'b0000000000010100;
        weights1[9716] <= 16'b0000000000000000;
        weights1[9717] <= 16'b0000000000000001;
        weights1[9718] <= 16'b1111111111111100;
        weights1[9719] <= 16'b0000000000000110;
        weights1[9720] <= 16'b1111111111101010;
        weights1[9721] <= 16'b0000000000000100;
        weights1[9722] <= 16'b0000000000000001;
        weights1[9723] <= 16'b0000000000010110;
        weights1[9724] <= 16'b1111111111101110;
        weights1[9725] <= 16'b1111111111111001;
        weights1[9726] <= 16'b1111111111111010;
        weights1[9727] <= 16'b0000000000000000;
        weights1[9728] <= 16'b1111111111111111;
        weights1[9729] <= 16'b0000000000000011;
        weights1[9730] <= 16'b0000000000000110;
        weights1[9731] <= 16'b0000000000000001;
        weights1[9732] <= 16'b1111111111111001;
        weights1[9733] <= 16'b1111111111111000;
        weights1[9734] <= 16'b0000000000000000;
        weights1[9735] <= 16'b1111111111111010;
        weights1[9736] <= 16'b1111111111110101;
        weights1[9737] <= 16'b1111111111110100;
        weights1[9738] <= 16'b1111111111111001;
        weights1[9739] <= 16'b1111111111110101;
        weights1[9740] <= 16'b1111111111111101;
        weights1[9741] <= 16'b0000000000001000;
        weights1[9742] <= 16'b0000000000010101;
        weights1[9743] <= 16'b0000000000010100;
        weights1[9744] <= 16'b0000000000010010;
        weights1[9745] <= 16'b1111111111111001;
        weights1[9746] <= 16'b0000000000001101;
        weights1[9747] <= 16'b1111111111111000;
        weights1[9748] <= 16'b1111111111111101;
        weights1[9749] <= 16'b1111111111110010;
        weights1[9750] <= 16'b1111111111111011;
        weights1[9751] <= 16'b1111111111110100;
        weights1[9752] <= 16'b0000000000000010;
        weights1[9753] <= 16'b1111111111110100;
        weights1[9754] <= 16'b1111111111110010;
        weights1[9755] <= 16'b0000000000001010;
        weights1[9756] <= 16'b1111111111111010;
        weights1[9757] <= 16'b1111111111111110;
        weights1[9758] <= 16'b1111111111111011;
        weights1[9759] <= 16'b0000000000000001;
        weights1[9760] <= 16'b1111111111110101;
        weights1[9761] <= 16'b0000000000000101;
        weights1[9762] <= 16'b1111111111111101;
        weights1[9763] <= 16'b0000000000000111;
        weights1[9764] <= 16'b0000000000000100;
        weights1[9765] <= 16'b1111111111111011;
        weights1[9766] <= 16'b1111111111111100;
        weights1[9767] <= 16'b0000000000001100;
        weights1[9768] <= 16'b1111111111110010;
        weights1[9769] <= 16'b1111111111111110;
        weights1[9770] <= 16'b0000000000000011;
        weights1[9771] <= 16'b0000000000001000;
        weights1[9772] <= 16'b0000000000010111;
        weights1[9773] <= 16'b0000000000001001;
        weights1[9774] <= 16'b0000000000000101;
        weights1[9775] <= 16'b0000000000001110;
        weights1[9776] <= 16'b1111111111110110;
        weights1[9777] <= 16'b1111111111101011;
        weights1[9778] <= 16'b1111111111111011;
        weights1[9779] <= 16'b1111111111100000;
        weights1[9780] <= 16'b1111111111100110;
        weights1[9781] <= 16'b1111111111101100;
        weights1[9782] <= 16'b1111111111011001;
        weights1[9783] <= 16'b1111111111101000;
        weights1[9784] <= 16'b1111111111110100;
        weights1[9785] <= 16'b1111111111110010;
        weights1[9786] <= 16'b1111111111111100;
        weights1[9787] <= 16'b1111111111011111;
        weights1[9788] <= 16'b1111111111110110;
        weights1[9789] <= 16'b1111111111110001;
        weights1[9790] <= 16'b1111111111111111;
        weights1[9791] <= 16'b1111111111111100;
        weights1[9792] <= 16'b1111111111111110;
        weights1[9793] <= 16'b1111111111110111;
        weights1[9794] <= 16'b1111111111111000;
        weights1[9795] <= 16'b1111111111101000;
        weights1[9796] <= 16'b1111111111110101;
        weights1[9797] <= 16'b1111111111101010;
        weights1[9798] <= 16'b1111111111101010;
        weights1[9799] <= 16'b1111111111111100;
        weights1[9800] <= 16'b0000000000010000;
        weights1[9801] <= 16'b0000000000000011;
        weights1[9802] <= 16'b0000000000000010;
        weights1[9803] <= 16'b0000000000001000;
        weights1[9804] <= 16'b0000000000001100;
        weights1[9805] <= 16'b1111111111011000;
        weights1[9806] <= 16'b0000000000010011;
        weights1[9807] <= 16'b1111111111111011;
        weights1[9808] <= 16'b1111111111111010;
        weights1[9809] <= 16'b1111111111101111;
        weights1[9810] <= 16'b1111111111110101;
        weights1[9811] <= 16'b1111111111111101;
        weights1[9812] <= 16'b1111111111111010;
        weights1[9813] <= 16'b0000000000000100;
        weights1[9814] <= 16'b0000000000000110;
        weights1[9815] <= 16'b0000000000001111;
        weights1[9816] <= 16'b0000000000000010;
        weights1[9817] <= 16'b0000000000000101;
        weights1[9818] <= 16'b1111111111111101;
        weights1[9819] <= 16'b1111111111111011;
        weights1[9820] <= 16'b0000000000001101;
        weights1[9821] <= 16'b1111111111101101;
        weights1[9822] <= 16'b0000000000001001;
        weights1[9823] <= 16'b1111111111010101;
        weights1[9824] <= 16'b1111111111101100;
        weights1[9825] <= 16'b1111111111010001;
        weights1[9826] <= 16'b1111111111100101;
        weights1[9827] <= 16'b1111111111100110;
        weights1[9828] <= 16'b0000000000001011;
        weights1[9829] <= 16'b0000000000001010;
        weights1[9830] <= 16'b0000000000010100;
        weights1[9831] <= 16'b0000000000010001;
        weights1[9832] <= 16'b0000000000010011;
        weights1[9833] <= 16'b0000000000010011;
        weights1[9834] <= 16'b0000000000000111;
        weights1[9835] <= 16'b1111111111110110;
        weights1[9836] <= 16'b0000000000000111;
        weights1[9837] <= 16'b0000000000000000;
        weights1[9838] <= 16'b0000000000001100;
        weights1[9839] <= 16'b1111111111111111;
        weights1[9840] <= 16'b0000000000100000;
        weights1[9841] <= 16'b0000000000011001;
        weights1[9842] <= 16'b0000000000010011;
        weights1[9843] <= 16'b0000000000010000;
        weights1[9844] <= 16'b0000000000001111;
        weights1[9845] <= 16'b0000000000001110;
        weights1[9846] <= 16'b1111111111110101;
        weights1[9847] <= 16'b0000000000000010;
        weights1[9848] <= 16'b0000000000000101;
        weights1[9849] <= 16'b1111111111101101;
        weights1[9850] <= 16'b1111111111110010;
        weights1[9851] <= 16'b1111111111100111;
        weights1[9852] <= 16'b1111111111010001;
        weights1[9853] <= 16'b1111111111011111;
        weights1[9854] <= 16'b1111111111010111;
        weights1[9855] <= 16'b1111111111011011;
        weights1[9856] <= 16'b1111111111110111;
        weights1[9857] <= 16'b1111111111111011;
        weights1[9858] <= 16'b0000000000010110;
        weights1[9859] <= 16'b0000000000011101;
        weights1[9860] <= 16'b0000000000000001;
        weights1[9861] <= 16'b0000000000100111;
        weights1[9862] <= 16'b0000000000011111;
        weights1[9863] <= 16'b0000000000001000;
        weights1[9864] <= 16'b1111111111110111;
        weights1[9865] <= 16'b1111111111111001;
        weights1[9866] <= 16'b0000000000001100;
        weights1[9867] <= 16'b0000000000000101;
        weights1[9868] <= 16'b0000000000000110;
        weights1[9869] <= 16'b0000000000001101;
        weights1[9870] <= 16'b0000000000010100;
        weights1[9871] <= 16'b1111111111111111;
        weights1[9872] <= 16'b0000000000001011;
        weights1[9873] <= 16'b1111111111111100;
        weights1[9874] <= 16'b0000000000001111;
        weights1[9875] <= 16'b1111111111110001;
        weights1[9876] <= 16'b1111111111111010;
        weights1[9877] <= 16'b1111111111011000;
        weights1[9878] <= 16'b1111111111010110;
        weights1[9879] <= 16'b1111111111010111;
        weights1[9880] <= 16'b1111111111011111;
        weights1[9881] <= 16'b1111111111101001;
        weights1[9882] <= 16'b1111111111101111;
        weights1[9883] <= 16'b1111111111101101;
        weights1[9884] <= 16'b1111111111100011;
        weights1[9885] <= 16'b1111111111110001;
        weights1[9886] <= 16'b0000000000000011;
        weights1[9887] <= 16'b0000000000000110;
        weights1[9888] <= 16'b0000000000000100;
        weights1[9889] <= 16'b1111111111111111;
        weights1[9890] <= 16'b1111111111111011;
        weights1[9891] <= 16'b0000000000001000;
        weights1[9892] <= 16'b0000000000010011;
        weights1[9893] <= 16'b0000000000001111;
        weights1[9894] <= 16'b0000000000010011;
        weights1[9895] <= 16'b1111111111110110;
        weights1[9896] <= 16'b0000000000010111;
        weights1[9897] <= 16'b0000000000011100;
        weights1[9898] <= 16'b0000000000011110;
        weights1[9899] <= 16'b0000000000010001;
        weights1[9900] <= 16'b1111111111111110;
        weights1[9901] <= 16'b1111111111111111;
        weights1[9902] <= 16'b1111111111111100;
        weights1[9903] <= 16'b1111111111101110;
        weights1[9904] <= 16'b1111111111011111;
        weights1[9905] <= 16'b1111111111010101;
        weights1[9906] <= 16'b1111111111100101;
        weights1[9907] <= 16'b1111111111101010;
        weights1[9908] <= 16'b1111111111111111;
        weights1[9909] <= 16'b0000000000010011;
        weights1[9910] <= 16'b1111111111111001;
        weights1[9911] <= 16'b0000000000001100;
        weights1[9912] <= 16'b1111111111011011;
        weights1[9913] <= 16'b1111111111000111;
        weights1[9914] <= 16'b1111111111010101;
        weights1[9915] <= 16'b1111111111100011;
        weights1[9916] <= 16'b1111111111101010;
        weights1[9917] <= 16'b0000000000001100;
        weights1[9918] <= 16'b0000000000000110;
        weights1[9919] <= 16'b1111111111111011;
        weights1[9920] <= 16'b1111111111111100;
        weights1[9921] <= 16'b1111111111111101;
        weights1[9922] <= 16'b0000000000001100;
        weights1[9923] <= 16'b1111111111111100;
        weights1[9924] <= 16'b0000000000100011;
        weights1[9925] <= 16'b0000000000100000;
        weights1[9926] <= 16'b0000000000001000;
        weights1[9927] <= 16'b0000000000010111;
        weights1[9928] <= 16'b0000000000000111;
        weights1[9929] <= 16'b1111111111101011;
        weights1[9930] <= 16'b1111111111100010;
        weights1[9931] <= 16'b1111111111010011;
        weights1[9932] <= 16'b1111111111010111;
        weights1[9933] <= 16'b1111111111100101;
        weights1[9934] <= 16'b1111111111110000;
        weights1[9935] <= 16'b0000000000001010;
        weights1[9936] <= 16'b0000000000000010;
        weights1[9937] <= 16'b0000000000100000;
        weights1[9938] <= 16'b0000000000011001;
        weights1[9939] <= 16'b0000000000000100;
        weights1[9940] <= 16'b1111111111011000;
        weights1[9941] <= 16'b1111111111000011;
        weights1[9942] <= 16'b1111111110111110;
        weights1[9943] <= 16'b1111111110110010;
        weights1[9944] <= 16'b1111111110111010;
        weights1[9945] <= 16'b1111111111100000;
        weights1[9946] <= 16'b1111111111101111;
        weights1[9947] <= 16'b1111111111111000;
        weights1[9948] <= 16'b0000000000000101;
        weights1[9949] <= 16'b0000000000001001;
        weights1[9950] <= 16'b1111111111111001;
        weights1[9951] <= 16'b0000000000001010;
        weights1[9952] <= 16'b1111111111110010;
        weights1[9953] <= 16'b0000000000001010;
        weights1[9954] <= 16'b1111111111111100;
        weights1[9955] <= 16'b1111111111100001;
        weights1[9956] <= 16'b1111111111001110;
        weights1[9957] <= 16'b1111111111010010;
        weights1[9958] <= 16'b1111111111011011;
        weights1[9959] <= 16'b1111111111010111;
        weights1[9960] <= 16'b1111111111100010;
        weights1[9961] <= 16'b1111111111110100;
        weights1[9962] <= 16'b0000000000001011;
        weights1[9963] <= 16'b0000000000010101;
        weights1[9964] <= 16'b0000000000010001;
        weights1[9965] <= 16'b0000000000100001;
        weights1[9966] <= 16'b0000000000011000;
        weights1[9967] <= 16'b0000000000001010;
        weights1[9968] <= 16'b1111111111011000;
        weights1[9969] <= 16'b1111111110111011;
        weights1[9970] <= 16'b1111111110101110;
        weights1[9971] <= 16'b1111111110011101;
        weights1[9972] <= 16'b1111111110000111;
        weights1[9973] <= 16'b1111111110000100;
        weights1[9974] <= 16'b1111111101100001;
        weights1[9975] <= 16'b1111111101011101;
        weights1[9976] <= 16'b1111111101001111;
        weights1[9977] <= 16'b1111111101101101;
        weights1[9978] <= 16'b1111111110000100;
        weights1[9979] <= 16'b1111111101110010;
        weights1[9980] <= 16'b1111111101010100;
        weights1[9981] <= 16'b1111111101111011;
        weights1[9982] <= 16'b1111111110001000;
        weights1[9983] <= 16'b1111111110100000;
        weights1[9984] <= 16'b1111111111001000;
        weights1[9985] <= 16'b1111111111010101;
        weights1[9986] <= 16'b1111111111101011;
        weights1[9987] <= 16'b1111111111111101;
        weights1[9988] <= 16'b0000000000001111;
        weights1[9989] <= 16'b0000000000010010;
        weights1[9990] <= 16'b0000000000010100;
        weights1[9991] <= 16'b0000000000010111;
        weights1[9992] <= 16'b0000000000011001;
        weights1[9993] <= 16'b0000000000011001;
        weights1[9994] <= 16'b0000000000010010;
        weights1[9995] <= 16'b0000000000001100;
        weights1[9996] <= 16'b1111111111011111;
        weights1[9997] <= 16'b1111111111000101;
        weights1[9998] <= 16'b1111111110101011;
        weights1[9999] <= 16'b1111111110101010;
        weights1[10000] <= 16'b1111111110011110;
        weights1[10001] <= 16'b1111111110100010;
        weights1[10002] <= 16'b1111111110000100;
        weights1[10003] <= 16'b1111111101101101;
        weights1[10004] <= 16'b1111111100110010;
        weights1[10005] <= 16'b1111111100100111;
        weights1[10006] <= 16'b1111111100011100;
        weights1[10007] <= 16'b1111111011111001;
        weights1[10008] <= 16'b1111111100010001;
        weights1[10009] <= 16'b1111111101000010;
        weights1[10010] <= 16'b1111111110000001;
        weights1[10011] <= 16'b1111111110110100;
        weights1[10012] <= 16'b1111111111100001;
        weights1[10013] <= 16'b1111111111011101;
        weights1[10014] <= 16'b0000000000000011;
        weights1[10015] <= 16'b0000000000011100;
        weights1[10016] <= 16'b0000000000000100;
        weights1[10017] <= 16'b0000000000010110;
        weights1[10018] <= 16'b0000000000110000;
        weights1[10019] <= 16'b0000000000101000;
        weights1[10020] <= 16'b0000000000010101;
        weights1[10021] <= 16'b0000000000011000;
        weights1[10022] <= 16'b0000000000010010;
        weights1[10023] <= 16'b0000000000001011;
        weights1[10024] <= 16'b1111111111100111;
        weights1[10025] <= 16'b1111111111001101;
        weights1[10026] <= 16'b1111111111000011;
        weights1[10027] <= 16'b1111111111000100;
        weights1[10028] <= 16'b1111111110111101;
        weights1[10029] <= 16'b1111111110111000;
        weights1[10030] <= 16'b1111111110110101;
        weights1[10031] <= 16'b1111111111000001;
        weights1[10032] <= 16'b1111111110110011;
        weights1[10033] <= 16'b1111111110001001;
        weights1[10034] <= 16'b1111111110001001;
        weights1[10035] <= 16'b1111111110101011;
        weights1[10036] <= 16'b1111111110111110;
        weights1[10037] <= 16'b1111111111010100;
        weights1[10038] <= 16'b1111111111011111;
        weights1[10039] <= 16'b1111111111100000;
        weights1[10040] <= 16'b0000000000000000;
        weights1[10041] <= 16'b0000000000001100;
        weights1[10042] <= 16'b0000000000011101;
        weights1[10043] <= 16'b1111111111111101;
        weights1[10044] <= 16'b0000000000010010;
        weights1[10045] <= 16'b0000000000010000;
        weights1[10046] <= 16'b0000000000011010;
        weights1[10047] <= 16'b0000000000011001;
        weights1[10048] <= 16'b0000000000010011;
        weights1[10049] <= 16'b0000000000001101;
        weights1[10050] <= 16'b0000000000001010;
        weights1[10051] <= 16'b0000000000010010;
        weights1[10052] <= 16'b1111111111111010;
        weights1[10053] <= 16'b1111111111101000;
        weights1[10054] <= 16'b1111111111011101;
        weights1[10055] <= 16'b1111111111101000;
        weights1[10056] <= 16'b1111111111110010;
        weights1[10057] <= 16'b1111111111010111;
        weights1[10058] <= 16'b1111111111100010;
        weights1[10059] <= 16'b1111111111111101;
        weights1[10060] <= 16'b0000000000000001;
        weights1[10061] <= 16'b1111111111111101;
        weights1[10062] <= 16'b0000000000011000;
        weights1[10063] <= 16'b0000000000101000;
        weights1[10064] <= 16'b0000000001001010;
        weights1[10065] <= 16'b0000000001001001;
        weights1[10066] <= 16'b0000000000110100;
        weights1[10067] <= 16'b0000000001000001;
        weights1[10068] <= 16'b0000000000011010;
        weights1[10069] <= 16'b0000000000010010;
        weights1[10070] <= 16'b0000000000001111;
        weights1[10071] <= 16'b0000000000100110;
        weights1[10072] <= 16'b0000000000001101;
        weights1[10073] <= 16'b0000000000010010;
        weights1[10074] <= 16'b0000000000001100;
        weights1[10075] <= 16'b1111111111110001;
        weights1[10076] <= 16'b0000000000011101;
        weights1[10077] <= 16'b0000000000000111;
        weights1[10078] <= 16'b0000000000001011;
        weights1[10079] <= 16'b0000000000001100;
        weights1[10080] <= 16'b0000000000000001;
        weights1[10081] <= 16'b0000000000000111;
        weights1[10082] <= 16'b1111111111101101;
        weights1[10083] <= 16'b1111111111110101;
        weights1[10084] <= 16'b0000000000000011;
        weights1[10085] <= 16'b0000000000010010;
        weights1[10086] <= 16'b1111111111111101;
        weights1[10087] <= 16'b0000000000010010;
        weights1[10088] <= 16'b0000000000110100;
        weights1[10089] <= 16'b0000000001100011;
        weights1[10090] <= 16'b0000000001101110;
        weights1[10091] <= 16'b0000000010000100;
        weights1[10092] <= 16'b0000000001001000;
        weights1[10093] <= 16'b0000000000101000;
        weights1[10094] <= 16'b0000000000101111;
        weights1[10095] <= 16'b0000000000110111;
        weights1[10096] <= 16'b0000000000001010;
        weights1[10097] <= 16'b0000000000010011;
        weights1[10098] <= 16'b0000000000001111;
        weights1[10099] <= 16'b0000000000011101;
        weights1[10100] <= 16'b0000000000010011;
        weights1[10101] <= 16'b0000000000000000;
        weights1[10102] <= 16'b0000000000001011;
        weights1[10103] <= 16'b0000000000011000;
        weights1[10104] <= 16'b0000000000001100;
        weights1[10105] <= 16'b0000000000000010;
        weights1[10106] <= 16'b0000000000000010;
        weights1[10107] <= 16'b1111111111111111;
        weights1[10108] <= 16'b1111111111111111;
        weights1[10109] <= 16'b1111111111111111;
        weights1[10110] <= 16'b0000000000010010;
        weights1[10111] <= 16'b0000000000011011;
        weights1[10112] <= 16'b0000000000011011;
        weights1[10113] <= 16'b0000000000101101;
        weights1[10114] <= 16'b0000000001010010;
        weights1[10115] <= 16'b0000000001000100;
        weights1[10116] <= 16'b0000000001011111;
        weights1[10117] <= 16'b0000000000111111;
        weights1[10118] <= 16'b0000000001101100;
        weights1[10119] <= 16'b0000000000110000;
        weights1[10120] <= 16'b0000000000110100;
        weights1[10121] <= 16'b0000000000101001;
        weights1[10122] <= 16'b0000000000001110;
        weights1[10123] <= 16'b0000000000011001;
        weights1[10124] <= 16'b0000000000010001;
        weights1[10125] <= 16'b0000000000001110;
        weights1[10126] <= 16'b0000000000001111;
        weights1[10127] <= 16'b0000000000100011;
        weights1[10128] <= 16'b0000000000001010;
        weights1[10129] <= 16'b0000000000001011;
        weights1[10130] <= 16'b0000000000001111;
        weights1[10131] <= 16'b0000000000100000;
        weights1[10132] <= 16'b0000000000100001;
        weights1[10133] <= 16'b0000000000000001;
        weights1[10134] <= 16'b0000000000000111;
        weights1[10135] <= 16'b0000000000000010;
        weights1[10136] <= 16'b1111111111111101;
        weights1[10137] <= 16'b0000000000000111;
        weights1[10138] <= 16'b0000000000010011;
        weights1[10139] <= 16'b0000000000011011;
        weights1[10140] <= 16'b0000000000011101;
        weights1[10141] <= 16'b0000000000101100;
        weights1[10142] <= 16'b0000000001001111;
        weights1[10143] <= 16'b0000000001010110;
        weights1[10144] <= 16'b0000000001001000;
        weights1[10145] <= 16'b0000000000011001;
        weights1[10146] <= 16'b0000000000010101;
        weights1[10147] <= 16'b0000000000000111;
        weights1[10148] <= 16'b0000000000000100;
        weights1[10149] <= 16'b0000000000011001;
        weights1[10150] <= 16'b0000000000001001;
        weights1[10151] <= 16'b0000000000011000;
        weights1[10152] <= 16'b0000000000000110;
        weights1[10153] <= 16'b0000000000001001;
        weights1[10154] <= 16'b0000000000001111;
        weights1[10155] <= 16'b0000000000000010;
        weights1[10156] <= 16'b0000000000010000;
        weights1[10157] <= 16'b0000000000000010;
        weights1[10158] <= 16'b1111111111111110;
        weights1[10159] <= 16'b1111111111111011;
        weights1[10160] <= 16'b0000000000001001;
        weights1[10161] <= 16'b0000000000001011;
        weights1[10162] <= 16'b0000000000000100;
        weights1[10163] <= 16'b1111111111111111;
        weights1[10164] <= 16'b0000000000000011;
        weights1[10165] <= 16'b0000000000001101;
        weights1[10166] <= 16'b0000000000011000;
        weights1[10167] <= 16'b0000000000011111;
        weights1[10168] <= 16'b0000000000101010;
        weights1[10169] <= 16'b0000000000110111;
        weights1[10170] <= 16'b0000000000111110;
        weights1[10171] <= 16'b0000000001000001;
        weights1[10172] <= 16'b0000000000101010;
        weights1[10173] <= 16'b0000000000100100;
        weights1[10174] <= 16'b0000000000101011;
        weights1[10175] <= 16'b0000000000100110;
        weights1[10176] <= 16'b0000000000110010;
        weights1[10177] <= 16'b0000000000100000;
        weights1[10178] <= 16'b0000000000101000;
        weights1[10179] <= 16'b0000000000010011;
        weights1[10180] <= 16'b0000000000011000;
        weights1[10181] <= 16'b0000000000000111;
        weights1[10182] <= 16'b0000000000010111;
        weights1[10183] <= 16'b0000000000000111;
        weights1[10184] <= 16'b0000000000000001;
        weights1[10185] <= 16'b0000000000001010;
        weights1[10186] <= 16'b0000000000001110;
        weights1[10187] <= 16'b0000000000010011;
        weights1[10188] <= 16'b0000000000001000;
        weights1[10189] <= 16'b0000000000000110;
        weights1[10190] <= 16'b1111111111111100;
        weights1[10191] <= 16'b1111111111111100;
        weights1[10192] <= 16'b0000000000000001;
        weights1[10193] <= 16'b0000000000000000;
        weights1[10194] <= 16'b0000000000000010;
        weights1[10195] <= 16'b0000000000000100;
        weights1[10196] <= 16'b0000000000001010;
        weights1[10197] <= 16'b0000000000000101;
        weights1[10198] <= 16'b0000000000000111;
        weights1[10199] <= 16'b0000000000001011;
        weights1[10200] <= 16'b0000000000001101;
        weights1[10201] <= 16'b0000000000001010;
        weights1[10202] <= 16'b0000000000011101;
        weights1[10203] <= 16'b0000000000010011;
        weights1[10204] <= 16'b1111111111111110;
        weights1[10205] <= 16'b0000000000000001;
        weights1[10206] <= 16'b1111111111111110;
        weights1[10207] <= 16'b0000000000010000;
        weights1[10208] <= 16'b0000000000000101;
        weights1[10209] <= 16'b0000000000000011;
        weights1[10210] <= 16'b0000000000000010;
        weights1[10211] <= 16'b0000000000001100;
        weights1[10212] <= 16'b0000000000000001;
        weights1[10213] <= 16'b0000000000000110;
        weights1[10214] <= 16'b1111111111111100;
        weights1[10215] <= 16'b0000000000010101;
        weights1[10216] <= 16'b0000000000010000;
        weights1[10217] <= 16'b0000000000001011;
        weights1[10218] <= 16'b0000000000000100;
        weights1[10219] <= 16'b0000000000000010;
        weights1[10220] <= 16'b0000000000000001;
        weights1[10221] <= 16'b0000000000000001;
        weights1[10222] <= 16'b0000000000000100;
        weights1[10223] <= 16'b0000000000000100;
        weights1[10224] <= 16'b0000000000010010;
        weights1[10225] <= 16'b0000000000010010;
        weights1[10226] <= 16'b0000000000010011;
        weights1[10227] <= 16'b0000000000000011;
        weights1[10228] <= 16'b0000000000000010;
        weights1[10229] <= 16'b0000000000001101;
        weights1[10230] <= 16'b0000000000001001;
        weights1[10231] <= 16'b1111111111111110;
        weights1[10232] <= 16'b0000000000001100;
        weights1[10233] <= 16'b0000000000001100;
        weights1[10234] <= 16'b1111111111111101;
        weights1[10235] <= 16'b0000000000000000;
        weights1[10236] <= 16'b0000000000001010;
        weights1[10237] <= 16'b0000000000000100;
        weights1[10238] <= 16'b1111111111110111;
        weights1[10239] <= 16'b0000000000001001;
        weights1[10240] <= 16'b0000000000000110;
        weights1[10241] <= 16'b1111111111111111;
        weights1[10242] <= 16'b0000000000000110;
        weights1[10243] <= 16'b0000000000000010;
        weights1[10244] <= 16'b0000000000001010;
        weights1[10245] <= 16'b0000000000000010;
        weights1[10246] <= 16'b1111111111111111;
        weights1[10247] <= 16'b0000000000000001;
        weights1[10248] <= 16'b0000000000000010;
        weights1[10249] <= 16'b0000000000000101;
        weights1[10250] <= 16'b0000000000000100;
        weights1[10251] <= 16'b0000000000000100;
        weights1[10252] <= 16'b0000000000000101;
        weights1[10253] <= 16'b1111111111111011;
        weights1[10254] <= 16'b0000000000010000;
        weights1[10255] <= 16'b0000000000010111;
        weights1[10256] <= 16'b0000000000001010;
        weights1[10257] <= 16'b0000000000011000;
        weights1[10258] <= 16'b0000000000010011;
        weights1[10259] <= 16'b0000000000001010;
        weights1[10260] <= 16'b0000000000001010;
        weights1[10261] <= 16'b0000000000000101;
        weights1[10262] <= 16'b0000000000000001;
        weights1[10263] <= 16'b0000000000001000;
        weights1[10264] <= 16'b0000000000001000;
        weights1[10265] <= 16'b1111111111111111;
        weights1[10266] <= 16'b1111111111111000;
        weights1[10267] <= 16'b0000000000000111;
        weights1[10268] <= 16'b0000000000000011;
        weights1[10269] <= 16'b0000000000001010;
        weights1[10270] <= 16'b0000000000000001;
        weights1[10271] <= 16'b1111111111111011;
        weights1[10272] <= 16'b1111111111111100;
        weights1[10273] <= 16'b0000000000000001;
        weights1[10274] <= 16'b0000000000000101;
        weights1[10275] <= 16'b0000000000000111;
        weights1[10276] <= 16'b0000000000000011;
        weights1[10277] <= 16'b0000000000000111;
        weights1[10278] <= 16'b0000000000001101;
        weights1[10279] <= 16'b0000000000001011;
        weights1[10280] <= 16'b0000000000000101;
        weights1[10281] <= 16'b0000000000001111;
        weights1[10282] <= 16'b0000000000001010;
        weights1[10283] <= 16'b0000000000010001;
        weights1[10284] <= 16'b1111111111111001;
        weights1[10285] <= 16'b1111111111110111;
        weights1[10286] <= 16'b0000000000000000;
        weights1[10287] <= 16'b0000000000010100;
        weights1[10288] <= 16'b0000000000000100;
        weights1[10289] <= 16'b1111111111101111;
        weights1[10290] <= 16'b0000000000001010;
        weights1[10291] <= 16'b0000000000000100;
        weights1[10292] <= 16'b1111111111110110;
        weights1[10293] <= 16'b0000000000000001;
        weights1[10294] <= 16'b1111111111110100;
        weights1[10295] <= 16'b1111111111110111;
        weights1[10296] <= 16'b0000000000001001;
        weights1[10297] <= 16'b0000000000000010;
        weights1[10298] <= 16'b1111111111111101;
        weights1[10299] <= 16'b0000000000001101;
        weights1[10300] <= 16'b1111111111111011;
        weights1[10301] <= 16'b0000000000001101;
        weights1[10302] <= 16'b0000000000001111;
        weights1[10303] <= 16'b0000000000001101;
        weights1[10304] <= 16'b0000000000000111;
        weights1[10305] <= 16'b0000000000001000;
        weights1[10306] <= 16'b0000000000010010;
        weights1[10307] <= 16'b0000000000000001;
        weights1[10308] <= 16'b0000000000000001;
        weights1[10309] <= 16'b0000000000000010;
        weights1[10310] <= 16'b1111111111101110;
        weights1[10311] <= 16'b0000000000001101;
        weights1[10312] <= 16'b0000000000000111;
        weights1[10313] <= 16'b1111111111101111;
        weights1[10314] <= 16'b0000000000000001;
        weights1[10315] <= 16'b1111111111110111;
        weights1[10316] <= 16'b0000000000000011;
        weights1[10317] <= 16'b0000000000001000;
        weights1[10318] <= 16'b0000000000000101;
        weights1[10319] <= 16'b0000000000000010;
        weights1[10320] <= 16'b0000000000001001;
        weights1[10321] <= 16'b0000000000000101;
        weights1[10322] <= 16'b0000000000010011;
        weights1[10323] <= 16'b0000000000010001;
        weights1[10324] <= 16'b1111111111111110;
        weights1[10325] <= 16'b0000000000000001;
        weights1[10326] <= 16'b1111111111111001;
        weights1[10327] <= 16'b1111111111111011;
        weights1[10328] <= 16'b0000000000001100;
        weights1[10329] <= 16'b0000000000000100;
        weights1[10330] <= 16'b1111111111111111;
        weights1[10331] <= 16'b0000000000000100;
        weights1[10332] <= 16'b0000000000001001;
        weights1[10333] <= 16'b0000000000001010;
        weights1[10334] <= 16'b0000000000010001;
        weights1[10335] <= 16'b0000000000000010;
        weights1[10336] <= 16'b1111111111111110;
        weights1[10337] <= 16'b0000000000000010;
        weights1[10338] <= 16'b1111111111111100;
        weights1[10339] <= 16'b1111111111111010;
        weights1[10340] <= 16'b0000000000000100;
        weights1[10341] <= 16'b0000000000000001;
        weights1[10342] <= 16'b0000000000000011;
        weights1[10343] <= 16'b0000000000000011;
        weights1[10344] <= 16'b0000000000010011;
        weights1[10345] <= 16'b0000000000000011;
        weights1[10346] <= 16'b1111111111111011;
        weights1[10347] <= 16'b0000000000000010;
        weights1[10348] <= 16'b0000000000001100;
        weights1[10349] <= 16'b1111111111110110;
        weights1[10350] <= 16'b1111111111110001;
        weights1[10351] <= 16'b0000000000000100;
        weights1[10352] <= 16'b1111111111111101;
        weights1[10353] <= 16'b1111111111111111;
        weights1[10354] <= 16'b1111111111100001;
        weights1[10355] <= 16'b0000000000100110;
        weights1[10356] <= 16'b0000000000000001;
        weights1[10357] <= 16'b1111111111101001;
        weights1[10358] <= 16'b1111111111110010;
        weights1[10359] <= 16'b0000000000000110;
        weights1[10360] <= 16'b0000000000000111;
        weights1[10361] <= 16'b0000000000000011;
        weights1[10362] <= 16'b0000000000000010;
        weights1[10363] <= 16'b0000000000000101;
        weights1[10364] <= 16'b1111111111101100;
        weights1[10365] <= 16'b1111111111101101;
        weights1[10366] <= 16'b0000000000001010;
        weights1[10367] <= 16'b1111111111101100;
        weights1[10368] <= 16'b1111111111111111;
        weights1[10369] <= 16'b1111111111111110;
        weights1[10370] <= 16'b0000000000000010;
        weights1[10371] <= 16'b0000000000001100;
        weights1[10372] <= 16'b1111111111101100;
        weights1[10373] <= 16'b1111111111111001;
        weights1[10374] <= 16'b1111111111111110;
        weights1[10375] <= 16'b1111111111111011;
        weights1[10376] <= 16'b0000000000001011;
        weights1[10377] <= 16'b1111111111111110;
        weights1[10378] <= 16'b0000000000010000;
        weights1[10379] <= 16'b0000000000000100;
        weights1[10380] <= 16'b0000000000000011;
        weights1[10381] <= 16'b0000000000000110;
        weights1[10382] <= 16'b0000000000000101;
        weights1[10383] <= 16'b1111111111110100;
        weights1[10384] <= 16'b1111111111111001;
        weights1[10385] <= 16'b1111111111110011;
        weights1[10386] <= 16'b0000000000010101;
        weights1[10387] <= 16'b0000000000000111;
        weights1[10388] <= 16'b1111111111111110;
        weights1[10389] <= 16'b1111111111110111;
        weights1[10390] <= 16'b1111111111110000;
        weights1[10391] <= 16'b1111111111101101;
        weights1[10392] <= 16'b1111111111110101;
        weights1[10393] <= 16'b0000000000001101;
        weights1[10394] <= 16'b1111111111101111;
        weights1[10395] <= 16'b0000000000010110;
        weights1[10396] <= 16'b1111111111111100;
        weights1[10397] <= 16'b1111111111110010;
        weights1[10398] <= 16'b1111111111110110;
        weights1[10399] <= 16'b0000000000001111;
        weights1[10400] <= 16'b0000000000010000;
        weights1[10401] <= 16'b0000000000000110;
        weights1[10402] <= 16'b0000000000010101;
        weights1[10403] <= 16'b0000000000001000;
        weights1[10404] <= 16'b0000000000001000;
        weights1[10405] <= 16'b0000000000011010;
        weights1[10406] <= 16'b0000000000001010;
        weights1[10407] <= 16'b0000000000010001;
        weights1[10408] <= 16'b0000000000001110;
        weights1[10409] <= 16'b1111111111111101;
        weights1[10410] <= 16'b0000000000000100;
        weights1[10411] <= 16'b0000000000000010;
        weights1[10412] <= 16'b0000000000000111;
        weights1[10413] <= 16'b1111111111111100;
        weights1[10414] <= 16'b1111111111110111;
        weights1[10415] <= 16'b0000000000000101;
        weights1[10416] <= 16'b1111111111111110;
        weights1[10417] <= 16'b1111111111110001;
        weights1[10418] <= 16'b0000000000000001;
        weights1[10419] <= 16'b1111111111101001;
        weights1[10420] <= 16'b1111111111111001;
        weights1[10421] <= 16'b0000000000000011;
        weights1[10422] <= 16'b1111111111110111;
        weights1[10423] <= 16'b1111111111110111;
        weights1[10424] <= 16'b1111111111110100;
        weights1[10425] <= 16'b0000000000001000;
        weights1[10426] <= 16'b1111111111111111;
        weights1[10427] <= 16'b0000000000000110;
        weights1[10428] <= 16'b0000000000000101;
        weights1[10429] <= 16'b1111111111111000;
        weights1[10430] <= 16'b0000000000000101;
        weights1[10431] <= 16'b0000000000000101;
        weights1[10432] <= 16'b0000000000001010;
        weights1[10433] <= 16'b1111111111111100;
        weights1[10434] <= 16'b1111111111111011;
        weights1[10435] <= 16'b0000000000000010;
        weights1[10436] <= 16'b0000000000001111;
        weights1[10437] <= 16'b0000000000010011;
        weights1[10438] <= 16'b0000000000001011;
        weights1[10439] <= 16'b0000000000010000;
        weights1[10440] <= 16'b0000000000011000;
        weights1[10441] <= 16'b0000000000000101;
        weights1[10442] <= 16'b1111111111111000;
        weights1[10443] <= 16'b0000000000000011;
        weights1[10444] <= 16'b1111111111110110;
        weights1[10445] <= 16'b1111111111101011;
        weights1[10446] <= 16'b1111111111101011;
        weights1[10447] <= 16'b1111111111110001;
        weights1[10448] <= 16'b0000000000000000;
        weights1[10449] <= 16'b0000000000001100;
        weights1[10450] <= 16'b0000000000000000;
        weights1[10451] <= 16'b0000000000001101;
        weights1[10452] <= 16'b0000000000010101;
        weights1[10453] <= 16'b0000000000001110;
        weights1[10454] <= 16'b1111111111110110;
        weights1[10455] <= 16'b0000000000000101;
        weights1[10456] <= 16'b0000000000000100;
        weights1[10457] <= 16'b0000000000001101;
        weights1[10458] <= 16'b1111111111111111;
        weights1[10459] <= 16'b0000000000000100;
        weights1[10460] <= 16'b1111111111111101;
        weights1[10461] <= 16'b0000000000000011;
        weights1[10462] <= 16'b1111111111111101;
        weights1[10463] <= 16'b0000000000000000;
        weights1[10464] <= 16'b0000000000001000;
        weights1[10465] <= 16'b0000000000010101;
        weights1[10466] <= 16'b0000000000010011;
        weights1[10467] <= 16'b0000000000001100;
        weights1[10468] <= 16'b0000000000000001;
        weights1[10469] <= 16'b0000000000001010;
        weights1[10470] <= 16'b0000000000000010;
        weights1[10471] <= 16'b0000000000000111;
        weights1[10472] <= 16'b1111111111101111;
        weights1[10473] <= 16'b1111111111100111;
        weights1[10474] <= 16'b1111111111011111;
        weights1[10475] <= 16'b1111111111110000;
        weights1[10476] <= 16'b0000000000000110;
        weights1[10477] <= 16'b1111111111110100;
        weights1[10478] <= 16'b1111111111111010;
        weights1[10479] <= 16'b0000000000000111;
        weights1[10480] <= 16'b0000000000000100;
        weights1[10481] <= 16'b1111111111101000;
        weights1[10482] <= 16'b0000000000001100;
        weights1[10483] <= 16'b1111111111110011;
        weights1[10484] <= 16'b1111111111100111;
        weights1[10485] <= 16'b1111111111111110;
        weights1[10486] <= 16'b1111111111110010;
        weights1[10487] <= 16'b1111111111111010;
        weights1[10488] <= 16'b1111111111111000;
        weights1[10489] <= 16'b1111111111111110;
        weights1[10490] <= 16'b1111111111111101;
        weights1[10491] <= 16'b1111111111101000;
        weights1[10492] <= 16'b1111111111111101;
        weights1[10493] <= 16'b1111111111111001;
        weights1[10494] <= 16'b1111111111101011;
        weights1[10495] <= 16'b0000000000000110;
        weights1[10496] <= 16'b1111111111111000;
        weights1[10497] <= 16'b0000000000001101;
        weights1[10498] <= 16'b0000000000010101;
        weights1[10499] <= 16'b0000000000001111;
        weights1[10500] <= 16'b1111111111100110;
        weights1[10501] <= 16'b1111111111010101;
        weights1[10502] <= 16'b1111111111001010;
        weights1[10503] <= 16'b1111111111011011;
        weights1[10504] <= 16'b1111111111100101;
        weights1[10505] <= 16'b1111111111110111;
        weights1[10506] <= 16'b1111111111110100;
        weights1[10507] <= 16'b1111111111110011;
        weights1[10508] <= 16'b1111111111111100;
        weights1[10509] <= 16'b1111111111110000;
        weights1[10510] <= 16'b1111111111101111;
        weights1[10511] <= 16'b0000000000011011;
        weights1[10512] <= 16'b0000000000010010;
        weights1[10513] <= 16'b0000000000001100;
        weights1[10514] <= 16'b0000000000000011;
        weights1[10515] <= 16'b0000000000001001;
        weights1[10516] <= 16'b1111111111111100;
        weights1[10517] <= 16'b1111111111111111;
        weights1[10518] <= 16'b1111111111111001;
        weights1[10519] <= 16'b0000000000000110;
        weights1[10520] <= 16'b1111111111011001;
        weights1[10521] <= 16'b1111111111100110;
        weights1[10522] <= 16'b0000000000000000;
        weights1[10523] <= 16'b1111111111110101;
        weights1[10524] <= 16'b0000000000000100;
        weights1[10525] <= 16'b0000000000000110;
        weights1[10526] <= 16'b1111111111111110;
        weights1[10527] <= 16'b0000000000000111;
        weights1[10528] <= 16'b1111111111011110;
        weights1[10529] <= 16'b1111111111000111;
        weights1[10530] <= 16'b1111111110101001;
        weights1[10531] <= 16'b1111111110110101;
        weights1[10532] <= 16'b1111111110111001;
        weights1[10533] <= 16'b1111111111100111;
        weights1[10534] <= 16'b1111111111011111;
        weights1[10535] <= 16'b0000000000011110;
        weights1[10536] <= 16'b1111111111110010;
        weights1[10537] <= 16'b0000000000010000;
        weights1[10538] <= 16'b0000000000011001;
        weights1[10539] <= 16'b0000000000001101;
        weights1[10540] <= 16'b0000000000000001;
        weights1[10541] <= 16'b0000000000010101;
        weights1[10542] <= 16'b0000000000010101;
        weights1[10543] <= 16'b0000000000010101;
        weights1[10544] <= 16'b0000000000001111;
        weights1[10545] <= 16'b0000000000000101;
        weights1[10546] <= 16'b1111111111111001;
        weights1[10547] <= 16'b0000000000000001;
        weights1[10548] <= 16'b0000000000001000;
        weights1[10549] <= 16'b1111111111110101;
        weights1[10550] <= 16'b1111111111100111;
        weights1[10551] <= 16'b1111111111101010;
        weights1[10552] <= 16'b0000000000001001;
        weights1[10553] <= 16'b1111111111111101;
        weights1[10554] <= 16'b0000000000000111;
        weights1[10555] <= 16'b0000000000000110;
        weights1[10556] <= 16'b1111111111011111;
        weights1[10557] <= 16'b1111111111001001;
        weights1[10558] <= 16'b1111111110100010;
        weights1[10559] <= 16'b1111111110011101;
        weights1[10560] <= 16'b1111111101111101;
        weights1[10561] <= 16'b1111111110000111;
        weights1[10562] <= 16'b1111111110100110;
        weights1[10563] <= 16'b1111111111110001;
        weights1[10564] <= 16'b0000000000010101;
        weights1[10565] <= 16'b0000000000011011;
        weights1[10566] <= 16'b0000000000001010;
        weights1[10567] <= 16'b0000000000010100;
        weights1[10568] <= 16'b0000000000000011;
        weights1[10569] <= 16'b0000000000011101;
        weights1[10570] <= 16'b0000000000011001;
        weights1[10571] <= 16'b0000000000001011;
        weights1[10572] <= 16'b0000000000001101;
        weights1[10573] <= 16'b0000000000000010;
        weights1[10574] <= 16'b0000000000000111;
        weights1[10575] <= 16'b0000000000000000;
        weights1[10576] <= 16'b1111111111110101;
        weights1[10577] <= 16'b0000000000001000;
        weights1[10578] <= 16'b1111111111110100;
        weights1[10579] <= 16'b1111111111101111;
        weights1[10580] <= 16'b1111111111100110;
        weights1[10581] <= 16'b1111111111110111;
        weights1[10582] <= 16'b0000000000010001;
        weights1[10583] <= 16'b0000000000010111;
        weights1[10584] <= 16'b1111111111101110;
        weights1[10585] <= 16'b1111111111011010;
        weights1[10586] <= 16'b1111111110101100;
        weights1[10587] <= 16'b1111111110011011;
        weights1[10588] <= 16'b1111111101100011;
        weights1[10589] <= 16'b1111111101000110;
        weights1[10590] <= 16'b1111111100101010;
        weights1[10591] <= 16'b1111111101011011;
        weights1[10592] <= 16'b1111111110100010;
        weights1[10593] <= 16'b1111111111110100;
        weights1[10594] <= 16'b0000000000001001;
        weights1[10595] <= 16'b0000000000010110;
        weights1[10596] <= 16'b0000000000101111;
        weights1[10597] <= 16'b0000000000100001;
        weights1[10598] <= 16'b0000000000010111;
        weights1[10599] <= 16'b0000000000000011;
        weights1[10600] <= 16'b0000000000010110;
        weights1[10601] <= 16'b1111111111110111;
        weights1[10602] <= 16'b0000000000000011;
        weights1[10603] <= 16'b1111111111111111;
        weights1[10604] <= 16'b1111111111110001;
        weights1[10605] <= 16'b1111111111111100;
        weights1[10606] <= 16'b0000000000000010;
        weights1[10607] <= 16'b1111111111111011;
        weights1[10608] <= 16'b1111111111100110;
        weights1[10609] <= 16'b1111111111111011;
        weights1[10610] <= 16'b1111111111111101;
        weights1[10611] <= 16'b0000000000001010;
        weights1[10612] <= 16'b0000000000000101;
        weights1[10613] <= 16'b1111111111110111;
        weights1[10614] <= 16'b1111111111011101;
        weights1[10615] <= 16'b1111111111010100;
        weights1[10616] <= 16'b1111111111001010;
        weights1[10617] <= 16'b1111111110001010;
        weights1[10618] <= 16'b1111111100111110;
        weights1[10619] <= 16'b1111111011110000;
        weights1[10620] <= 16'b1111111011101000;
        weights1[10621] <= 16'b1111111101000100;
        weights1[10622] <= 16'b1111111110111010;
        weights1[10623] <= 16'b1111111111111100;
        weights1[10624] <= 16'b0000000000100010;
        weights1[10625] <= 16'b0000000000011100;
        weights1[10626] <= 16'b0000000000011010;
        weights1[10627] <= 16'b0000000000011011;
        weights1[10628] <= 16'b0000000000000111;
        weights1[10629] <= 16'b0000000000000100;
        weights1[10630] <= 16'b1111111111110111;
        weights1[10631] <= 16'b0000000000000111;
        weights1[10632] <= 16'b1111111111111111;
        weights1[10633] <= 16'b0000000000000101;
        weights1[10634] <= 16'b0000000000000000;
        weights1[10635] <= 16'b0000000000001010;
        weights1[10636] <= 16'b1111111111110000;
        weights1[10637] <= 16'b1111111111111010;
        weights1[10638] <= 16'b1111111111101001;
        weights1[10639] <= 16'b0000000000000001;
        weights1[10640] <= 16'b0000000000010110;
        weights1[10641] <= 16'b0000000000010100;
        weights1[10642] <= 16'b0000000000010010;
        weights1[10643] <= 16'b0000000000101110;
        weights1[10644] <= 16'b0000000000001011;
        weights1[10645] <= 16'b0000000000001100;
        weights1[10646] <= 16'b1111111111110000;
        weights1[10647] <= 16'b1111111110100000;
        weights1[10648] <= 16'b1111111100011011;
        weights1[10649] <= 16'b1111111010110000;
        weights1[10650] <= 16'b1111111011010000;
        weights1[10651] <= 16'b1111111100100010;
        weights1[10652] <= 16'b1111111101111110;
        weights1[10653] <= 16'b1111111111010111;
        weights1[10654] <= 16'b1111111111111000;
        weights1[10655] <= 16'b1111111111111011;
        weights1[10656] <= 16'b1111111111111110;
        weights1[10657] <= 16'b1111111111111001;
        weights1[10658] <= 16'b0000000000000100;
        weights1[10659] <= 16'b0000000000010000;
        weights1[10660] <= 16'b1111111111111001;
        weights1[10661] <= 16'b0000000000001010;
        weights1[10662] <= 16'b0000000000000010;
        weights1[10663] <= 16'b0000000000000010;
        weights1[10664] <= 16'b1111111111111000;
        weights1[10665] <= 16'b1111111111110100;
        weights1[10666] <= 16'b1111111111110101;
        weights1[10667] <= 16'b1111111111111001;
        weights1[10668] <= 16'b0000000000011100;
        weights1[10669] <= 16'b0000000000011001;
        weights1[10670] <= 16'b0000000000100110;
        weights1[10671] <= 16'b0000000000110001;
        weights1[10672] <= 16'b0000000000010111;
        weights1[10673] <= 16'b0000000000101110;
        weights1[10674] <= 16'b0000000000110000;
        weights1[10675] <= 16'b0000000000101101;
        weights1[10676] <= 16'b0000000000011111;
        weights1[10677] <= 16'b1111111110111011;
        weights1[10678] <= 16'b1111111101100011;
        weights1[10679] <= 16'b1111111101000111;
        weights1[10680] <= 16'b1111111100110100;
        weights1[10681] <= 16'b1111111101110001;
        weights1[10682] <= 16'b1111111110011111;
        weights1[10683] <= 16'b1111111111010010;
        weights1[10684] <= 16'b1111111111100000;
        weights1[10685] <= 16'b1111111111100101;
        weights1[10686] <= 16'b1111111111110010;
        weights1[10687] <= 16'b1111111111110001;
        weights1[10688] <= 16'b1111111111111011;
        weights1[10689] <= 16'b1111111111111001;
        weights1[10690] <= 16'b1111111111110101;
        weights1[10691] <= 16'b0000000000000011;
        weights1[10692] <= 16'b0000000000001000;
        weights1[10693] <= 16'b0000000000001000;
        weights1[10694] <= 16'b1111111111111101;
        weights1[10695] <= 16'b1111111111111011;
        weights1[10696] <= 16'b0000000000011010;
        weights1[10697] <= 16'b1111111111111011;
        weights1[10698] <= 16'b0000000000100010;
        weights1[10699] <= 16'b0000000000100010;
        weights1[10700] <= 16'b0000000000101001;
        weights1[10701] <= 16'b0000000001011011;
        weights1[10702] <= 16'b0000000001101010;
        weights1[10703] <= 16'b0000000001001111;
        weights1[10704] <= 16'b0000000001100100;
        weights1[10705] <= 16'b0000000000111000;
        weights1[10706] <= 16'b0000000000000100;
        weights1[10707] <= 16'b1111111111010011;
        weights1[10708] <= 16'b1111111110101001;
        weights1[10709] <= 16'b1111111111000110;
        weights1[10710] <= 16'b1111111111000110;
        weights1[10711] <= 16'b1111111111011010;
        weights1[10712] <= 16'b1111111111100010;
        weights1[10713] <= 16'b1111111111101100;
        weights1[10714] <= 16'b1111111111110011;
        weights1[10715] <= 16'b1111111111111101;
        weights1[10716] <= 16'b1111111111110011;
        weights1[10717] <= 16'b0000000000001100;
        weights1[10718] <= 16'b0000000000010001;
        weights1[10719] <= 16'b1111111111111110;
        weights1[10720] <= 16'b1111111111101101;
        weights1[10721] <= 16'b0000000000001111;
        weights1[10722] <= 16'b0000000000000101;
        weights1[10723] <= 16'b0000000000000000;
        weights1[10724] <= 16'b1111111111111010;
        weights1[10725] <= 16'b1111111111111101;
        weights1[10726] <= 16'b0000000000001111;
        weights1[10727] <= 16'b0000000000100000;
        weights1[10728] <= 16'b0000000000110100;
        weights1[10729] <= 16'b0000000000111011;
        weights1[10730] <= 16'b0000000001000010;
        weights1[10731] <= 16'b0000000001001010;
        weights1[10732] <= 16'b0000000001010110;
        weights1[10733] <= 16'b0000000001101011;
        weights1[10734] <= 16'b0000000001000111;
        weights1[10735] <= 16'b0000000000101011;
        weights1[10736] <= 16'b0000000000010000;
        weights1[10737] <= 16'b1111111111110001;
        weights1[10738] <= 16'b1111111111100011;
        weights1[10739] <= 16'b1111111111110000;
        weights1[10740] <= 16'b1111111111100110;
        weights1[10741] <= 16'b1111111111011111;
        weights1[10742] <= 16'b0000000000000100;
        weights1[10743] <= 16'b1111111111100011;
        weights1[10744] <= 16'b1111111111111110;
        weights1[10745] <= 16'b0000000000000000;
        weights1[10746] <= 16'b0000000000000111;
        weights1[10747] <= 16'b1111111111111000;
        weights1[10748] <= 16'b0000000000000010;
        weights1[10749] <= 16'b1111111111111100;
        weights1[10750] <= 16'b0000000000000000;
        weights1[10751] <= 16'b1111111111110111;
        weights1[10752] <= 16'b1111111111110011;
        weights1[10753] <= 16'b1111111111011110;
        weights1[10754] <= 16'b1111111111111111;
        weights1[10755] <= 16'b1111111111111001;
        weights1[10756] <= 16'b0000000000100111;
        weights1[10757] <= 16'b0000000000001100;
        weights1[10758] <= 16'b0000000000010010;
        weights1[10759] <= 16'b0000000000001101;
        weights1[10760] <= 16'b0000000000001110;
        weights1[10761] <= 16'b0000000000010000;
        weights1[10762] <= 16'b0000000000100010;
        weights1[10763] <= 16'b0000000000011100;
        weights1[10764] <= 16'b0000000000101011;
        weights1[10765] <= 16'b1111111111111011;
        weights1[10766] <= 16'b1111111111110111;
        weights1[10767] <= 16'b1111111111111100;
        weights1[10768] <= 16'b1111111111111101;
        weights1[10769] <= 16'b0000000000000100;
        weights1[10770] <= 16'b1111111111101100;
        weights1[10771] <= 16'b0000000000001001;
        weights1[10772] <= 16'b1111111111110010;
        weights1[10773] <= 16'b0000000000000111;
        weights1[10774] <= 16'b1111111111101110;
        weights1[10775] <= 16'b0000000000000000;
        weights1[10776] <= 16'b0000000000000100;
        weights1[10777] <= 16'b1111111111111100;
        weights1[10778] <= 16'b1111111111111100;
        weights1[10779] <= 16'b1111111111111110;
        weights1[10780] <= 16'b1111111111101101;
        weights1[10781] <= 16'b1111111111010111;
        weights1[10782] <= 16'b1111111111000111;
        weights1[10783] <= 16'b1111111111010110;
        weights1[10784] <= 16'b1111111111111101;
        weights1[10785] <= 16'b0000000000001110;
        weights1[10786] <= 16'b0000000000001010;
        weights1[10787] <= 16'b0000000000001011;
        weights1[10788] <= 16'b0000000000010100;
        weights1[10789] <= 16'b1111111111111000;
        weights1[10790] <= 16'b0000000000010010;
        weights1[10791] <= 16'b0000000000011010;
        weights1[10792] <= 16'b0000000000010110;
        weights1[10793] <= 16'b0000000000011100;
        weights1[10794] <= 16'b0000000000100010;
        weights1[10795] <= 16'b0000000000001110;
        weights1[10796] <= 16'b1111111111111011;
        weights1[10797] <= 16'b0000000000000011;
        weights1[10798] <= 16'b1111111111111000;
        weights1[10799] <= 16'b0000000000000011;
        weights1[10800] <= 16'b0000000000000000;
        weights1[10801] <= 16'b1111111111110100;
        weights1[10802] <= 16'b0000000000001011;
        weights1[10803] <= 16'b1111111111110111;
        weights1[10804] <= 16'b1111111111110100;
        weights1[10805] <= 16'b1111111111111001;
        weights1[10806] <= 16'b1111111111101110;
        weights1[10807] <= 16'b1111111111110010;
        weights1[10808] <= 16'b1111111111101100;
        weights1[10809] <= 16'b1111111111011000;
        weights1[10810] <= 16'b1111111111000011;
        weights1[10811] <= 16'b1111111110111011;
        weights1[10812] <= 16'b1111111111000111;
        weights1[10813] <= 16'b1111111111000110;
        weights1[10814] <= 16'b1111111111110100;
        weights1[10815] <= 16'b1111111111101110;
        weights1[10816] <= 16'b0000000000000000;
        weights1[10817] <= 16'b0000000000011010;
        weights1[10818] <= 16'b0000000000000111;
        weights1[10819] <= 16'b0000000000000110;
        weights1[10820] <= 16'b0000000000000100;
        weights1[10821] <= 16'b0000000000001010;
        weights1[10822] <= 16'b0000000000000000;
        weights1[10823] <= 16'b0000000000001001;
        weights1[10824] <= 16'b0000000000001010;
        weights1[10825] <= 16'b1111111111111001;
        weights1[10826] <= 16'b0000000000001110;
        weights1[10827] <= 16'b1111111111111000;
        weights1[10828] <= 16'b1111111111110111;
        weights1[10829] <= 16'b1111111111110111;
        weights1[10830] <= 16'b1111111111101110;
        weights1[10831] <= 16'b0000000000001101;
        weights1[10832] <= 16'b1111111111110110;
        weights1[10833] <= 16'b1111111111111111;
        weights1[10834] <= 16'b1111111111101111;
        weights1[10835] <= 16'b1111111111111000;
        weights1[10836] <= 16'b1111111111110110;
        weights1[10837] <= 16'b1111111111100110;
        weights1[10838] <= 16'b1111111111011001;
        weights1[10839] <= 16'b1111111111001111;
        weights1[10840] <= 16'b1111111111001011;
        weights1[10841] <= 16'b1111111111100101;
        weights1[10842] <= 16'b1111111111101110;
        weights1[10843] <= 16'b1111111111111011;
        weights1[10844] <= 16'b1111111111111001;
        weights1[10845] <= 16'b1111111111111100;
        weights1[10846] <= 16'b0000000000110110;
        weights1[10847] <= 16'b0000000000011000;
        weights1[10848] <= 16'b0000000000001100;
        weights1[10849] <= 16'b0000000000001111;
        weights1[10850] <= 16'b0000000000001111;
        weights1[10851] <= 16'b0000000000000111;
        weights1[10852] <= 16'b1111111111110111;
        weights1[10853] <= 16'b0000000000000011;
        weights1[10854] <= 16'b0000000000001111;
        weights1[10855] <= 16'b0000000000000111;
        weights1[10856] <= 16'b0000000000010000;
        weights1[10857] <= 16'b0000000000000110;
        weights1[10858] <= 16'b1111111111111001;
        weights1[10859] <= 16'b1111111111101101;
        weights1[10860] <= 16'b1111111111110110;
        weights1[10861] <= 16'b1111111111110110;
        weights1[10862] <= 16'b1111111111110100;
        weights1[10863] <= 16'b1111111111110110;
        weights1[10864] <= 16'b1111111111111010;
        weights1[10865] <= 16'b1111111111110011;
        weights1[10866] <= 16'b1111111111101101;
        weights1[10867] <= 16'b1111111111011011;
        weights1[10868] <= 16'b1111111111011110;
        weights1[10869] <= 16'b1111111111010110;
        weights1[10870] <= 16'b1111111111011010;
        weights1[10871] <= 16'b1111111111111100;
        weights1[10872] <= 16'b0000000000000000;
        weights1[10873] <= 16'b1111111111111110;
        weights1[10874] <= 16'b0000000000000001;
        weights1[10875] <= 16'b1111111111111110;
        weights1[10876] <= 16'b0000000000010000;
        weights1[10877] <= 16'b1111111111111000;
        weights1[10878] <= 16'b0000000000000101;
        weights1[10879] <= 16'b0000000000000101;
        weights1[10880] <= 16'b1111111111110101;
        weights1[10881] <= 16'b0000000000000010;
        weights1[10882] <= 16'b0000000000000011;
        weights1[10883] <= 16'b1111111111101100;
        weights1[10884] <= 16'b1111111111110011;
        weights1[10885] <= 16'b0000000000000110;
        weights1[10886] <= 16'b1111111111011111;
        weights1[10887] <= 16'b1111111111101001;
        weights1[10888] <= 16'b1111111111110001;
        weights1[10889] <= 16'b1111111111110011;
        weights1[10890] <= 16'b1111111111111001;
        weights1[10891] <= 16'b1111111111111101;
        weights1[10892] <= 16'b1111111111111111;
        weights1[10893] <= 16'b1111111111111101;
        weights1[10894] <= 16'b1111111111111000;
        weights1[10895] <= 16'b1111111111111011;
        weights1[10896] <= 16'b1111111111101101;
        weights1[10897] <= 16'b1111111111011111;
        weights1[10898] <= 16'b1111111111100110;
        weights1[10899] <= 16'b1111111111110111;
        weights1[10900] <= 16'b1111111111111011;
        weights1[10901] <= 16'b1111111111100000;
        weights1[10902] <= 16'b1111111111111111;
        weights1[10903] <= 16'b1111111111101010;
        weights1[10904] <= 16'b1111111111110011;
        weights1[10905] <= 16'b0000000000001101;
        weights1[10906] <= 16'b0000000000010100;
        weights1[10907] <= 16'b0000000000000110;
        weights1[10908] <= 16'b0000000000000110;
        weights1[10909] <= 16'b0000000000001110;
        weights1[10910] <= 16'b0000000000000010;
        weights1[10911] <= 16'b1111111111111001;
        weights1[10912] <= 16'b1111111111110110;
        weights1[10913] <= 16'b1111111111101000;
        weights1[10914] <= 16'b1111111111011011;
        weights1[10915] <= 16'b1111111111101011;
        weights1[10916] <= 16'b1111111111110101;
        weights1[10917] <= 16'b1111111111110101;
        weights1[10918] <= 16'b1111111111111010;
        weights1[10919] <= 16'b0000000000000000;
        weights1[10920] <= 16'b1111111111111110;
        weights1[10921] <= 16'b1111111111111100;
        weights1[10922] <= 16'b0000000000000001;
        weights1[10923] <= 16'b0000000000000000;
        weights1[10924] <= 16'b1111111111111010;
        weights1[10925] <= 16'b1111111111110111;
        weights1[10926] <= 16'b1111111111101011;
        weights1[10927] <= 16'b1111111111011001;
        weights1[10928] <= 16'b1111111111100011;
        weights1[10929] <= 16'b1111111111100110;
        weights1[10930] <= 16'b1111111111110100;
        weights1[10931] <= 16'b1111111111100110;
        weights1[10932] <= 16'b1111111111111000;
        weights1[10933] <= 16'b1111111111111000;
        weights1[10934] <= 16'b1111111111100111;
        weights1[10935] <= 16'b1111111111110110;
        weights1[10936] <= 16'b0000000000000010;
        weights1[10937] <= 16'b1111111111111110;
        weights1[10938] <= 16'b1111111111101111;
        weights1[10939] <= 16'b1111111111101100;
        weights1[10940] <= 16'b1111111111101111;
        weights1[10941] <= 16'b1111111111100000;
        weights1[10942] <= 16'b1111111111101001;
        weights1[10943] <= 16'b1111111111111000;
        weights1[10944] <= 16'b1111111111111000;
        weights1[10945] <= 16'b1111111111111001;
        weights1[10946] <= 16'b1111111111111110;
        weights1[10947] <= 16'b0000000000000000;
        weights1[10948] <= 16'b0000000000000001;
        weights1[10949] <= 16'b0000000000000000;
        weights1[10950] <= 16'b0000000000000010;
        weights1[10951] <= 16'b0000000000001001;
        weights1[10952] <= 16'b0000000000000110;
        weights1[10953] <= 16'b0000000000000100;
        weights1[10954] <= 16'b0000000000000110;
        weights1[10955] <= 16'b1111111111111010;
        weights1[10956] <= 16'b1111111111100111;
        weights1[10957] <= 16'b1111111111101001;
        weights1[10958] <= 16'b1111111111011011;
        weights1[10959] <= 16'b1111111111011000;
        weights1[10960] <= 16'b1111111111100111;
        weights1[10961] <= 16'b1111111111100000;
        weights1[10962] <= 16'b1111111111101001;
        weights1[10963] <= 16'b1111111111101110;
        weights1[10964] <= 16'b1111111111100111;
        weights1[10965] <= 16'b1111111111100001;
        weights1[10966] <= 16'b1111111111110010;
        weights1[10967] <= 16'b1111111111110110;
        weights1[10968] <= 16'b1111111111110011;
        weights1[10969] <= 16'b1111111111101110;
        weights1[10970] <= 16'b1111111111110010;
        weights1[10971] <= 16'b1111111111110110;
        weights1[10972] <= 16'b1111111111111011;
        weights1[10973] <= 16'b1111111111111100;
        weights1[10974] <= 16'b0000000000000000;
        weights1[10975] <= 16'b0000000000000000;
        weights1[10976] <= 16'b0000000000000000;
        weights1[10977] <= 16'b0000000000000000;
        weights1[10978] <= 16'b0000000000000000;
        weights1[10979] <= 16'b0000000000000000;
        weights1[10980] <= 16'b1111111111111011;
        weights1[10981] <= 16'b1111111111111001;
        weights1[10982] <= 16'b1111111111111010;
        weights1[10983] <= 16'b1111111111111010;
        weights1[10984] <= 16'b1111111111110011;
        weights1[10985] <= 16'b1111111111101010;
        weights1[10986] <= 16'b1111111111110001;
        weights1[10987] <= 16'b1111111111110100;
        weights1[10988] <= 16'b1111111111110110;
        weights1[10989] <= 16'b1111111111111101;
        weights1[10990] <= 16'b1111111111110010;
        weights1[10991] <= 16'b1111111111111011;
        weights1[10992] <= 16'b0000000000001111;
        weights1[10993] <= 16'b0000000000000011;
        weights1[10994] <= 16'b1111111111111111;
        weights1[10995] <= 16'b1111111111111001;
        weights1[10996] <= 16'b1111111111110010;
        weights1[10997] <= 16'b1111111111111110;
        weights1[10998] <= 16'b0000000000000011;
        weights1[10999] <= 16'b0000000000000001;
        weights1[11000] <= 16'b1111111111111101;
        weights1[11001] <= 16'b1111111111111101;
        weights1[11002] <= 16'b1111111111111100;
        weights1[11003] <= 16'b1111111111111101;
        weights1[11004] <= 16'b0000000000000000;
        weights1[11005] <= 16'b0000000000000000;
        weights1[11006] <= 16'b1111111111111011;
        weights1[11007] <= 16'b1111111111111000;
        weights1[11008] <= 16'b1111111111111111;
        weights1[11009] <= 16'b1111111111110110;
        weights1[11010] <= 16'b1111111111110110;
        weights1[11011] <= 16'b1111111111110110;
        weights1[11012] <= 16'b1111111111111111;
        weights1[11013] <= 16'b1111111111101110;
        weights1[11014] <= 16'b1111111111110101;
        weights1[11015] <= 16'b1111111111110001;
        weights1[11016] <= 16'b1111111111110101;
        weights1[11017] <= 16'b1111111111111000;
        weights1[11018] <= 16'b0000000000000000;
        weights1[11019] <= 16'b1111111111111110;
        weights1[11020] <= 16'b1111111111111111;
        weights1[11021] <= 16'b1111111111110011;
        weights1[11022] <= 16'b0000000000000101;
        weights1[11023] <= 16'b1111111111111010;
        weights1[11024] <= 16'b1111111111111101;
        weights1[11025] <= 16'b1111111111111010;
        weights1[11026] <= 16'b0000000000000101;
        weights1[11027] <= 16'b1111111111110111;
        weights1[11028] <= 16'b1111111111110110;
        weights1[11029] <= 16'b1111111111111110;
        weights1[11030] <= 16'b1111111111111110;
        weights1[11031] <= 16'b1111111111111111;
        weights1[11032] <= 16'b1111111111111110;
        weights1[11033] <= 16'b1111111111111101;
        weights1[11034] <= 16'b1111111111110111;
        weights1[11035] <= 16'b1111111111111010;
        weights1[11036] <= 16'b1111111111110011;
        weights1[11037] <= 16'b1111111111111010;
        weights1[11038] <= 16'b1111111111111010;
        weights1[11039] <= 16'b1111111111111001;
        weights1[11040] <= 16'b1111111111111111;
        weights1[11041] <= 16'b0000000000000001;
        weights1[11042] <= 16'b1111111111110111;
        weights1[11043] <= 16'b1111111111111101;
        weights1[11044] <= 16'b1111111111111010;
        weights1[11045] <= 16'b0000000000000011;
        weights1[11046] <= 16'b1111111111111101;
        weights1[11047] <= 16'b0000000000001001;
        weights1[11048] <= 16'b1111111111111001;
        weights1[11049] <= 16'b1111111111111010;
        weights1[11050] <= 16'b1111111111110010;
        weights1[11051] <= 16'b1111111111111101;
        weights1[11052] <= 16'b0000000000000111;
        weights1[11053] <= 16'b1111111111111100;
        weights1[11054] <= 16'b1111111111110110;
        weights1[11055] <= 16'b0000000000000011;
        weights1[11056] <= 16'b1111111111111001;
        weights1[11057] <= 16'b0000000000001000;
        weights1[11058] <= 16'b1111111111111111;
        weights1[11059] <= 16'b1111111111111100;
        weights1[11060] <= 16'b1111111111111111;
        weights1[11061] <= 16'b1111111111111101;
        weights1[11062] <= 16'b0000000000000001;
        weights1[11063] <= 16'b0000000000000101;
        weights1[11064] <= 16'b1111111111111001;
        weights1[11065] <= 16'b1111111111111111;
        weights1[11066] <= 16'b0000000000001111;
        weights1[11067] <= 16'b1111111111111111;
        weights1[11068] <= 16'b1111111111111111;
        weights1[11069] <= 16'b0000000000000001;
        weights1[11070] <= 16'b1111111111111011;
        weights1[11071] <= 16'b1111111111111110;
        weights1[11072] <= 16'b1111111111110010;
        weights1[11073] <= 16'b1111111111110110;
        weights1[11074] <= 16'b1111111111110100;
        weights1[11075] <= 16'b0000000000000000;
        weights1[11076] <= 16'b1111111111101011;
        weights1[11077] <= 16'b0000000000010010;
        weights1[11078] <= 16'b0000000000010100;
        weights1[11079] <= 16'b0000000000000100;
        weights1[11080] <= 16'b1111111111111001;
        weights1[11081] <= 16'b1111111111101100;
        weights1[11082] <= 16'b1111111111111000;
        weights1[11083] <= 16'b1111111111101111;
        weights1[11084] <= 16'b1111111111111101;
        weights1[11085] <= 16'b1111111111110101;
        weights1[11086] <= 16'b0000000000000000;
        weights1[11087] <= 16'b0000000000000100;
        weights1[11088] <= 16'b1111111111111110;
        weights1[11089] <= 16'b1111111111111100;
        weights1[11090] <= 16'b1111111111111100;
        weights1[11091] <= 16'b0000000000000011;
        weights1[11092] <= 16'b1111111111111001;
        weights1[11093] <= 16'b0000000000001011;
        weights1[11094] <= 16'b0000000000000000;
        weights1[11095] <= 16'b1111111111110100;
        weights1[11096] <= 16'b1111111111111110;
        weights1[11097] <= 16'b1111111111111011;
        weights1[11098] <= 16'b1111111111111001;
        weights1[11099] <= 16'b1111111111111110;
        weights1[11100] <= 16'b0000000000000011;
        weights1[11101] <= 16'b0000000000001100;
        weights1[11102] <= 16'b1111111111110101;
        weights1[11103] <= 16'b0000000000001110;
        weights1[11104] <= 16'b0000000000010010;
        weights1[11105] <= 16'b1111111111101011;
        weights1[11106] <= 16'b1111111111110110;
        weights1[11107] <= 16'b0000000000000010;
        weights1[11108] <= 16'b0000000000000101;
        weights1[11109] <= 16'b0000000000001011;
        weights1[11110] <= 16'b0000000000000000;
        weights1[11111] <= 16'b1111111111111011;
        weights1[11112] <= 16'b0000000000001011;
        weights1[11113] <= 16'b1111111111111100;
        weights1[11114] <= 16'b1111111111111101;
        weights1[11115] <= 16'b0000000000000110;
        weights1[11116] <= 16'b0000000000000100;
        weights1[11117] <= 16'b1111111111111011;
        weights1[11118] <= 16'b0000000000000010;
        weights1[11119] <= 16'b1111111111111010;
        weights1[11120] <= 16'b1111111111111100;
        weights1[11121] <= 16'b0000000000001000;
        weights1[11122] <= 16'b0000000000000010;
        weights1[11123] <= 16'b1111111111111110;
        weights1[11124] <= 16'b0000000000001010;
        weights1[11125] <= 16'b0000000000000001;
        weights1[11126] <= 16'b1111111111111001;
        weights1[11127] <= 16'b1111111111111001;
        weights1[11128] <= 16'b0000000000001001;
        weights1[11129] <= 16'b0000000000000110;
        weights1[11130] <= 16'b1111111111110111;
        weights1[11131] <= 16'b1111111111110101;
        weights1[11132] <= 16'b0000000000000100;
        weights1[11133] <= 16'b1111111111111001;
        weights1[11134] <= 16'b0000000000001011;
        weights1[11135] <= 16'b1111111111111011;
        weights1[11136] <= 16'b1111111111111110;
        weights1[11137] <= 16'b1111111111111101;
        weights1[11138] <= 16'b1111111111110101;
        weights1[11139] <= 16'b1111111111111010;
        weights1[11140] <= 16'b0000000000000111;
        weights1[11141] <= 16'b0000000000000101;
        weights1[11142] <= 16'b0000000000000010;
        weights1[11143] <= 16'b0000000000000010;
        weights1[11144] <= 16'b0000000000000101;
        weights1[11145] <= 16'b1111111111111101;
        weights1[11146] <= 16'b1111111111110110;
        weights1[11147] <= 16'b0000000000001001;
        weights1[11148] <= 16'b1111111111111111;
        weights1[11149] <= 16'b1111111111101110;
        weights1[11150] <= 16'b0000000000000011;
        weights1[11151] <= 16'b0000000000000001;
        weights1[11152] <= 16'b1111111111111001;
        weights1[11153] <= 16'b0000000000001111;
        weights1[11154] <= 16'b1111111111110110;
        weights1[11155] <= 16'b1111111111111110;
        weights1[11156] <= 16'b1111111111110010;
        weights1[11157] <= 16'b1111111111101101;
        weights1[11158] <= 16'b0000000000000000;
        weights1[11159] <= 16'b0000000000000101;
        weights1[11160] <= 16'b1111111111111011;
        weights1[11161] <= 16'b0000000000000001;
        weights1[11162] <= 16'b0000000000010000;
        weights1[11163] <= 16'b1111111111110011;
        weights1[11164] <= 16'b0000000000000100;
        weights1[11165] <= 16'b1111111111110100;
        weights1[11166] <= 16'b1111111111111100;
        weights1[11167] <= 16'b0000000000001101;
        weights1[11168] <= 16'b0000000000000001;
        weights1[11169] <= 16'b1111111111111111;
        weights1[11170] <= 16'b0000000000000100;
        weights1[11171] <= 16'b0000000000001000;
        weights1[11172] <= 16'b0000000000000000;
        weights1[11173] <= 16'b1111111111111100;
        weights1[11174] <= 16'b0000000000000001;
        weights1[11175] <= 16'b1111111111110111;
        weights1[11176] <= 16'b0000000000000100;
        weights1[11177] <= 16'b1111111111111011;
        weights1[11178] <= 16'b0000000000001011;
        weights1[11179] <= 16'b0000000000001001;
        weights1[11180] <= 16'b1111111111111000;
        weights1[11181] <= 16'b1111111111110111;
        weights1[11182] <= 16'b0000000000000011;
        weights1[11183] <= 16'b1111111111110111;
        weights1[11184] <= 16'b1111111111111001;
        weights1[11185] <= 16'b1111111111111010;
        weights1[11186] <= 16'b0000000000000011;
        weights1[11187] <= 16'b1111111111110010;
        weights1[11188] <= 16'b1111111111111100;
        weights1[11189] <= 16'b1111111111111111;
        weights1[11190] <= 16'b0000000000000001;
        weights1[11191] <= 16'b1111111111101100;
        weights1[11192] <= 16'b0000000000001111;
        weights1[11193] <= 16'b1111111111101111;
        weights1[11194] <= 16'b0000000000001110;
        weights1[11195] <= 16'b0000000000001011;
        weights1[11196] <= 16'b1111111111110111;
        weights1[11197] <= 16'b0000000000001010;
        weights1[11198] <= 16'b0000000000000111;
        weights1[11199] <= 16'b1111111111111110;
        weights1[11200] <= 16'b0000000000001000;
        weights1[11201] <= 16'b0000000000000110;
        weights1[11202] <= 16'b0000000000001011;
        weights1[11203] <= 16'b0000000000001000;
        weights1[11204] <= 16'b1111111111110110;
        weights1[11205] <= 16'b0000000000010000;
        weights1[11206] <= 16'b0000000000000110;
        weights1[11207] <= 16'b0000000000000111;
        weights1[11208] <= 16'b1111111111110101;
        weights1[11209] <= 16'b1111111111111010;
        weights1[11210] <= 16'b1111111111110111;
        weights1[11211] <= 16'b0000000000000001;
        weights1[11212] <= 16'b0000000000001001;
        weights1[11213] <= 16'b0000000000001010;
        weights1[11214] <= 16'b0000000000000010;
        weights1[11215] <= 16'b0000000000001010;
        weights1[11216] <= 16'b1111111111101110;
        weights1[11217] <= 16'b0000000000001011;
        weights1[11218] <= 16'b0000000000000110;
        weights1[11219] <= 16'b1111111111111010;
        weights1[11220] <= 16'b0000000000001101;
        weights1[11221] <= 16'b0000000000000010;
        weights1[11222] <= 16'b0000000000000010;
        weights1[11223] <= 16'b0000000000000000;
        weights1[11224] <= 16'b0000000000001000;
        weights1[11225] <= 16'b1111111111111001;
        weights1[11226] <= 16'b1111111111111111;
        weights1[11227] <= 16'b1111111111101111;
        weights1[11228] <= 16'b0000000000001010;
        weights1[11229] <= 16'b0000000000000101;
        weights1[11230] <= 16'b0000000000000100;
        weights1[11231] <= 16'b1111111111111101;
        weights1[11232] <= 16'b1111111111110111;
        weights1[11233] <= 16'b0000000000000000;
        weights1[11234] <= 16'b1111111111111011;
        weights1[11235] <= 16'b0000000000001011;
        weights1[11236] <= 16'b0000000000001100;
        weights1[11237] <= 16'b0000000000011001;
        weights1[11238] <= 16'b0000000000000010;
        weights1[11239] <= 16'b1111111111101110;
        weights1[11240] <= 16'b1111111111111111;
        weights1[11241] <= 16'b0000000000000110;
        weights1[11242] <= 16'b1111111111111110;
        weights1[11243] <= 16'b0000000000000010;
        weights1[11244] <= 16'b1111111111110111;
        weights1[11245] <= 16'b1111111111111010;
        weights1[11246] <= 16'b1111111111111100;
        weights1[11247] <= 16'b1111111111110110;
        weights1[11248] <= 16'b1111111111110111;
        weights1[11249] <= 16'b1111111111101010;
        weights1[11250] <= 16'b0000000000000110;
        weights1[11251] <= 16'b1111111111111111;
        weights1[11252] <= 16'b1111111111111101;
        weights1[11253] <= 16'b0000000000001100;
        weights1[11254] <= 16'b0000000000000110;
        weights1[11255] <= 16'b1111111111111110;
        weights1[11256] <= 16'b0000000000010000;
        weights1[11257] <= 16'b0000000000000100;
        weights1[11258] <= 16'b0000000000001001;
        weights1[11259] <= 16'b0000000000000001;
        weights1[11260] <= 16'b1111111111111100;
        weights1[11261] <= 16'b0000000000000001;
        weights1[11262] <= 16'b1111111111110100;
        weights1[11263] <= 16'b1111111111111010;
        weights1[11264] <= 16'b0000000000000011;
        weights1[11265] <= 16'b0000000000000010;
        weights1[11266] <= 16'b1111111111101001;
        weights1[11267] <= 16'b0000000000000100;
        weights1[11268] <= 16'b0000000000001100;
        weights1[11269] <= 16'b1111111111111010;
        weights1[11270] <= 16'b0000000000001110;
        weights1[11271] <= 16'b0000000000000011;
        weights1[11272] <= 16'b1111111111101011;
        weights1[11273] <= 16'b0000000000001110;
        weights1[11274] <= 16'b1111111111110110;
        weights1[11275] <= 16'b1111111111111001;
        weights1[11276] <= 16'b0000000000001010;
        weights1[11277] <= 16'b0000000000001010;
        weights1[11278] <= 16'b1111111111111000;
        weights1[11279] <= 16'b0000000000000101;
        weights1[11280] <= 16'b1111111111111100;
        weights1[11281] <= 16'b1111111111111011;
        weights1[11282] <= 16'b0000000000000001;
        weights1[11283] <= 16'b0000000000000111;
        weights1[11284] <= 16'b0000000000001101;
        weights1[11285] <= 16'b0000000000001000;
        weights1[11286] <= 16'b0000000000010001;
        weights1[11287] <= 16'b0000000000001001;
        weights1[11288] <= 16'b0000000000000111;
        weights1[11289] <= 16'b0000000000001100;
        weights1[11290] <= 16'b0000000000010110;
        weights1[11291] <= 16'b1111111111110101;
        weights1[11292] <= 16'b0000000000001000;
        weights1[11293] <= 16'b0000000000001011;
        weights1[11294] <= 16'b0000000000000011;
        weights1[11295] <= 16'b0000000000000010;
        weights1[11296] <= 16'b0000000000000110;
        weights1[11297] <= 16'b1111111111101100;
        weights1[11298] <= 16'b0000000000000000;
        weights1[11299] <= 16'b0000000000001011;
        weights1[11300] <= 16'b0000000000000011;
        weights1[11301] <= 16'b0000000000000111;
        weights1[11302] <= 16'b1111111111111100;
        weights1[11303] <= 16'b1111111111111101;
        weights1[11304] <= 16'b1111111111111001;
        weights1[11305] <= 16'b0000000000000010;
        weights1[11306] <= 16'b0000000000001100;
        weights1[11307] <= 16'b0000000000000110;
        weights1[11308] <= 16'b0000000000000011;
        weights1[11309] <= 16'b1111111111111010;
        weights1[11310] <= 16'b1111111111110010;
        weights1[11311] <= 16'b0000000000000101;
        weights1[11312] <= 16'b0000000000000010;
        weights1[11313] <= 16'b0000000000000010;
        weights1[11314] <= 16'b1111111111111111;
        weights1[11315] <= 16'b0000000000001011;
        weights1[11316] <= 16'b0000000000010011;
        weights1[11317] <= 16'b1111111111111100;
        weights1[11318] <= 16'b1111111111111001;
        weights1[11319] <= 16'b0000000000001100;
        weights1[11320] <= 16'b0000000000000100;
        weights1[11321] <= 16'b0000000000000001;
        weights1[11322] <= 16'b1111111111110101;
        weights1[11323] <= 16'b0000000000000011;
        weights1[11324] <= 16'b0000000000000111;
        weights1[11325] <= 16'b1111111111111101;
        weights1[11326] <= 16'b1111111111111010;
        weights1[11327] <= 16'b1111111111111111;
        weights1[11328] <= 16'b0000000000000111;
        weights1[11329] <= 16'b1111111111101101;
        weights1[11330] <= 16'b1111111111111100;
        weights1[11331] <= 16'b0000000000000111;
        weights1[11332] <= 16'b0000000000000000;
        weights1[11333] <= 16'b0000000000000010;
        weights1[11334] <= 16'b1111111111101110;
        weights1[11335] <= 16'b1111111111110011;
        weights1[11336] <= 16'b1111111111111011;
        weights1[11337] <= 16'b1111111111111011;
        weights1[11338] <= 16'b1111111111111010;
        weights1[11339] <= 16'b1111111111111011;
        weights1[11340] <= 16'b0000000000000100;
        weights1[11341] <= 16'b1111111111110101;
        weights1[11342] <= 16'b0000000000000011;
        weights1[11343] <= 16'b0000000000000111;
        weights1[11344] <= 16'b0000000000000000;
        weights1[11345] <= 16'b1111111111111101;
        weights1[11346] <= 16'b1111111111111111;
        weights1[11347] <= 16'b0000000000001001;
        weights1[11348] <= 16'b0000000000000100;
        weights1[11349] <= 16'b0000000000001000;
        weights1[11350] <= 16'b1111111111111001;
        weights1[11351] <= 16'b0000000000010011;
        weights1[11352] <= 16'b1111111111110011;
        weights1[11353] <= 16'b1111111111111100;
        weights1[11354] <= 16'b1111111111111111;
        weights1[11355] <= 16'b0000000000000111;
        weights1[11356] <= 16'b1111111111111101;
        weights1[11357] <= 16'b0000000000000110;
        weights1[11358] <= 16'b0000000000000000;
        weights1[11359] <= 16'b1111111111110101;
        weights1[11360] <= 16'b1111111111111011;
        weights1[11361] <= 16'b0000000000010000;
        weights1[11362] <= 16'b0000000000001110;
        weights1[11363] <= 16'b1111111111110010;
        weights1[11364] <= 16'b0000000000000100;
        weights1[11365] <= 16'b0000000000000001;
        weights1[11366] <= 16'b0000000000001001;
        weights1[11367] <= 16'b1111111111110110;
        weights1[11368] <= 16'b0000000000000001;
        weights1[11369] <= 16'b0000000000000011;
        weights1[11370] <= 16'b0000000000001110;
        weights1[11371] <= 16'b1111111111110101;
        weights1[11372] <= 16'b0000000000001001;
        weights1[11373] <= 16'b0000000000000000;
        weights1[11374] <= 16'b0000000000000010;
        weights1[11375] <= 16'b1111111111111100;
        weights1[11376] <= 16'b1111111111111000;
        weights1[11377] <= 16'b1111111111111111;
        weights1[11378] <= 16'b0000000000001000;
        weights1[11379] <= 16'b1111111111111000;
        weights1[11380] <= 16'b1111111111111000;
        weights1[11381] <= 16'b1111111111110101;
        weights1[11382] <= 16'b1111111111111101;
        weights1[11383] <= 16'b1111111111110110;
        weights1[11384] <= 16'b1111111111110110;
        weights1[11385] <= 16'b0000000000001001;
        weights1[11386] <= 16'b1111111111111100;
        weights1[11387] <= 16'b0000000000000110;
        weights1[11388] <= 16'b1111111111111111;
        weights1[11389] <= 16'b1111111111111111;
        weights1[11390] <= 16'b0000000000000101;
        weights1[11391] <= 16'b0000000000000101;
        weights1[11392] <= 16'b1111111111101100;
        weights1[11393] <= 16'b0000000000010111;
        weights1[11394] <= 16'b1111111111101101;
        weights1[11395] <= 16'b1111111111110111;
        weights1[11396] <= 16'b1111111111111110;
        weights1[11397] <= 16'b0000000000000100;
        weights1[11398] <= 16'b1111111111111010;
        weights1[11399] <= 16'b1111111111111100;
        weights1[11400] <= 16'b0000000000000111;
        weights1[11401] <= 16'b1111111111111101;
        weights1[11402] <= 16'b1111111111111110;
        weights1[11403] <= 16'b1111111111111100;
        weights1[11404] <= 16'b0000000000001110;
        weights1[11405] <= 16'b0000000000001100;
        weights1[11406] <= 16'b0000000000001010;
        weights1[11407] <= 16'b1111111111111000;
        weights1[11408] <= 16'b1111111111111110;
        weights1[11409] <= 16'b0000000000000000;
        weights1[11410] <= 16'b0000000000001000;
        weights1[11411] <= 16'b0000000000000110;
        weights1[11412] <= 16'b0000000000000001;
        weights1[11413] <= 16'b0000000000000101;
        weights1[11414] <= 16'b1111111111111111;
        weights1[11415] <= 16'b0000000000000011;
        weights1[11416] <= 16'b0000000000001000;
        weights1[11417] <= 16'b0000000000000111;
        weights1[11418] <= 16'b1111111111111111;
        weights1[11419] <= 16'b0000000000000010;
        weights1[11420] <= 16'b1111111111111011;
        weights1[11421] <= 16'b0000000000000001;
        weights1[11422] <= 16'b0000000000000000;
        weights1[11423] <= 16'b1111111111111011;
        weights1[11424] <= 16'b1111111111110010;
        weights1[11425] <= 16'b1111111111110011;
        weights1[11426] <= 16'b1111111111110001;
        weights1[11427] <= 16'b1111111111101000;
        weights1[11428] <= 16'b1111111111110111;
        weights1[11429] <= 16'b1111111111101011;
        weights1[11430] <= 16'b1111111111101110;
        weights1[11431] <= 16'b0000000000001100;
        weights1[11432] <= 16'b0000000000010010;
        weights1[11433] <= 16'b0000000000000101;
        weights1[11434] <= 16'b0000000000000110;
        weights1[11435] <= 16'b1111111111110011;
        weights1[11436] <= 16'b1111111111110000;
        weights1[11437] <= 16'b1111111111111000;
        weights1[11438] <= 16'b1111111111111101;
        weights1[11439] <= 16'b0000000000000001;
        weights1[11440] <= 16'b0000000000000010;
        weights1[11441] <= 16'b1111111111111100;
        weights1[11442] <= 16'b1111111111110000;
        weights1[11443] <= 16'b0000000000000011;
        weights1[11444] <= 16'b0000000000001010;
        weights1[11445] <= 16'b0000000000001110;
        weights1[11446] <= 16'b0000000000011010;
        weights1[11447] <= 16'b0000000000010111;
        weights1[11448] <= 16'b0000000000000100;
        weights1[11449] <= 16'b1111111111110010;
        weights1[11450] <= 16'b1111111111111011;
        weights1[11451] <= 16'b1111111111111011;
        weights1[11452] <= 16'b1111111111101100;
        weights1[11453] <= 16'b1111111111101110;
        weights1[11454] <= 16'b1111111111100111;
        weights1[11455] <= 16'b1111111111101110;
        weights1[11456] <= 16'b1111111111110101;
        weights1[11457] <= 16'b1111111111101110;
        weights1[11458] <= 16'b0000000000010000;
        weights1[11459] <= 16'b0000000000010000;
        weights1[11460] <= 16'b0000000000011111;
        weights1[11461] <= 16'b0000000000000011;
        weights1[11462] <= 16'b1111111111110110;
        weights1[11463] <= 16'b1111111111100101;
        weights1[11464] <= 16'b1111111111101000;
        weights1[11465] <= 16'b1111111111111001;
        weights1[11466] <= 16'b0000000000001110;
        weights1[11467] <= 16'b0000000000000110;
        weights1[11468] <= 16'b0000000000001101;
        weights1[11469] <= 16'b1111111111110000;
        weights1[11470] <= 16'b1111111111111000;
        weights1[11471] <= 16'b1111111111111000;
        weights1[11472] <= 16'b1111111111111101;
        weights1[11473] <= 16'b1111111111111111;
        weights1[11474] <= 16'b0000000000100110;
        weights1[11475] <= 16'b0000000000010111;
        weights1[11476] <= 16'b0000000000010010;
        weights1[11477] <= 16'b0000000000000011;
        weights1[11478] <= 16'b1111111111111010;
        weights1[11479] <= 16'b1111111111111011;
        weights1[11480] <= 16'b1111111111101000;
        weights1[11481] <= 16'b1111111111011101;
        weights1[11482] <= 16'b1111111111010100;
        weights1[11483] <= 16'b1111111111110010;
        weights1[11484] <= 16'b1111111111111000;
        weights1[11485] <= 16'b0000000000000101;
        weights1[11486] <= 16'b0000000000100011;
        weights1[11487] <= 16'b0000000000110011;
        weights1[11488] <= 16'b0000000000101000;
        weights1[11489] <= 16'b1111111111111111;
        weights1[11490] <= 16'b1111111111101001;
        weights1[11491] <= 16'b1111111111101001;
        weights1[11492] <= 16'b1111111111001111;
        weights1[11493] <= 16'b0000000000000010;
        weights1[11494] <= 16'b0000000000011010;
        weights1[11495] <= 16'b0000000000101110;
        weights1[11496] <= 16'b1111111111110110;
        weights1[11497] <= 16'b1111111111110100;
        weights1[11498] <= 16'b1111111111101111;
        weights1[11499] <= 16'b1111111111100101;
        weights1[11500] <= 16'b0000000000001101;
        weights1[11501] <= 16'b0000000000001000;
        weights1[11502] <= 16'b0000000000011110;
        weights1[11503] <= 16'b0000000000010001;
        weights1[11504] <= 16'b0000000000010010;
        weights1[11505] <= 16'b0000000000010110;
        weights1[11506] <= 16'b0000000000001100;
        weights1[11507] <= 16'b0000000000000000;
        weights1[11508] <= 16'b1111111111100010;
        weights1[11509] <= 16'b1111111111011110;
        weights1[11510] <= 16'b1111111111110010;
        weights1[11511] <= 16'b1111111111101111;
        weights1[11512] <= 16'b0000000000000101;
        weights1[11513] <= 16'b0000000000011111;
        weights1[11514] <= 16'b0000000000101101;
        weights1[11515] <= 16'b0000000000100011;
        weights1[11516] <= 16'b0000000000010101;
        weights1[11517] <= 16'b1111111111101101;
        weights1[11518] <= 16'b1111111111011111;
        weights1[11519] <= 16'b1111111110111010;
        weights1[11520] <= 16'b1111111111010110;
        weights1[11521] <= 16'b0000000000010011;
        weights1[11522] <= 16'b0000000000100100;
        weights1[11523] <= 16'b0000000000100101;
        weights1[11524] <= 16'b1111111111110010;
        weights1[11525] <= 16'b1111111111010100;
        weights1[11526] <= 16'b1111111111100001;
        weights1[11527] <= 16'b1111111111100000;
        weights1[11528] <= 16'b1111111111111000;
        weights1[11529] <= 16'b1111111111110001;
        weights1[11530] <= 16'b0000000000011111;
        weights1[11531] <= 16'b0000000000100101;
        weights1[11532] <= 16'b0000000000010111;
        weights1[11533] <= 16'b0000000000011000;
        weights1[11534] <= 16'b0000000000001100;
        weights1[11535] <= 16'b0000000000000011;
        weights1[11536] <= 16'b1111111111101001;
        weights1[11537] <= 16'b1111111111110111;
        weights1[11538] <= 16'b0000000000000011;
        weights1[11539] <= 16'b0000000000010001;
        weights1[11540] <= 16'b0000000000111010;
        weights1[11541] <= 16'b0000000000101111;
        weights1[11542] <= 16'b0000000000101010;
        weights1[11543] <= 16'b0000000000000010;
        weights1[11544] <= 16'b1111111111111011;
        weights1[11545] <= 16'b1111111111010111;
        weights1[11546] <= 16'b1111111111000001;
        weights1[11547] <= 16'b1111111110110001;
        weights1[11548] <= 16'b1111111111101100;
        weights1[11549] <= 16'b0000000000010011;
        weights1[11550] <= 16'b0000000000110110;
        weights1[11551] <= 16'b0000000000101101;
        weights1[11552] <= 16'b0000000000000010;
        weights1[11553] <= 16'b1111111111010100;
        weights1[11554] <= 16'b1111111111001100;
        weights1[11555] <= 16'b1111111111011010;
        weights1[11556] <= 16'b1111111111011101;
        weights1[11557] <= 16'b1111111111110011;
        weights1[11558] <= 16'b0000000000100111;
        weights1[11559] <= 16'b0000000000100011;
        weights1[11560] <= 16'b0000000000110100;
        weights1[11561] <= 16'b0000000000010101;
        weights1[11562] <= 16'b0000000000000110;
        weights1[11563] <= 16'b0000000000000000;
        weights1[11564] <= 16'b0000000000001010;
        weights1[11565] <= 16'b0000000000010010;
        weights1[11566] <= 16'b0000000000011111;
        weights1[11567] <= 16'b0000000000100101;
        weights1[11568] <= 16'b0000000000101101;
        weights1[11569] <= 16'b0000000000110100;
        weights1[11570] <= 16'b0000000000101010;
        weights1[11571] <= 16'b1111111111110101;
        weights1[11572] <= 16'b1111111111011001;
        weights1[11573] <= 16'b1111111110011000;
        weights1[11574] <= 16'b1111111110001111;
        weights1[11575] <= 16'b1111111111000011;
        weights1[11576] <= 16'b0000000000000100;
        weights1[11577] <= 16'b0000000000101011;
        weights1[11578] <= 16'b0000000000111110;
        weights1[11579] <= 16'b0000000000100111;
        weights1[11580] <= 16'b0000000000000000;
        weights1[11581] <= 16'b1111111111010101;
        weights1[11582] <= 16'b1111111110011010;
        weights1[11583] <= 16'b1111111110111101;
        weights1[11584] <= 16'b1111111110111111;
        weights1[11585] <= 16'b1111111111111010;
        weights1[11586] <= 16'b0000000000001110;
        weights1[11587] <= 16'b0000000000101101;
        weights1[11588] <= 16'b0000000000101110;
        weights1[11589] <= 16'b0000000000011001;
        weights1[11590] <= 16'b0000000000001111;
        weights1[11591] <= 16'b0000000000001001;
        weights1[11592] <= 16'b0000000000010111;
        weights1[11593] <= 16'b0000000000011010;
        weights1[11594] <= 16'b0000000000101101;
        weights1[11595] <= 16'b0000000000101101;
        weights1[11596] <= 16'b0000000000101011;
        weights1[11597] <= 16'b0000000000011011;
        weights1[11598] <= 16'b1111111111111010;
        weights1[11599] <= 16'b1111111110110001;
        weights1[11600] <= 16'b1111111110000111;
        weights1[11601] <= 16'b1111111101110001;
        weights1[11602] <= 16'b1111111110000011;
        weights1[11603] <= 16'b1111111111010100;
        weights1[11604] <= 16'b0000000000100010;
        weights1[11605] <= 16'b0000000000101100;
        weights1[11606] <= 16'b0000000000100100;
        weights1[11607] <= 16'b0000000001000001;
        weights1[11608] <= 16'b1111111111110101;
        weights1[11609] <= 16'b1111111110111100;
        weights1[11610] <= 16'b1111111110100000;
        weights1[11611] <= 16'b1111111111000100;
        weights1[11612] <= 16'b1111111110111111;
        weights1[11613] <= 16'b1111111111001010;
        weights1[11614] <= 16'b1111111111110110;
        weights1[11615] <= 16'b0000000000010100;
        weights1[11616] <= 16'b0000000000100001;
        weights1[11617] <= 16'b0000000000011110;
        weights1[11618] <= 16'b0000000000010010;
        weights1[11619] <= 16'b0000000000001111;
        weights1[11620] <= 16'b0000000000001110;
        weights1[11621] <= 16'b0000000000011001;
        weights1[11622] <= 16'b0000000000011101;
        weights1[11623] <= 16'b0000000000001011;
        weights1[11624] <= 16'b0000000000000010;
        weights1[11625] <= 16'b1111111111000001;
        weights1[11626] <= 16'b1111111110101101;
        weights1[11627] <= 16'b1111111110000100;
        weights1[11628] <= 16'b1111111101101100;
        weights1[11629] <= 16'b1111111100111110;
        weights1[11630] <= 16'b1111111110110000;
        weights1[11631] <= 16'b0000000000010000;
        weights1[11632] <= 16'b0000000000110101;
        weights1[11633] <= 16'b0000000000111011;
        weights1[11634] <= 16'b0000000000111000;
        weights1[11635] <= 16'b0000000000101111;
        weights1[11636] <= 16'b0000000000010011;
        weights1[11637] <= 16'b1111111111001100;
        weights1[11638] <= 16'b1111111110100100;
        weights1[11639] <= 16'b1111111110111001;
        weights1[11640] <= 16'b1111111110111101;
        weights1[11641] <= 16'b1111111111000000;
        weights1[11642] <= 16'b1111111111101011;
        weights1[11643] <= 16'b0000000000000000;
        weights1[11644] <= 16'b0000000000010110;
        weights1[11645] <= 16'b0000000000001110;
        weights1[11646] <= 16'b0000000000011010;
        weights1[11647] <= 16'b0000000000010100;
        weights1[11648] <= 16'b0000000000001010;
        weights1[11649] <= 16'b0000000000000101;
        weights1[11650] <= 16'b0000000000000010;
        weights1[11651] <= 16'b1111111111110111;
        weights1[11652] <= 16'b1111111111011110;
        weights1[11653] <= 16'b1111111110110011;
        weights1[11654] <= 16'b1111111110100010;
        weights1[11655] <= 16'b1111111101111110;
        weights1[11656] <= 16'b1111111101001111;
        weights1[11657] <= 16'b1111111110000101;
        weights1[11658] <= 16'b0000000000010010;
        weights1[11659] <= 16'b0000000000110111;
        weights1[11660] <= 16'b0000000000110011;
        weights1[11661] <= 16'b0000000000010110;
        weights1[11662] <= 16'b0000000000001101;
        weights1[11663] <= 16'b0000000001000011;
        weights1[11664] <= 16'b1111111111100000;
        weights1[11665] <= 16'b1111111110101101;
        weights1[11666] <= 16'b1111111101101111;
        weights1[11667] <= 16'b1111111110101001;
        weights1[11668] <= 16'b1111111110111110;
        weights1[11669] <= 16'b1111111111000000;
        weights1[11670] <= 16'b1111111111011000;
        weights1[11671] <= 16'b1111111111101001;
        weights1[11672] <= 16'b1111111111111001;
        weights1[11673] <= 16'b0000000000000001;
        weights1[11674] <= 16'b0000000000001010;
        weights1[11675] <= 16'b0000000000001100;
        weights1[11676] <= 16'b1111111111111100;
        weights1[11677] <= 16'b1111111111110011;
        weights1[11678] <= 16'b1111111111101100;
        weights1[11679] <= 16'b1111111111010010;
        weights1[11680] <= 16'b1111111111001000;
        weights1[11681] <= 16'b1111111110110001;
        weights1[11682] <= 16'b1111111110000110;
        weights1[11683] <= 16'b1111111101111110;
        weights1[11684] <= 16'b1111111101110101;
        weights1[11685] <= 16'b1111111111001010;
        weights1[11686] <= 16'b0000000000000000;
        weights1[11687] <= 16'b0000000000100100;
        weights1[11688] <= 16'b0000000000101000;
        weights1[11689] <= 16'b0000000000011010;
        weights1[11690] <= 16'b0000000000110110;
        weights1[11691] <= 16'b0000000000111001;
        weights1[11692] <= 16'b0000000000001100;
        weights1[11693] <= 16'b1111111111000100;
        weights1[11694] <= 16'b1111111110100000;
        weights1[11695] <= 16'b1111111110101101;
        weights1[11696] <= 16'b1111111110111100;
        weights1[11697] <= 16'b1111111110110111;
        weights1[11698] <= 16'b1111111111001100;
        weights1[11699] <= 16'b1111111111011100;
        weights1[11700] <= 16'b1111111111101011;
        weights1[11701] <= 16'b0000000000000000;
        weights1[11702] <= 16'b0000000000001001;
        weights1[11703] <= 16'b0000000000001000;
        weights1[11704] <= 16'b1111111111110111;
        weights1[11705] <= 16'b1111111111101011;
        weights1[11706] <= 16'b1111111111100000;
        weights1[11707] <= 16'b1111111111001110;
        weights1[11708] <= 16'b1111111110111001;
        weights1[11709] <= 16'b1111111110110100;
        weights1[11710] <= 16'b1111111110100011;
        weights1[11711] <= 16'b1111111110010101;
        weights1[11712] <= 16'b1111111110111110;
        weights1[11713] <= 16'b1111111111111101;
        weights1[11714] <= 16'b0000000000011110;
        weights1[11715] <= 16'b0000000000101001;
        weights1[11716] <= 16'b0000000000101100;
        weights1[11717] <= 16'b0000000000100101;
        weights1[11718] <= 16'b0000000000101000;
        weights1[11719] <= 16'b0000000000010001;
        weights1[11720] <= 16'b1111111111101011;
        weights1[11721] <= 16'b1111111111001100;
        weights1[11722] <= 16'b1111111110101111;
        weights1[11723] <= 16'b1111111110111010;
        weights1[11724] <= 16'b1111111111000011;
        weights1[11725] <= 16'b1111111111000001;
        weights1[11726] <= 16'b1111111111011001;
        weights1[11727] <= 16'b1111111111011110;
        weights1[11728] <= 16'b1111111111101111;
        weights1[11729] <= 16'b1111111111111110;
        weights1[11730] <= 16'b0000000000000111;
        weights1[11731] <= 16'b0000000000000010;
        weights1[11732] <= 16'b1111111111111010;
        weights1[11733] <= 16'b1111111111110010;
        weights1[11734] <= 16'b1111111111100010;
        weights1[11735] <= 16'b1111111111001100;
        weights1[11736] <= 16'b1111111110110010;
        weights1[11737] <= 16'b1111111110100011;
        weights1[11738] <= 16'b1111111110010111;
        weights1[11739] <= 16'b1111111110100101;
        weights1[11740] <= 16'b1111111111100000;
        weights1[11741] <= 16'b0000000000000000;
        weights1[11742] <= 16'b0000000000101000;
        weights1[11743] <= 16'b0000000000100100;
        weights1[11744] <= 16'b0000000000110010;
        weights1[11745] <= 16'b0000000000101111;
        weights1[11746] <= 16'b0000000000011110;
        weights1[11747] <= 16'b0000000000010000;
        weights1[11748] <= 16'b0000000000000110;
        weights1[11749] <= 16'b1111111111010011;
        weights1[11750] <= 16'b1111111111000101;
        weights1[11751] <= 16'b1111111110110110;
        weights1[11752] <= 16'b1111111111000000;
        weights1[11753] <= 16'b1111111111001001;
        weights1[11754] <= 16'b1111111111011010;
        weights1[11755] <= 16'b1111111111100011;
        weights1[11756] <= 16'b1111111111110001;
        weights1[11757] <= 16'b0000000000000001;
        weights1[11758] <= 16'b0000000000001000;
        weights1[11759] <= 16'b0000000000001000;
        weights1[11760] <= 16'b0000000000000000;
        weights1[11761] <= 16'b0000000000000000;
        weights1[11762] <= 16'b0000000000000000;
        weights1[11763] <= 16'b0000000000000000;
        weights1[11764] <= 16'b0000000000000000;
        weights1[11765] <= 16'b1111111111111110;
        weights1[11766] <= 16'b0000000000000000;
        weights1[11767] <= 16'b0000000000000000;
        weights1[11768] <= 16'b0000000000000000;
        weights1[11769] <= 16'b0000000000000000;
        weights1[11770] <= 16'b0000000000000010;
        weights1[11771] <= 16'b0000000000000010;
        weights1[11772] <= 16'b0000000000000100;
        weights1[11773] <= 16'b0000000000000110;
        weights1[11774] <= 16'b0000000000001001;
        weights1[11775] <= 16'b0000000000001010;
        weights1[11776] <= 16'b0000000000000110;
        weights1[11777] <= 16'b0000000000001000;
        weights1[11778] <= 16'b0000000000000010;
        weights1[11779] <= 16'b1111111111111111;
        weights1[11780] <= 16'b0000000000000011;
        weights1[11781] <= 16'b0000000000000100;
        weights1[11782] <= 16'b0000000000000011;
        weights1[11783] <= 16'b0000000000000001;
        weights1[11784] <= 16'b0000000000000000;
        weights1[11785] <= 16'b1111111111111111;
        weights1[11786] <= 16'b0000000000000000;
        weights1[11787] <= 16'b0000000000000000;
        weights1[11788] <= 16'b0000000000000000;
        weights1[11789] <= 16'b0000000000000000;
        weights1[11790] <= 16'b0000000000000000;
        weights1[11791] <= 16'b1111111111111111;
        weights1[11792] <= 16'b1111111111111110;
        weights1[11793] <= 16'b1111111111111110;
        weights1[11794] <= 16'b1111111111111100;
        weights1[11795] <= 16'b1111111111111111;
        weights1[11796] <= 16'b1111111111111111;
        weights1[11797] <= 16'b0000000000000010;
        weights1[11798] <= 16'b0000000000000001;
        weights1[11799] <= 16'b0000000000000100;
        weights1[11800] <= 16'b0000000000001001;
        weights1[11801] <= 16'b0000000000001110;
        weights1[11802] <= 16'b0000000000001100;
        weights1[11803] <= 16'b0000000000001101;
        weights1[11804] <= 16'b0000000000001010;
        weights1[11805] <= 16'b0000000000001000;
        weights1[11806] <= 16'b0000000000001101;
        weights1[11807] <= 16'b0000000000000101;
        weights1[11808] <= 16'b0000000000000110;
        weights1[11809] <= 16'b0000000000001010;
        weights1[11810] <= 16'b0000000000000111;
        weights1[11811] <= 16'b0000000000000100;
        weights1[11812] <= 16'b1111111111111111;
        weights1[11813] <= 16'b1111111111111110;
        weights1[11814] <= 16'b1111111111111110;
        weights1[11815] <= 16'b0000000000000001;
        weights1[11816] <= 16'b0000000000000000;
        weights1[11817] <= 16'b0000000000000000;
        weights1[11818] <= 16'b0000000000000000;
        weights1[11819] <= 16'b1111111111111111;
        weights1[11820] <= 16'b1111111111111110;
        weights1[11821] <= 16'b1111111111111100;
        weights1[11822] <= 16'b1111111111111101;
        weights1[11823] <= 16'b0000000000000000;
        weights1[11824] <= 16'b1111111111111110;
        weights1[11825] <= 16'b1111111111111111;
        weights1[11826] <= 16'b0000000000000001;
        weights1[11827] <= 16'b0000000000000101;
        weights1[11828] <= 16'b0000000000001111;
        weights1[11829] <= 16'b0000000000010001;
        weights1[11830] <= 16'b0000000000001000;
        weights1[11831] <= 16'b0000000000001000;
        weights1[11832] <= 16'b0000000000000100;
        weights1[11833] <= 16'b0000000000001001;
        weights1[11834] <= 16'b0000000000001110;
        weights1[11835] <= 16'b0000000000001111;
        weights1[11836] <= 16'b0000000000000000;
        weights1[11837] <= 16'b0000000000000101;
        weights1[11838] <= 16'b0000000000001000;
        weights1[11839] <= 16'b0000000000001010;
        weights1[11840] <= 16'b0000000000000101;
        weights1[11841] <= 16'b0000000000000001;
        weights1[11842] <= 16'b0000000000000001;
        weights1[11843] <= 16'b0000000000000001;
        weights1[11844] <= 16'b1111111111111111;
        weights1[11845] <= 16'b1111111111111111;
        weights1[11846] <= 16'b1111111111111110;
        weights1[11847] <= 16'b1111111111111101;
        weights1[11848] <= 16'b1111111111111011;
        weights1[11849] <= 16'b1111111111110010;
        weights1[11850] <= 16'b1111111111110100;
        weights1[11851] <= 16'b1111111111111101;
        weights1[11852] <= 16'b1111111111111111;
        weights1[11853] <= 16'b1111111111111011;
        weights1[11854] <= 16'b1111111111111011;
        weights1[11855] <= 16'b1111111111110101;
        weights1[11856] <= 16'b1111111111110100;
        weights1[11857] <= 16'b1111111111110111;
        weights1[11858] <= 16'b1111111111110000;
        weights1[11859] <= 16'b1111111111111001;
        weights1[11860] <= 16'b1111111111111100;
        weights1[11861] <= 16'b1111111111110001;
        weights1[11862] <= 16'b1111111111110111;
        weights1[11863] <= 16'b1111111111111011;
        weights1[11864] <= 16'b1111111111110100;
        weights1[11865] <= 16'b1111111111111000;
        weights1[11866] <= 16'b0000000000000101;
        weights1[11867] <= 16'b0000000000000111;
        weights1[11868] <= 16'b0000000000000011;
        weights1[11869] <= 16'b0000000000000100;
        weights1[11870] <= 16'b1111111111111101;
        weights1[11871] <= 16'b1111111111111110;
        weights1[11872] <= 16'b1111111111111111;
        weights1[11873] <= 16'b1111111111111110;
        weights1[11874] <= 16'b1111111111111101;
        weights1[11875] <= 16'b1111111111111101;
        weights1[11876] <= 16'b1111111111111100;
        weights1[11877] <= 16'b1111111111111010;
        weights1[11878] <= 16'b1111111111110101;
        weights1[11879] <= 16'b1111111111110111;
        weights1[11880] <= 16'b1111111111111010;
        weights1[11881] <= 16'b0000000000000110;
        weights1[11882] <= 16'b0000000000001000;
        weights1[11883] <= 16'b1111111111111100;
        weights1[11884] <= 16'b1111111111111110;
        weights1[11885] <= 16'b0000000000000111;
        weights1[11886] <= 16'b0000000000000111;
        weights1[11887] <= 16'b1111111111111000;
        weights1[11888] <= 16'b1111111111111000;
        weights1[11889] <= 16'b1111111111111001;
        weights1[11890] <= 16'b1111111111110000;
        weights1[11891] <= 16'b1111111111111110;
        weights1[11892] <= 16'b1111111111101011;
        weights1[11893] <= 16'b1111111111110100;
        weights1[11894] <= 16'b0000000000000000;
        weights1[11895] <= 16'b1111111111111001;
        weights1[11896] <= 16'b1111111111111011;
        weights1[11897] <= 16'b1111111111111001;
        weights1[11898] <= 16'b1111111111111101;
        weights1[11899] <= 16'b1111111111111100;
        weights1[11900] <= 16'b1111111111111110;
        weights1[11901] <= 16'b1111111111111010;
        weights1[11902] <= 16'b1111111111111011;
        weights1[11903] <= 16'b1111111111110100;
        weights1[11904] <= 16'b1111111111111001;
        weights1[11905] <= 16'b1111111111110101;
        weights1[11906] <= 16'b0000000000000000;
        weights1[11907] <= 16'b1111111111111001;
        weights1[11908] <= 16'b1111111111100011;
        weights1[11909] <= 16'b0000000000000100;
        weights1[11910] <= 16'b1111111111111110;
        weights1[11911] <= 16'b0000000000010011;
        weights1[11912] <= 16'b0000000000000111;
        weights1[11913] <= 16'b1111111111011100;
        weights1[11914] <= 16'b1111111111111000;
        weights1[11915] <= 16'b1111111111111100;
        weights1[11916] <= 16'b0000000000001100;
        weights1[11917] <= 16'b0000000000001100;
        weights1[11918] <= 16'b0000000000001101;
        weights1[11919] <= 16'b0000000000000000;
        weights1[11920] <= 16'b0000000000001111;
        weights1[11921] <= 16'b0000000000000101;
        weights1[11922] <= 16'b1111111111110111;
        weights1[11923] <= 16'b1111111111110010;
        weights1[11924] <= 16'b1111111111101011;
        weights1[11925] <= 16'b1111111111110000;
        weights1[11926] <= 16'b1111111111111000;
        weights1[11927] <= 16'b1111111111111010;
        weights1[11928] <= 16'b1111111111111100;
        weights1[11929] <= 16'b1111111111111000;
        weights1[11930] <= 16'b1111111111110111;
        weights1[11931] <= 16'b1111111111111001;
        weights1[11932] <= 16'b1111111111101101;
        weights1[11933] <= 16'b1111111111011011;
        weights1[11934] <= 16'b0000000000001101;
        weights1[11935] <= 16'b1111111111101110;
        weights1[11936] <= 16'b1111111111110010;
        weights1[11937] <= 16'b0000000000001001;
        weights1[11938] <= 16'b0000000000100000;
        weights1[11939] <= 16'b1111111111110000;
        weights1[11940] <= 16'b1111111111101101;
        weights1[11941] <= 16'b1111111111111110;
        weights1[11942] <= 16'b1111111111101001;
        weights1[11943] <= 16'b1111111111111110;
        weights1[11944] <= 16'b1111111111110110;
        weights1[11945] <= 16'b1111111111101111;
        weights1[11946] <= 16'b0000000000011011;
        weights1[11947] <= 16'b1111111111110111;
        weights1[11948] <= 16'b0000000000001110;
        weights1[11949] <= 16'b0000000000010100;
        weights1[11950] <= 16'b0000000000001100;
        weights1[11951] <= 16'b1111111111111011;
        weights1[11952] <= 16'b0000000000001101;
        weights1[11953] <= 16'b1111111111110100;
        weights1[11954] <= 16'b0000000000000001;
        weights1[11955] <= 16'b1111111111111111;
        weights1[11956] <= 16'b1111111111111000;
        weights1[11957] <= 16'b1111111111110101;
        weights1[11958] <= 16'b1111111111110001;
        weights1[11959] <= 16'b1111111111101110;
        weights1[11960] <= 16'b1111111111110010;
        weights1[11961] <= 16'b1111111111111010;
        weights1[11962] <= 16'b0000000000001000;
        weights1[11963] <= 16'b0000000000000111;
        weights1[11964] <= 16'b0000000000001111;
        weights1[11965] <= 16'b1111111111110101;
        weights1[11966] <= 16'b1111111111110111;
        weights1[11967] <= 16'b0000000000000101;
        weights1[11968] <= 16'b1111111111111011;
        weights1[11969] <= 16'b1111111111110011;
        weights1[11970] <= 16'b1111111111111111;
        weights1[11971] <= 16'b0000000000010010;
        weights1[11972] <= 16'b1111111111111100;
        weights1[11973] <= 16'b1111111111111011;
        weights1[11974] <= 16'b0000000000001100;
        weights1[11975] <= 16'b1111111111110000;
        weights1[11976] <= 16'b1111111111111101;
        weights1[11977] <= 16'b0000000000011001;
        weights1[11978] <= 16'b1111111111110010;
        weights1[11979] <= 16'b1111111111101100;
        weights1[11980] <= 16'b1111111111110110;
        weights1[11981] <= 16'b1111111111111011;
        weights1[11982] <= 16'b0000000000000010;
        weights1[11983] <= 16'b1111111111111111;
        weights1[11984] <= 16'b1111111111111001;
        weights1[11985] <= 16'b1111111111111011;
        weights1[11986] <= 16'b1111111111110011;
        weights1[11987] <= 16'b1111111111101110;
        weights1[11988] <= 16'b1111111111111000;
        weights1[11989] <= 16'b1111111111101000;
        weights1[11990] <= 16'b0000000000010001;
        weights1[11991] <= 16'b0000000000001011;
        weights1[11992] <= 16'b1111111111010001;
        weights1[11993] <= 16'b1111111111100100;
        weights1[11994] <= 16'b1111111111110111;
        weights1[11995] <= 16'b1111111111111000;
        weights1[11996] <= 16'b0000000000000100;
        weights1[11997] <= 16'b0000000000010001;
        weights1[11998] <= 16'b1111111111110101;
        weights1[11999] <= 16'b1111111111100011;
        weights1[12000] <= 16'b0000000000001001;
        weights1[12001] <= 16'b0000000000000100;
        weights1[12002] <= 16'b1111111111110101;
        weights1[12003] <= 16'b0000000000001000;
        weights1[12004] <= 16'b0000000000000100;
        weights1[12005] <= 16'b1111111111101000;
        weights1[12006] <= 16'b0000000000000010;
        weights1[12007] <= 16'b1111111111101011;
        weights1[12008] <= 16'b1111111111110011;
        weights1[12009] <= 16'b1111111111111011;
        weights1[12010] <= 16'b0000000000000000;
        weights1[12011] <= 16'b1111111111111111;
        weights1[12012] <= 16'b1111111111111111;
        weights1[12013] <= 16'b1111111111110111;
        weights1[12014] <= 16'b1111111111101110;
        weights1[12015] <= 16'b1111111111110000;
        weights1[12016] <= 16'b1111111111110010;
        weights1[12017] <= 16'b1111111111100010;
        weights1[12018] <= 16'b1111111111101011;
        weights1[12019] <= 16'b1111111111111000;
        weights1[12020] <= 16'b1111111111111100;
        weights1[12021] <= 16'b0000000000000011;
        weights1[12022] <= 16'b1111111111110001;
        weights1[12023] <= 16'b1111111111111010;
        weights1[12024] <= 16'b1111111111111100;
        weights1[12025] <= 16'b1111111111111001;
        weights1[12026] <= 16'b1111111111110000;
        weights1[12027] <= 16'b1111111111111111;
        weights1[12028] <= 16'b0000000000000001;
        weights1[12029] <= 16'b1111111111101001;
        weights1[12030] <= 16'b0000000000000001;
        weights1[12031] <= 16'b1111111111110010;
        weights1[12032] <= 16'b0000000000000000;
        weights1[12033] <= 16'b0000000000000100;
        weights1[12034] <= 16'b0000000000001001;
        weights1[12035] <= 16'b0000000000000100;
        weights1[12036] <= 16'b1111111111101110;
        weights1[12037] <= 16'b0000000000000101;
        weights1[12038] <= 16'b0000000000010000;
        weights1[12039] <= 16'b0000000000000100;
        weights1[12040] <= 16'b1111111111111000;
        weights1[12041] <= 16'b1111111111101110;
        weights1[12042] <= 16'b1111111111111000;
        weights1[12043] <= 16'b0000000000000001;
        weights1[12044] <= 16'b1111111111111110;
        weights1[12045] <= 16'b1111111111110001;
        weights1[12046] <= 16'b1111111111111101;
        weights1[12047] <= 16'b1111111111111010;
        weights1[12048] <= 16'b1111111111101001;
        weights1[12049] <= 16'b0000000000001010;
        weights1[12050] <= 16'b1111111111101110;
        weights1[12051] <= 16'b1111111111110110;
        weights1[12052] <= 16'b1111111111111010;
        weights1[12053] <= 16'b1111111111111101;
        weights1[12054] <= 16'b1111111111111000;
        weights1[12055] <= 16'b1111111111110110;
        weights1[12056] <= 16'b0000000000001010;
        weights1[12057] <= 16'b1111111111111100;
        weights1[12058] <= 16'b0000000000000000;
        weights1[12059] <= 16'b1111111111111101;
        weights1[12060] <= 16'b1111111111111111;
        weights1[12061] <= 16'b1111111111111100;
        weights1[12062] <= 16'b1111111111111000;
        weights1[12063] <= 16'b0000000000000000;
        weights1[12064] <= 16'b1111111111100111;
        weights1[12065] <= 16'b1111111111111010;
        weights1[12066] <= 16'b1111111111110111;
        weights1[12067] <= 16'b1111111111110110;
        weights1[12068] <= 16'b1111111111110100;
        weights1[12069] <= 16'b1111111111110010;
        weights1[12070] <= 16'b1111111111110001;
        weights1[12071] <= 16'b1111111111110100;
        weights1[12072] <= 16'b0000000000000100;
        weights1[12073] <= 16'b1111111111101111;
        weights1[12074] <= 16'b0000000000001110;
        weights1[12075] <= 16'b1111111111100101;
        weights1[12076] <= 16'b1111111111101110;
        weights1[12077] <= 16'b1111111111110100;
        weights1[12078] <= 16'b1111111111110111;
        weights1[12079] <= 16'b1111111111110110;
        weights1[12080] <= 16'b1111111111101110;
        weights1[12081] <= 16'b1111111111111011;
        weights1[12082] <= 16'b1111111111100001;
        weights1[12083] <= 16'b1111111111111000;
        weights1[12084] <= 16'b1111111111100001;
        weights1[12085] <= 16'b1111111111110101;
        weights1[12086] <= 16'b1111111111101101;
        weights1[12087] <= 16'b0000000000000001;
        weights1[12088] <= 16'b1111111111110001;
        weights1[12089] <= 16'b0000000000000000;
        weights1[12090] <= 16'b1111111111110101;
        weights1[12091] <= 16'b1111111111101100;
        weights1[12092] <= 16'b1111111111100111;
        weights1[12093] <= 16'b1111111111101100;
        weights1[12094] <= 16'b1111111111110100;
        weights1[12095] <= 16'b1111111111111001;
        weights1[12096] <= 16'b1111111111110111;
        weights1[12097] <= 16'b1111111111110101;
        weights1[12098] <= 16'b1111111111111101;
        weights1[12099] <= 16'b1111111111110011;
        weights1[12100] <= 16'b1111111111111111;
        weights1[12101] <= 16'b1111111111111001;
        weights1[12102] <= 16'b1111111111110000;
        weights1[12103] <= 16'b1111111111101001;
        weights1[12104] <= 16'b0000000000000110;
        weights1[12105] <= 16'b0000000000000100;
        weights1[12106] <= 16'b1111111111110001;
        weights1[12107] <= 16'b1111111111101011;
        weights1[12108] <= 16'b0000000000000011;
        weights1[12109] <= 16'b1111111111101101;
        weights1[12110] <= 16'b1111111111101110;
        weights1[12111] <= 16'b1111111111110010;
        weights1[12112] <= 16'b1111111111110100;
        weights1[12113] <= 16'b1111111111100000;
        weights1[12114] <= 16'b1111111111011011;
        weights1[12115] <= 16'b1111111111111000;
        weights1[12116] <= 16'b1111111111100101;
        weights1[12117] <= 16'b1111111111110100;
        weights1[12118] <= 16'b1111111111100001;
        weights1[12119] <= 16'b1111111111011100;
        weights1[12120] <= 16'b1111111111011000;
        weights1[12121] <= 16'b1111111111101100;
        weights1[12122] <= 16'b1111111111101011;
        weights1[12123] <= 16'b1111111111110010;
        weights1[12124] <= 16'b1111111111101110;
        weights1[12125] <= 16'b0000000000000000;
        weights1[12126] <= 16'b1111111111111000;
        weights1[12127] <= 16'b1111111111110010;
        weights1[12128] <= 16'b1111111111110110;
        weights1[12129] <= 16'b1111111111100000;
        weights1[12130] <= 16'b0000000000000011;
        weights1[12131] <= 16'b1111111111110111;
        weights1[12132] <= 16'b1111111111100000;
        weights1[12133] <= 16'b1111111111100010;
        weights1[12134] <= 16'b1111111111110000;
        weights1[12135] <= 16'b1111111111100110;
        weights1[12136] <= 16'b1111111111101111;
        weights1[12137] <= 16'b0000000000001010;
        weights1[12138] <= 16'b0000000000000011;
        weights1[12139] <= 16'b1111111111101000;
        weights1[12140] <= 16'b1111111111110000;
        weights1[12141] <= 16'b1111111111111001;
        weights1[12142] <= 16'b0000000000000000;
        weights1[12143] <= 16'b1111111111101111;
        weights1[12144] <= 16'b1111111111100111;
        weights1[12145] <= 16'b1111111111010110;
        weights1[12146] <= 16'b1111111111011011;
        weights1[12147] <= 16'b1111111111011011;
        weights1[12148] <= 16'b1111111111011010;
        weights1[12149] <= 16'b1111111111110001;
        weights1[12150] <= 16'b1111111111101100;
        weights1[12151] <= 16'b1111111111111000;
        weights1[12152] <= 16'b1111111111110111;
        weights1[12153] <= 16'b1111111111111111;
        weights1[12154] <= 16'b1111111111110000;
        weights1[12155] <= 16'b1111111111101010;
        weights1[12156] <= 16'b0000000000010010;
        weights1[12157] <= 16'b1111111111100010;
        weights1[12158] <= 16'b1111111111101010;
        weights1[12159] <= 16'b1111111111101001;
        weights1[12160] <= 16'b1111111111100110;
        weights1[12161] <= 16'b1111111111110101;
        weights1[12162] <= 16'b1111111111111110;
        weights1[12163] <= 16'b1111111111110000;
        weights1[12164] <= 16'b1111111111101100;
        weights1[12165] <= 16'b1111111111110001;
        weights1[12166] <= 16'b1111111111111100;
        weights1[12167] <= 16'b0000000000001011;
        weights1[12168] <= 16'b1111111111110011;
        weights1[12169] <= 16'b1111111111101001;
        weights1[12170] <= 16'b1111111111100100;
        weights1[12171] <= 16'b1111111111110110;
        weights1[12172] <= 16'b1111111111101110;
        weights1[12173] <= 16'b1111111111101000;
        weights1[12174] <= 16'b1111111111001000;
        weights1[12175] <= 16'b1111111111011010;
        weights1[12176] <= 16'b1111111111100100;
        weights1[12177] <= 16'b1111111111100010;
        weights1[12178] <= 16'b1111111111100111;
        weights1[12179] <= 16'b0000000000000101;
        weights1[12180] <= 16'b1111111111111001;
        weights1[12181] <= 16'b0000000000000101;
        weights1[12182] <= 16'b1111111111101110;
        weights1[12183] <= 16'b1111111111110001;
        weights1[12184] <= 16'b1111111111111101;
        weights1[12185] <= 16'b1111111111110010;
        weights1[12186] <= 16'b1111111111110000;
        weights1[12187] <= 16'b1111111111101010;
        weights1[12188] <= 16'b0000000000001010;
        weights1[12189] <= 16'b1111111111101100;
        weights1[12190] <= 16'b1111111111110111;
        weights1[12191] <= 16'b0000000000001000;
        weights1[12192] <= 16'b0000000000001010;
        weights1[12193] <= 16'b1111111111110111;
        weights1[12194] <= 16'b1111111111110011;
        weights1[12195] <= 16'b0000000000001111;
        weights1[12196] <= 16'b0000000000000010;
        weights1[12197] <= 16'b1111111111111100;
        weights1[12198] <= 16'b1111111111010100;
        weights1[12199] <= 16'b1111111111101001;
        weights1[12200] <= 16'b1111111111100000;
        weights1[12201] <= 16'b1111111111101110;
        weights1[12202] <= 16'b1111111111100000;
        weights1[12203] <= 16'b1111111111101010;
        weights1[12204] <= 16'b1111111111011100;
        weights1[12205] <= 16'b1111111111010111;
        weights1[12206] <= 16'b1111111111111110;
        weights1[12207] <= 16'b0000000000011011;
        weights1[12208] <= 16'b1111111111110000;
        weights1[12209] <= 16'b1111111111101111;
        weights1[12210] <= 16'b1111111111101001;
        weights1[12211] <= 16'b1111111111100110;
        weights1[12212] <= 16'b1111111111101101;
        weights1[12213] <= 16'b1111111111100010;
        weights1[12214] <= 16'b1111111111111100;
        weights1[12215] <= 16'b1111111111111111;
        weights1[12216] <= 16'b0000000000001000;
        weights1[12217] <= 16'b0000000000010100;
        weights1[12218] <= 16'b0000000000001010;
        weights1[12219] <= 16'b1111111111111100;
        weights1[12220] <= 16'b1111111111110100;
        weights1[12221] <= 16'b1111111111110010;
        weights1[12222] <= 16'b1111111111110011;
        weights1[12223] <= 16'b1111111111110011;
        weights1[12224] <= 16'b1111111111101110;
        weights1[12225] <= 16'b1111111111111000;
        weights1[12226] <= 16'b1111111111111100;
        weights1[12227] <= 16'b1111111111111101;
        weights1[12228] <= 16'b1111111111100000;
        weights1[12229] <= 16'b1111111111110011;
        weights1[12230] <= 16'b1111111111101000;
        weights1[12231] <= 16'b1111111111110001;
        weights1[12232] <= 16'b1111111111101111;
        weights1[12233] <= 16'b1111111111110010;
        weights1[12234] <= 16'b0000000000100000;
        weights1[12235] <= 16'b0000000000101001;
        weights1[12236] <= 16'b1111111111110001;
        weights1[12237] <= 16'b1111111111101011;
        weights1[12238] <= 16'b1111111111110001;
        weights1[12239] <= 16'b1111111111010100;
        weights1[12240] <= 16'b1111111111011100;
        weights1[12241] <= 16'b1111111111101011;
        weights1[12242] <= 16'b0000000000001001;
        weights1[12243] <= 16'b0000000000000000;
        weights1[12244] <= 16'b1111111111110101;
        weights1[12245] <= 16'b1111111111111111;
        weights1[12246] <= 16'b1111111111111111;
        weights1[12247] <= 16'b1111111111110000;
        weights1[12248] <= 16'b1111111111111110;
        weights1[12249] <= 16'b1111111111111010;
        weights1[12250] <= 16'b1111111111111010;
        weights1[12251] <= 16'b1111111111101011;
        weights1[12252] <= 16'b1111111111111100;
        weights1[12253] <= 16'b0000000000000000;
        weights1[12254] <= 16'b0000000000000000;
        weights1[12255] <= 16'b1111111111111101;
        weights1[12256] <= 16'b1111111111100110;
        weights1[12257] <= 16'b1111111111111010;
        weights1[12258] <= 16'b1111111111101011;
        weights1[12259] <= 16'b1111111111101100;
        weights1[12260] <= 16'b0000000000000100;
        weights1[12261] <= 16'b0000000000011000;
        weights1[12262] <= 16'b0000000000100100;
        weights1[12263] <= 16'b0000000000111101;
        weights1[12264] <= 16'b1111111111111010;
        weights1[12265] <= 16'b1111111111101011;
        weights1[12266] <= 16'b1111111111111100;
        weights1[12267] <= 16'b1111111111110101;
        weights1[12268] <= 16'b1111111111111001;
        weights1[12269] <= 16'b0000000000000001;
        weights1[12270] <= 16'b1111111111111000;
        weights1[12271] <= 16'b1111111111111110;
        weights1[12272] <= 16'b1111111111111110;
        weights1[12273] <= 16'b1111111111111110;
        weights1[12274] <= 16'b1111111111111010;
        weights1[12275] <= 16'b1111111111110100;
        weights1[12276] <= 16'b1111111111111001;
        weights1[12277] <= 16'b1111111111111010;
        weights1[12278] <= 16'b1111111111100000;
        weights1[12279] <= 16'b1111111111111001;
        weights1[12280] <= 16'b1111111111111000;
        weights1[12281] <= 16'b0000000000001101;
        weights1[12282] <= 16'b0000000000010000;
        weights1[12283] <= 16'b1111111111111110;
        weights1[12284] <= 16'b1111111111011010;
        weights1[12285] <= 16'b1111111111011100;
        weights1[12286] <= 16'b1111111111110101;
        weights1[12287] <= 16'b1111111111110000;
        weights1[12288] <= 16'b0000000000000010;
        weights1[12289] <= 16'b0000000000110011;
        weights1[12290] <= 16'b0000000000111000;
        weights1[12291] <= 16'b0000000000101110;
        weights1[12292] <= 16'b0000000000001000;
        weights1[12293] <= 16'b1111111111111100;
        weights1[12294] <= 16'b1111111111101111;
        weights1[12295] <= 16'b1111111111111100;
        weights1[12296] <= 16'b0000000000001000;
        weights1[12297] <= 16'b1111111111110111;
        weights1[12298] <= 16'b0000000000000001;
        weights1[12299] <= 16'b1111111111110101;
        weights1[12300] <= 16'b1111111111111101;
        weights1[12301] <= 16'b1111111111011110;
        weights1[12302] <= 16'b1111111111110100;
        weights1[12303] <= 16'b1111111111111110;
        weights1[12304] <= 16'b0000000000000111;
        weights1[12305] <= 16'b1111111111111011;
        weights1[12306] <= 16'b1111111111100011;
        weights1[12307] <= 16'b1111111111100110;
        weights1[12308] <= 16'b1111111111110001;
        weights1[12309] <= 16'b1111111111110001;
        weights1[12310] <= 16'b1111111111111010;
        weights1[12311] <= 16'b1111111111110010;
        weights1[12312] <= 16'b1111111111101000;
        weights1[12313] <= 16'b1111111111110110;
        weights1[12314] <= 16'b0000000000001101;
        weights1[12315] <= 16'b0000000000010101;
        weights1[12316] <= 16'b0000000000011110;
        weights1[12317] <= 16'b0000000001001000;
        weights1[12318] <= 16'b0000000000110110;
        weights1[12319] <= 16'b0000000000100100;
        weights1[12320] <= 16'b0000000000010111;
        weights1[12321] <= 16'b0000000000001110;
        weights1[12322] <= 16'b0000000000001110;
        weights1[12323] <= 16'b0000000000010010;
        weights1[12324] <= 16'b0000000000001111;
        weights1[12325] <= 16'b1111111111101111;
        weights1[12326] <= 16'b1111111111111110;
        weights1[12327] <= 16'b0000000000011011;
        weights1[12328] <= 16'b1111111111101001;
        weights1[12329] <= 16'b0000000000001001;
        weights1[12330] <= 16'b1111111111100110;
        weights1[12331] <= 16'b1111111111100101;
        weights1[12332] <= 16'b1111111111101000;
        weights1[12333] <= 16'b1111111111010001;
        weights1[12334] <= 16'b1111111111101101;
        weights1[12335] <= 16'b1111111111101000;
        weights1[12336] <= 16'b1111111111011101;
        weights1[12337] <= 16'b1111111111010010;
        weights1[12338] <= 16'b1111111111101010;
        weights1[12339] <= 16'b0000000000001010;
        weights1[12340] <= 16'b1111111111101011;
        weights1[12341] <= 16'b0000000000001110;
        weights1[12342] <= 16'b0000000000100001;
        weights1[12343] <= 16'b0000000000110110;
        weights1[12344] <= 16'b0000000000111110;
        weights1[12345] <= 16'b0000000001010011;
        weights1[12346] <= 16'b0000000000111000;
        weights1[12347] <= 16'b0000000000100111;
        weights1[12348] <= 16'b0000000000101000;
        weights1[12349] <= 16'b0000000000101101;
        weights1[12350] <= 16'b0000000000100001;
        weights1[12351] <= 16'b0000000000100100;
        weights1[12352] <= 16'b0000000000010100;
        weights1[12353] <= 16'b1111111111111000;
        weights1[12354] <= 16'b1111111111111100;
        weights1[12355] <= 16'b0000000000001001;
        weights1[12356] <= 16'b0000000000000000;
        weights1[12357] <= 16'b1111111111100110;
        weights1[12358] <= 16'b1111111111010000;
        weights1[12359] <= 16'b1111111111011100;
        weights1[12360] <= 16'b1111111111010100;
        weights1[12361] <= 16'b0000000000001001;
        weights1[12362] <= 16'b0000000000000000;
        weights1[12363] <= 16'b0000000000000011;
        weights1[12364] <= 16'b1111111111100111;
        weights1[12365] <= 16'b1111111111100010;
        weights1[12366] <= 16'b1111111111111001;
        weights1[12367] <= 16'b0000000000010011;
        weights1[12368] <= 16'b0000000000101011;
        weights1[12369] <= 16'b0000000000111001;
        weights1[12370] <= 16'b0000000001100001;
        weights1[12371] <= 16'b0000000001010001;
        weights1[12372] <= 16'b0000000001100010;
        weights1[12373] <= 16'b0000000001010110;
        weights1[12374] <= 16'b0000000000110011;
        weights1[12375] <= 16'b0000000000110000;
        weights1[12376] <= 16'b0000000000110011;
        weights1[12377] <= 16'b0000000001000010;
        weights1[12378] <= 16'b0000000001000011;
        weights1[12379] <= 16'b0000000000110000;
        weights1[12380] <= 16'b0000000000100001;
        weights1[12381] <= 16'b0000000000110101;
        weights1[12382] <= 16'b0000000000101100;
        weights1[12383] <= 16'b0000000000001100;
        weights1[12384] <= 16'b0000000000001001;
        weights1[12385] <= 16'b0000000000101111;
        weights1[12386] <= 16'b0000000000001000;
        weights1[12387] <= 16'b0000000000011011;
        weights1[12388] <= 16'b0000000000100010;
        weights1[12389] <= 16'b0000000000000000;
        weights1[12390] <= 16'b0000000000101001;
        weights1[12391] <= 16'b0000000000110110;
        weights1[12392] <= 16'b0000000001001010;
        weights1[12393] <= 16'b0000000000101111;
        weights1[12394] <= 16'b0000000000111010;
        weights1[12395] <= 16'b0000000001011011;
        weights1[12396] <= 16'b0000000001011101;
        weights1[12397] <= 16'b0000000001101011;
        weights1[12398] <= 16'b0000000001100000;
        weights1[12399] <= 16'b0000000001100010;
        weights1[12400] <= 16'b0000000001010000;
        weights1[12401] <= 16'b0000000001010001;
        weights1[12402] <= 16'b0000000000110100;
        weights1[12403] <= 16'b0000000000101010;
        weights1[12404] <= 16'b0000000000110010;
        weights1[12405] <= 16'b0000000000111111;
        weights1[12406] <= 16'b0000000001001011;
        weights1[12407] <= 16'b0000000001011011;
        weights1[12408] <= 16'b0000000001001100;
        weights1[12409] <= 16'b0000000001011011;
        weights1[12410] <= 16'b0000000001011100;
        weights1[12411] <= 16'b0000000001001100;
        weights1[12412] <= 16'b0000000001101010;
        weights1[12413] <= 16'b0000000001101010;
        weights1[12414] <= 16'b0000000001010100;
        weights1[12415] <= 16'b0000000001101100;
        weights1[12416] <= 16'b0000000001100101;
        weights1[12417] <= 16'b0000000001000001;
        weights1[12418] <= 16'b0000000001001110;
        weights1[12419] <= 16'b0000000001011110;
        weights1[12420] <= 16'b0000000001100010;
        weights1[12421] <= 16'b0000000001101010;
        weights1[12422] <= 16'b0000000001101000;
        weights1[12423] <= 16'b0000000001100011;
        weights1[12424] <= 16'b0000000001010100;
        weights1[12425] <= 16'b0000000001000001;
        weights1[12426] <= 16'b0000000001010011;
        weights1[12427] <= 16'b0000000000101111;
        weights1[12428] <= 16'b0000000000110011;
        weights1[12429] <= 16'b0000000000111101;
        weights1[12430] <= 16'b0000000000100101;
        weights1[12431] <= 16'b0000000000011010;
        weights1[12432] <= 16'b0000000000101010;
        weights1[12433] <= 16'b0000000000111010;
        weights1[12434] <= 16'b0000000000111010;
        weights1[12435] <= 16'b0000000001001111;
        weights1[12436] <= 16'b0000000001000110;
        weights1[12437] <= 16'b0000000001010000;
        weights1[12438] <= 16'b0000000001000100;
        weights1[12439] <= 16'b0000000001010011;
        weights1[12440] <= 16'b0000000001100010;
        weights1[12441] <= 16'b0000000001001111;
        weights1[12442] <= 16'b0000000001110000;
        weights1[12443] <= 16'b0000000001101101;
        weights1[12444] <= 16'b0000000001011110;
        weights1[12445] <= 16'b0000000001010000;
        weights1[12446] <= 16'b0000000001001000;
        weights1[12447] <= 16'b0000000001001100;
        weights1[12448] <= 16'b0000000001011011;
        weights1[12449] <= 16'b0000000001001001;
        weights1[12450] <= 16'b0000000001000111;
        weights1[12451] <= 16'b0000000001000100;
        weights1[12452] <= 16'b0000000000110111;
        weights1[12453] <= 16'b0000000000101100;
        weights1[12454] <= 16'b0000000000111010;
        weights1[12455] <= 16'b0000000000010110;
        weights1[12456] <= 16'b0000000000101100;
        weights1[12457] <= 16'b0000000000110010;
        weights1[12458] <= 16'b0000000000011111;
        weights1[12459] <= 16'b0000000000001001;
        weights1[12460] <= 16'b0000000000011000;
        weights1[12461] <= 16'b0000000000101011;
        weights1[12462] <= 16'b0000000000100101;
        weights1[12463] <= 16'b0000000000101110;
        weights1[12464] <= 16'b0000000000110001;
        weights1[12465] <= 16'b0000000000100011;
        weights1[12466] <= 16'b0000000000101101;
        weights1[12467] <= 16'b0000000000011110;
        weights1[12468] <= 16'b0000000000110100;
        weights1[12469] <= 16'b0000000000101001;
        weights1[12470] <= 16'b0000000000111111;
        weights1[12471] <= 16'b0000000000110111;
        weights1[12472] <= 16'b0000000001001010;
        weights1[12473] <= 16'b0000000000110100;
        weights1[12474] <= 16'b0000000001000101;
        weights1[12475] <= 16'b0000000000110111;
        weights1[12476] <= 16'b0000000000110011;
        weights1[12477] <= 16'b0000000000011111;
        weights1[12478] <= 16'b0000000000010110;
        weights1[12479] <= 16'b0000000000100001;
        weights1[12480] <= 16'b0000000000110011;
        weights1[12481] <= 16'b0000000000010100;
        weights1[12482] <= 16'b0000000000011001;
        weights1[12483] <= 16'b0000000000010110;
        weights1[12484] <= 16'b0000000000011110;
        weights1[12485] <= 16'b0000000000011110;
        weights1[12486] <= 16'b0000000000010000;
        weights1[12487] <= 16'b0000000000000010;
        weights1[12488] <= 16'b0000000000000100;
        weights1[12489] <= 16'b0000000000000111;
        weights1[12490] <= 16'b0000000000010000;
        weights1[12491] <= 16'b0000000000010110;
        weights1[12492] <= 16'b0000000000010100;
        weights1[12493] <= 16'b0000000000011101;
        weights1[12494] <= 16'b0000000000010101;
        weights1[12495] <= 16'b0000000000011010;
        weights1[12496] <= 16'b0000000000010010;
        weights1[12497] <= 16'b0000000000010010;
        weights1[12498] <= 16'b0000000000100000;
        weights1[12499] <= 16'b0000000000001110;
        weights1[12500] <= 16'b0000000000100011;
        weights1[12501] <= 16'b0000000000011011;
        weights1[12502] <= 16'b0000000000010111;
        weights1[12503] <= 16'b0000000000010001;
        weights1[12504] <= 16'b0000000000001110;
        weights1[12505] <= 16'b0000000000001111;
        weights1[12506] <= 16'b0000000000100011;
        weights1[12507] <= 16'b0000000000011001;
        weights1[12508] <= 16'b0000000000010101;
        weights1[12509] <= 16'b0000000000011111;
        weights1[12510] <= 16'b0000000000010111;
        weights1[12511] <= 16'b0000000000010100;
        weights1[12512] <= 16'b0000000000010100;
        weights1[12513] <= 16'b0000000000000010;
        weights1[12514] <= 16'b0000000000000110;
        weights1[12515] <= 16'b1111111111111100;
        weights1[12516] <= 16'b1111111111111011;
        weights1[12517] <= 16'b0000000000000001;
        weights1[12518] <= 16'b0000000000000001;
        weights1[12519] <= 16'b1111111111111111;
        weights1[12520] <= 16'b0000000000001010;
        weights1[12521] <= 16'b0000000000010111;
        weights1[12522] <= 16'b0000000000001100;
        weights1[12523] <= 16'b0000000000001110;
        weights1[12524] <= 16'b0000000000001101;
        weights1[12525] <= 16'b0000000000001100;
        weights1[12526] <= 16'b0000000000011010;
        weights1[12527] <= 16'b0000000000011100;
        weights1[12528] <= 16'b0000000000010010;
        weights1[12529] <= 16'b0000000000010010;
        weights1[12530] <= 16'b0000000000010101;
        weights1[12531] <= 16'b0000000000100011;
        weights1[12532] <= 16'b0000000000001111;
        weights1[12533] <= 16'b0000000000001000;
        weights1[12534] <= 16'b0000000000101010;
        weights1[12535] <= 16'b0000000000101001;
        weights1[12536] <= 16'b0000000000001100;
        weights1[12537] <= 16'b0000000000001001;
        weights1[12538] <= 16'b0000000000010010;
        weights1[12539] <= 16'b0000000000000111;
        weights1[12540] <= 16'b0000000000000101;
        weights1[12541] <= 16'b0000000000001001;
        weights1[12542] <= 16'b1111111111111110;
        weights1[12543] <= 16'b1111111111111001;
        weights1[12544] <= 16'b0000000000000000;
        weights1[12545] <= 16'b1111111111111111;
        weights1[12546] <= 16'b1111111111111101;
        weights1[12547] <= 16'b1111111111111010;
        weights1[12548] <= 16'b1111111111110001;
        weights1[12549] <= 16'b1111111111110001;
        weights1[12550] <= 16'b1111111111101010;
        weights1[12551] <= 16'b1111111111101000;
        weights1[12552] <= 16'b1111111111101011;
        weights1[12553] <= 16'b1111111111100000;
        weights1[12554] <= 16'b1111111111011011;
        weights1[12555] <= 16'b1111111111011001;
        weights1[12556] <= 16'b1111111111011100;
        weights1[12557] <= 16'b1111111111011010;
        weights1[12558] <= 16'b1111111111100001;
        weights1[12559] <= 16'b1111111111100000;
        weights1[12560] <= 16'b1111111111011100;
        weights1[12561] <= 16'b1111111111101001;
        weights1[12562] <= 16'b1111111111100111;
        weights1[12563] <= 16'b1111111111100110;
        weights1[12564] <= 16'b1111111111101111;
        weights1[12565] <= 16'b1111111111101101;
        weights1[12566] <= 16'b1111111111110110;
        weights1[12567] <= 16'b1111111111111000;
        weights1[12568] <= 16'b1111111111110101;
        weights1[12569] <= 16'b1111111111111001;
        weights1[12570] <= 16'b1111111111111101;
        weights1[12571] <= 16'b1111111111111111;
        weights1[12572] <= 16'b0000000000000000;
        weights1[12573] <= 16'b1111111111111101;
        weights1[12574] <= 16'b1111111111110111;
        weights1[12575] <= 16'b1111111111110001;
        weights1[12576] <= 16'b1111111111101010;
        weights1[12577] <= 16'b1111111111100101;
        weights1[12578] <= 16'b1111111111100000;
        weights1[12579] <= 16'b1111111111011000;
        weights1[12580] <= 16'b1111111111011110;
        weights1[12581] <= 16'b1111111111001111;
        weights1[12582] <= 16'b1111111111001010;
        weights1[12583] <= 16'b1111111111001001;
        weights1[12584] <= 16'b1111111111000110;
        weights1[12585] <= 16'b1111111111000111;
        weights1[12586] <= 16'b1111111111001001;
        weights1[12587] <= 16'b1111111111000100;
        weights1[12588] <= 16'b1111111111000101;
        weights1[12589] <= 16'b1111111111010001;
        weights1[12590] <= 16'b1111111111010111;
        weights1[12591] <= 16'b1111111111010111;
        weights1[12592] <= 16'b1111111111011000;
        weights1[12593] <= 16'b1111111111011110;
        weights1[12594] <= 16'b1111111111100001;
        weights1[12595] <= 16'b1111111111101011;
        weights1[12596] <= 16'b1111111111101100;
        weights1[12597] <= 16'b1111111111110011;
        weights1[12598] <= 16'b1111111111111100;
        weights1[12599] <= 16'b1111111111111110;
        weights1[12600] <= 16'b0000000000000000;
        weights1[12601] <= 16'b1111111111111011;
        weights1[12602] <= 16'b1111111111101110;
        weights1[12603] <= 16'b1111111111101011;
        weights1[12604] <= 16'b1111111111100101;
        weights1[12605] <= 16'b1111111111011101;
        weights1[12606] <= 16'b1111111111010000;
        weights1[12607] <= 16'b1111111111001000;
        weights1[12608] <= 16'b1111111111001010;
        weights1[12609] <= 16'b1111111110111101;
        weights1[12610] <= 16'b1111111110111000;
        weights1[12611] <= 16'b1111111110101010;
        weights1[12612] <= 16'b1111111110100011;
        weights1[12613] <= 16'b1111111110101100;
        weights1[12614] <= 16'b1111111110101001;
        weights1[12615] <= 16'b1111111110001111;
        weights1[12616] <= 16'b1111111110100111;
        weights1[12617] <= 16'b1111111110101001;
        weights1[12618] <= 16'b1111111110101101;
        weights1[12619] <= 16'b1111111110101100;
        weights1[12620] <= 16'b1111111111000101;
        weights1[12621] <= 16'b1111111111010010;
        weights1[12622] <= 16'b1111111111010100;
        weights1[12623] <= 16'b1111111111011000;
        weights1[12624] <= 16'b1111111111100011;
        weights1[12625] <= 16'b1111111111110000;
        weights1[12626] <= 16'b1111111111111100;
        weights1[12627] <= 16'b1111111111110111;
        weights1[12628] <= 16'b0000000000000001;
        weights1[12629] <= 16'b1111111111111001;
        weights1[12630] <= 16'b1111111111110010;
        weights1[12631] <= 16'b1111111111100100;
        weights1[12632] <= 16'b1111111111100010;
        weights1[12633] <= 16'b1111111111010101;
        weights1[12634] <= 16'b1111111111000110;
        weights1[12635] <= 16'b1111111110110110;
        weights1[12636] <= 16'b1111111111000110;
        weights1[12637] <= 16'b1111111110101101;
        weights1[12638] <= 16'b1111111110011110;
        weights1[12639] <= 16'b1111111110100000;
        weights1[12640] <= 16'b1111111110001010;
        weights1[12641] <= 16'b1111111101110001;
        weights1[12642] <= 16'b1111111110011111;
        weights1[12643] <= 16'b1111111110011010;
        weights1[12644] <= 16'b1111111110111110;
        weights1[12645] <= 16'b1111111111000001;
        weights1[12646] <= 16'b1111111110101001;
        weights1[12647] <= 16'b1111111111000111;
        weights1[12648] <= 16'b1111111111000011;
        weights1[12649] <= 16'b1111111111010101;
        weights1[12650] <= 16'b1111111111011010;
        weights1[12651] <= 16'b1111111111001011;
        weights1[12652] <= 16'b1111111111100001;
        weights1[12653] <= 16'b1111111111100111;
        weights1[12654] <= 16'b1111111111110010;
        weights1[12655] <= 16'b1111111111110101;
        weights1[12656] <= 16'b0000000000000001;
        weights1[12657] <= 16'b1111111111111001;
        weights1[12658] <= 16'b1111111111110010;
        weights1[12659] <= 16'b1111111111100011;
        weights1[12660] <= 16'b1111111111011111;
        weights1[12661] <= 16'b1111111111001011;
        weights1[12662] <= 16'b1111111111010111;
        weights1[12663] <= 16'b1111111111001101;
        weights1[12664] <= 16'b1111111111001010;
        weights1[12665] <= 16'b1111111111100100;
        weights1[12666] <= 16'b1111111111010110;
        weights1[12667] <= 16'b1111111111100001;
        weights1[12668] <= 16'b1111111111100101;
        weights1[12669] <= 16'b1111111111011010;
        weights1[12670] <= 16'b1111111111011101;
        weights1[12671] <= 16'b1111111111111001;
        weights1[12672] <= 16'b1111111111110000;
        weights1[12673] <= 16'b1111111111101100;
        weights1[12674] <= 16'b1111111111101100;
        weights1[12675] <= 16'b1111111111100011;
        weights1[12676] <= 16'b0000000000000001;
        weights1[12677] <= 16'b1111111111011110;
        weights1[12678] <= 16'b1111111111101100;
        weights1[12679] <= 16'b1111111111101011;
        weights1[12680] <= 16'b1111111111010110;
        weights1[12681] <= 16'b1111111111001011;
        weights1[12682] <= 16'b1111111111101001;
        weights1[12683] <= 16'b1111111111110001;
        weights1[12684] <= 16'b0000000000000101;
        weights1[12685] <= 16'b1111111111111111;
        weights1[12686] <= 16'b1111111111110001;
        weights1[12687] <= 16'b1111111111110001;
        weights1[12688] <= 16'b1111111111111000;
        weights1[12689] <= 16'b1111111111111000;
        weights1[12690] <= 16'b0000000000000101;
        weights1[12691] <= 16'b0000000000001001;
        weights1[12692] <= 16'b0000000000010101;
        weights1[12693] <= 16'b0000000000001110;
        weights1[12694] <= 16'b0000000000000101;
        weights1[12695] <= 16'b0000000000110110;
        weights1[12696] <= 16'b0000000000111010;
        weights1[12697] <= 16'b0000000000011100;
        weights1[12698] <= 16'b0000000000011100;
        weights1[12699] <= 16'b0000000000100100;
        weights1[12700] <= 16'b0000000000001111;
        weights1[12701] <= 16'b0000000000000101;
        weights1[12702] <= 16'b0000000000000010;
        weights1[12703] <= 16'b0000000000000110;
        weights1[12704] <= 16'b1111111111110010;
        weights1[12705] <= 16'b1111111111110110;
        weights1[12706] <= 16'b1111111111110100;
        weights1[12707] <= 16'b1111111111110110;
        weights1[12708] <= 16'b1111111111101001;
        weights1[12709] <= 16'b1111111111000101;
        weights1[12710] <= 16'b1111111111010110;
        weights1[12711] <= 16'b1111111111100010;
        weights1[12712] <= 16'b0000000000000100;
        weights1[12713] <= 16'b0000000000000100;
        weights1[12714] <= 16'b0000000000000010;
        weights1[12715] <= 16'b0000000000010000;
        weights1[12716] <= 16'b0000000000011101;
        weights1[12717] <= 16'b0000000000110010;
        weights1[12718] <= 16'b0000000001000010;
        weights1[12719] <= 16'b0000000001010010;
        weights1[12720] <= 16'b0000000001010100;
        weights1[12721] <= 16'b0000000001001001;
        weights1[12722] <= 16'b0000000000110100;
        weights1[12723] <= 16'b0000000000101000;
        weights1[12724] <= 16'b0000000000011101;
        weights1[12725] <= 16'b0000000000111101;
        weights1[12726] <= 16'b0000000000101100;
        weights1[12727] <= 16'b0000000000101100;
        weights1[12728] <= 16'b0000000000001111;
        weights1[12729] <= 16'b0000000000010000;
        weights1[12730] <= 16'b0000000000101000;
        weights1[12731] <= 16'b0000000000011011;
        weights1[12732] <= 16'b0000000000000000;
        weights1[12733] <= 16'b0000000000010001;
        weights1[12734] <= 16'b0000000000010101;
        weights1[12735] <= 16'b1111111111110011;
        weights1[12736] <= 16'b1111111111101111;
        weights1[12737] <= 16'b1111111111101101;
        weights1[12738] <= 16'b1111111111101001;
        weights1[12739] <= 16'b1111111111100100;
        weights1[12740] <= 16'b0000000000000111;
        weights1[12741] <= 16'b0000000000010101;
        weights1[12742] <= 16'b0000000000100100;
        weights1[12743] <= 16'b0000000000101010;
        weights1[12744] <= 16'b0000000001000101;
        weights1[12745] <= 16'b0000000000111100;
        weights1[12746] <= 16'b0000000001000010;
        weights1[12747] <= 16'b0000000001001100;
        weights1[12748] <= 16'b0000000000100110;
        weights1[12749] <= 16'b0000000000100100;
        weights1[12750] <= 16'b0000000001001000;
        weights1[12751] <= 16'b0000000000111100;
        weights1[12752] <= 16'b0000000000111000;
        weights1[12753] <= 16'b0000000000101011;
        weights1[12754] <= 16'b0000000000100010;
        weights1[12755] <= 16'b0000000000001110;
        weights1[12756] <= 16'b0000000000011110;
        weights1[12757] <= 16'b0000000000100001;
        weights1[12758] <= 16'b0000000000011001;
        weights1[12759] <= 16'b1111111111111101;
        weights1[12760] <= 16'b0000000000011101;
        weights1[12761] <= 16'b0000000000001110;
        weights1[12762] <= 16'b0000000000100100;
        weights1[12763] <= 16'b0000000000001110;
        weights1[12764] <= 16'b0000000000000101;
        weights1[12765] <= 16'b0000000000000010;
        weights1[12766] <= 16'b1111111111100001;
        weights1[12767] <= 16'b1111111111100101;
        weights1[12768] <= 16'b0000000000010011;
        weights1[12769] <= 16'b0000000000011110;
        weights1[12770] <= 16'b0000000000101000;
        weights1[12771] <= 16'b0000000000101111;
        weights1[12772] <= 16'b0000000000110111;
        weights1[12773] <= 16'b0000000000101111;
        weights1[12774] <= 16'b0000000000110101;
        weights1[12775] <= 16'b0000000000001101;
        weights1[12776] <= 16'b0000000000100110;
        weights1[12777] <= 16'b0000000000110110;
        weights1[12778] <= 16'b0000000000111001;
        weights1[12779] <= 16'b0000000000101110;
        weights1[12780] <= 16'b0000000001001001;
        weights1[12781] <= 16'b0000000000110011;
        weights1[12782] <= 16'b0000000001001101;
        weights1[12783] <= 16'b0000000000111000;
        weights1[12784] <= 16'b0000000001010110;
        weights1[12785] <= 16'b0000000000100110;
        weights1[12786] <= 16'b0000000000110110;
        weights1[12787] <= 16'b0000000000011011;
        weights1[12788] <= 16'b0000000000010111;
        weights1[12789] <= 16'b1111111111111111;
        weights1[12790] <= 16'b0000000000000111;
        weights1[12791] <= 16'b1111111111111110;
        weights1[12792] <= 16'b0000000000001111;
        weights1[12793] <= 16'b1111111111110100;
        weights1[12794] <= 16'b1111111111101010;
        weights1[12795] <= 16'b1111111111101001;
        weights1[12796] <= 16'b0000000000010001;
        weights1[12797] <= 16'b0000000000011010;
        weights1[12798] <= 16'b0000000000010001;
        weights1[12799] <= 16'b0000000000100100;
        weights1[12800] <= 16'b0000000000001011;
        weights1[12801] <= 16'b0000000000010100;
        weights1[12802] <= 16'b0000000000010101;
        weights1[12803] <= 16'b1111111111110000;
        weights1[12804] <= 16'b1111111111100101;
        weights1[12805] <= 16'b1111111111100100;
        weights1[12806] <= 16'b1111111111111100;
        weights1[12807] <= 16'b1111111111101001;
        weights1[12808] <= 16'b0000000000000001;
        weights1[12809] <= 16'b0000000000010100;
        weights1[12810] <= 16'b0000000000001101;
        weights1[12811] <= 16'b0000000000011110;
        weights1[12812] <= 16'b0000000000011111;
        weights1[12813] <= 16'b0000000000100010;
        weights1[12814] <= 16'b0000000000101000;
        weights1[12815] <= 16'b0000000000000111;
        weights1[12816] <= 16'b0000000000101001;
        weights1[12817] <= 16'b0000000000010000;
        weights1[12818] <= 16'b0000000000001010;
        weights1[12819] <= 16'b0000000000011100;
        weights1[12820] <= 16'b1111111111111110;
        weights1[12821] <= 16'b0000000000010010;
        weights1[12822] <= 16'b0000000000000111;
        weights1[12823] <= 16'b1111111111101100;
        weights1[12824] <= 16'b0000000000001101;
        weights1[12825] <= 16'b0000000000000000;
        weights1[12826] <= 16'b1111111111111011;
        weights1[12827] <= 16'b1111111111111011;
        weights1[12828] <= 16'b1111111111100001;
        weights1[12829] <= 16'b1111111111111011;
        weights1[12830] <= 16'b1111111111110001;
        weights1[12831] <= 16'b1111111111110000;
        weights1[12832] <= 16'b1111111111011000;
        weights1[12833] <= 16'b1111111111011101;
        weights1[12834] <= 16'b1111111111010100;
        weights1[12835] <= 16'b1111111111000101;
        weights1[12836] <= 16'b1111111111011111;
        weights1[12837] <= 16'b1111111111000011;
        weights1[12838] <= 16'b1111111111011010;
        weights1[12839] <= 16'b1111111111100100;
        weights1[12840] <= 16'b0000000000011000;
        weights1[12841] <= 16'b1111111111110101;
        weights1[12842] <= 16'b0000000000101011;
        weights1[12843] <= 16'b0000000000100011;
        weights1[12844] <= 16'b0000000000100100;
        weights1[12845] <= 16'b0000000000100101;
        weights1[12846] <= 16'b0000000000100100;
        weights1[12847] <= 16'b0000000000011101;
        weights1[12848] <= 16'b0000000000010011;
        weights1[12849] <= 16'b0000000000100000;
        weights1[12850] <= 16'b0000000000000100;
        weights1[12851] <= 16'b0000000000000100;
        weights1[12852] <= 16'b0000000000000000;
        weights1[12853] <= 16'b1111111111111000;
        weights1[12854] <= 16'b1111111111110000;
        weights1[12855] <= 16'b1111111111010010;
        weights1[12856] <= 16'b1111111111001101;
        weights1[12857] <= 16'b1111111111100101;
        weights1[12858] <= 16'b1111111111000000;
        weights1[12859] <= 16'b1111111111000111;
        weights1[12860] <= 16'b1111111111100110;
        weights1[12861] <= 16'b1111111111010001;
        weights1[12862] <= 16'b1111111111011001;
        weights1[12863] <= 16'b1111111111011010;
        weights1[12864] <= 16'b1111111111010101;
        weights1[12865] <= 16'b1111111111100000;
        weights1[12866] <= 16'b1111111111011000;
        weights1[12867] <= 16'b1111111111000011;
        weights1[12868] <= 16'b1111111111100100;
        weights1[12869] <= 16'b0000000000000001;
        weights1[12870] <= 16'b0000000000001000;
        weights1[12871] <= 16'b0000000000000111;
        weights1[12872] <= 16'b0000000000010111;
        weights1[12873] <= 16'b0000000000010001;
        weights1[12874] <= 16'b0000000000101011;
        weights1[12875] <= 16'b0000000000101001;
        weights1[12876] <= 16'b0000000000010100;
        weights1[12877] <= 16'b0000000000010101;
        weights1[12878] <= 16'b0000000000010011;
        weights1[12879] <= 16'b0000000000000100;
        weights1[12880] <= 16'b1111111111110110;
        weights1[12881] <= 16'b1111111111100111;
        weights1[12882] <= 16'b1111111111101001;
        weights1[12883] <= 16'b1111111111011100;
        weights1[12884] <= 16'b1111111111011000;
        weights1[12885] <= 16'b1111111111000111;
        weights1[12886] <= 16'b1111111110110110;
        weights1[12887] <= 16'b1111111111101100;
        weights1[12888] <= 16'b1111111111101111;
        weights1[12889] <= 16'b0000000000000011;
        weights1[12890] <= 16'b1111111111101100;
        weights1[12891] <= 16'b1111111111110010;
        weights1[12892] <= 16'b1111111111101000;
        weights1[12893] <= 16'b1111111111011001;
        weights1[12894] <= 16'b1111111111010111;
        weights1[12895] <= 16'b1111111111101010;
        weights1[12896] <= 16'b1111111111100000;
        weights1[12897] <= 16'b1111111111110010;
        weights1[12898] <= 16'b0000000000001111;
        weights1[12899] <= 16'b0000000000001011;
        weights1[12900] <= 16'b0000000000000010;
        weights1[12901] <= 16'b0000000000001101;
        weights1[12902] <= 16'b0000000000001011;
        weights1[12903] <= 16'b0000000000000001;
        weights1[12904] <= 16'b1111111111110010;
        weights1[12905] <= 16'b0000000000011101;
        weights1[12906] <= 16'b0000000000001000;
        weights1[12907] <= 16'b0000000000000110;
        weights1[12908] <= 16'b1111111111101000;
        weights1[12909] <= 16'b1111111111011111;
        weights1[12910] <= 16'b1111111111011111;
        weights1[12911] <= 16'b1111111111011101;
        weights1[12912] <= 16'b1111111111011101;
        weights1[12913] <= 16'b1111111111011000;
        weights1[12914] <= 16'b1111111111000010;
        weights1[12915] <= 16'b1111111111101110;
        weights1[12916] <= 16'b0000000000001001;
        weights1[12917] <= 16'b1111111111111101;
        weights1[12918] <= 16'b1111111111111110;
        weights1[12919] <= 16'b0000000000000101;
        weights1[12920] <= 16'b0000000000001000;
        weights1[12921] <= 16'b1111111111111001;
        weights1[12922] <= 16'b1111111111100011;
        weights1[12923] <= 16'b0000000000000001;
        weights1[12924] <= 16'b0000000000001010;
        weights1[12925] <= 16'b1111111111101100;
        weights1[12926] <= 16'b0000000000000100;
        weights1[12927] <= 16'b0000000000000001;
        weights1[12928] <= 16'b0000000000010001;
        weights1[12929] <= 16'b0000000000011001;
        weights1[12930] <= 16'b0000000000000001;
        weights1[12931] <= 16'b0000000000001111;
        weights1[12932] <= 16'b0000000000000101;
        weights1[12933] <= 16'b0000000000001011;
        weights1[12934] <= 16'b0000000000001001;
        weights1[12935] <= 16'b0000000000001100;
        weights1[12936] <= 16'b1111111111100110;
        weights1[12937] <= 16'b1111111111011100;
        weights1[12938] <= 16'b1111111111101000;
        weights1[12939] <= 16'b1111111111100010;
        weights1[12940] <= 16'b0000000000000111;
        weights1[12941] <= 16'b1111111111011011;
        weights1[12942] <= 16'b1111111111011010;
        weights1[12943] <= 16'b1111111111111110;
        weights1[12944] <= 16'b1111111111110010;
        weights1[12945] <= 16'b1111111111100101;
        weights1[12946] <= 16'b1111111111111001;
        weights1[12947] <= 16'b0000000000000010;
        weights1[12948] <= 16'b1111111111111101;
        weights1[12949] <= 16'b0000000000001010;
        weights1[12950] <= 16'b0000000000000100;
        weights1[12951] <= 16'b1111111111110100;
        weights1[12952] <= 16'b1111111111100100;
        weights1[12953] <= 16'b1111111111101110;
        weights1[12954] <= 16'b1111111111100111;
        weights1[12955] <= 16'b1111111111111001;
        weights1[12956] <= 16'b1111111111110111;
        weights1[12957] <= 16'b0000000000001000;
        weights1[12958] <= 16'b0000000000011001;
        weights1[12959] <= 16'b1111111111111101;
        weights1[12960] <= 16'b0000000000011110;
        weights1[12961] <= 16'b0000000000000110;
        weights1[12962] <= 16'b0000000000001000;
        weights1[12963] <= 16'b0000000000001011;
        weights1[12964] <= 16'b1111111111110100;
        weights1[12965] <= 16'b1111111111101001;
        weights1[12966] <= 16'b1111111111100010;
        weights1[12967] <= 16'b1111111111101001;
        weights1[12968] <= 16'b0000000000001000;
        weights1[12969] <= 16'b0000000000000010;
        weights1[12970] <= 16'b0000000000001100;
        weights1[12971] <= 16'b1111111111101010;
        weights1[12972] <= 16'b1111111111110000;
        weights1[12973] <= 16'b1111111111111000;
        weights1[12974] <= 16'b0000000000001000;
        weights1[12975] <= 16'b1111111111110001;
        weights1[12976] <= 16'b0000000000000110;
        weights1[12977] <= 16'b1111111111111110;
        weights1[12978] <= 16'b0000000000001000;
        weights1[12979] <= 16'b1111111111110100;
        weights1[12980] <= 16'b1111111111110010;
        weights1[12981] <= 16'b0000000000000101;
        weights1[12982] <= 16'b1111111111111001;
        weights1[12983] <= 16'b1111111111011111;
        weights1[12984] <= 16'b1111111111111000;
        weights1[12985] <= 16'b1111111111111010;
        weights1[12986] <= 16'b0000000000011010;
        weights1[12987] <= 16'b0000000000000100;
        weights1[12988] <= 16'b0000000000000110;
        weights1[12989] <= 16'b1111111111110111;
        weights1[12990] <= 16'b1111111111110100;
        weights1[12991] <= 16'b0000000000000110;
        weights1[12992] <= 16'b1111111111111010;
        weights1[12993] <= 16'b1111111111111101;
        weights1[12994] <= 16'b1111111111111000;
        weights1[12995] <= 16'b1111111111111010;
        weights1[12996] <= 16'b1111111111111010;
        weights1[12997] <= 16'b0000000000010010;
        weights1[12998] <= 16'b1111111111110110;
        weights1[12999] <= 16'b1111111111111001;
        weights1[13000] <= 16'b0000000000000011;
        weights1[13001] <= 16'b1111111111111100;
        weights1[13002] <= 16'b0000000000010010;
        weights1[13003] <= 16'b0000000000010111;
        weights1[13004] <= 16'b1111111111111001;
        weights1[13005] <= 16'b0000000000000001;
        weights1[13006] <= 16'b1111111111110110;
        weights1[13007] <= 16'b0000000000000100;
        weights1[13008] <= 16'b0000000000001000;
        weights1[13009] <= 16'b1111111111101100;
        weights1[13010] <= 16'b1111111111101000;
        weights1[13011] <= 16'b1111111111011000;
        weights1[13012] <= 16'b0000000000000101;
        weights1[13013] <= 16'b1111111111111110;
        weights1[13014] <= 16'b0000000000000011;
        weights1[13015] <= 16'b0000000000001111;
        weights1[13016] <= 16'b0000000000001011;
        weights1[13017] <= 16'b0000000000000011;
        weights1[13018] <= 16'b0000000000000000;
        weights1[13019] <= 16'b0000000000000001;
        weights1[13020] <= 16'b1111111111110110;
        weights1[13021] <= 16'b0000000000000010;
        weights1[13022] <= 16'b1111111111111100;
        weights1[13023] <= 16'b1111111111111101;
        weights1[13024] <= 16'b0000000000011101;
        weights1[13025] <= 16'b0000000000010010;
        weights1[13026] <= 16'b0000000000000111;
        weights1[13027] <= 16'b1111111111111100;
        weights1[13028] <= 16'b0000000000001000;
        weights1[13029] <= 16'b0000000000000011;
        weights1[13030] <= 16'b1111111111100100;
        weights1[13031] <= 16'b0000000000000001;
        weights1[13032] <= 16'b0000000000000010;
        weights1[13033] <= 16'b1111111111100110;
        weights1[13034] <= 16'b1111111111101110;
        weights1[13035] <= 16'b1111111111111101;
        weights1[13036] <= 16'b0000000000000000;
        weights1[13037] <= 16'b1111111111111100;
        weights1[13038] <= 16'b1111111111110111;
        weights1[13039] <= 16'b1111111111110010;
        weights1[13040] <= 16'b1111111111101110;
        weights1[13041] <= 16'b1111111111110001;
        weights1[13042] <= 16'b1111111111110000;
        weights1[13043] <= 16'b0000000000001001;
        weights1[13044] <= 16'b0000000000000000;
        weights1[13045] <= 16'b1111111111111011;
        weights1[13046] <= 16'b1111111111111101;
        weights1[13047] <= 16'b0000000000000111;
        weights1[13048] <= 16'b1111111111110111;
        weights1[13049] <= 16'b0000000000000001;
        weights1[13050] <= 16'b0000000000001000;
        weights1[13051] <= 16'b1111111111111001;
        weights1[13052] <= 16'b0000000000001110;
        weights1[13053] <= 16'b0000000000010011;
        weights1[13054] <= 16'b0000000000010000;
        weights1[13055] <= 16'b1111111111110110;
        weights1[13056] <= 16'b0000000000001111;
        weights1[13057] <= 16'b0000000000000110;
        weights1[13058] <= 16'b0000000000000100;
        weights1[13059] <= 16'b1111111111111010;
        weights1[13060] <= 16'b0000000000000101;
        weights1[13061] <= 16'b0000000000001001;
        weights1[13062] <= 16'b1111111111100101;
        weights1[13063] <= 16'b1111111111110000;
        weights1[13064] <= 16'b0000000000001001;
        weights1[13065] <= 16'b0000000000010000;
        weights1[13066] <= 16'b0000000000010111;
        weights1[13067] <= 16'b0000000000001000;
        weights1[13068] <= 16'b1111111111110110;
        weights1[13069] <= 16'b1111111111101011;
        weights1[13070] <= 16'b0000000000001100;
        weights1[13071] <= 16'b0000000000000011;
        weights1[13072] <= 16'b0000000000000111;
        weights1[13073] <= 16'b1111111111111000;
        weights1[13074] <= 16'b1111111111111011;
        weights1[13075] <= 16'b0000000000001111;
        weights1[13076] <= 16'b1111111111111011;
        weights1[13077] <= 16'b1111111111110101;
        weights1[13078] <= 16'b0000000000000111;
        weights1[13079] <= 16'b1111111111111101;
        weights1[13080] <= 16'b1111111111111100;
        weights1[13081] <= 16'b0000000000000110;
        weights1[13082] <= 16'b1111111111111001;
        weights1[13083] <= 16'b1111111111111110;
        weights1[13084] <= 16'b0000000000010010;
        weights1[13085] <= 16'b0000000000000100;
        weights1[13086] <= 16'b0000000000000100;
        weights1[13087] <= 16'b1111111111110010;
        weights1[13088] <= 16'b0000000000011010;
        weights1[13089] <= 16'b1111111111101011;
        weights1[13090] <= 16'b1111111111111110;
        weights1[13091] <= 16'b0000000000000100;
        weights1[13092] <= 16'b1111111111101110;
        weights1[13093] <= 16'b1111111111111101;
        weights1[13094] <= 16'b1111111111110000;
        weights1[13095] <= 16'b0000000000001111;
        weights1[13096] <= 16'b0000000000001100;
        weights1[13097] <= 16'b0000000000000111;
        weights1[13098] <= 16'b0000000000000010;
        weights1[13099] <= 16'b0000000000011111;
        weights1[13100] <= 16'b0000000000001010;
        weights1[13101] <= 16'b0000000000000010;
        weights1[13102] <= 16'b0000000000000001;
        weights1[13103] <= 16'b1111111111110110;
        weights1[13104] <= 16'b0000000000000110;
        weights1[13105] <= 16'b0000000000001100;
        weights1[13106] <= 16'b1111111111111001;
        weights1[13107] <= 16'b1111111111111111;
        weights1[13108] <= 16'b0000000000010000;
        weights1[13109] <= 16'b1111111111111110;
        weights1[13110] <= 16'b1111111111111111;
        weights1[13111] <= 16'b0000000000011101;
        weights1[13112] <= 16'b0000000000001001;
        weights1[13113] <= 16'b1111111111110111;
        weights1[13114] <= 16'b0000000000001000;
        weights1[13115] <= 16'b1111111111110111;
        weights1[13116] <= 16'b1111111111111011;
        weights1[13117] <= 16'b1111111111100111;
        weights1[13118] <= 16'b0000000000000110;
        weights1[13119] <= 16'b1111111111110110;
        weights1[13120] <= 16'b1111111111111110;
        weights1[13121] <= 16'b1111111111110000;
        weights1[13122] <= 16'b0000000000000001;
        weights1[13123] <= 16'b0000000000000101;
        weights1[13124] <= 16'b1111111111111010;
        weights1[13125] <= 16'b0000000000011101;
        weights1[13126] <= 16'b1111111111101001;
        weights1[13127] <= 16'b0000000000000100;
        weights1[13128] <= 16'b0000000000000111;
        weights1[13129] <= 16'b0000000000000100;
        weights1[13130] <= 16'b1111111111110111;
        weights1[13131] <= 16'b1111111111111011;
        weights1[13132] <= 16'b1111111111111110;
        weights1[13133] <= 16'b1111111111111110;
        weights1[13134] <= 16'b1111111111111001;
        weights1[13135] <= 16'b1111111111100011;
        weights1[13136] <= 16'b0000000000001101;
        weights1[13137] <= 16'b0000000000001111;
        weights1[13138] <= 16'b0000000000000101;
        weights1[13139] <= 16'b1111111111110111;
        weights1[13140] <= 16'b1111111111110101;
        weights1[13141] <= 16'b0000000000001111;
        weights1[13142] <= 16'b1111111111111111;
        weights1[13143] <= 16'b0000000000010010;
        weights1[13144] <= 16'b0000000000001100;
        weights1[13145] <= 16'b0000000000000000;
        weights1[13146] <= 16'b1111111111111110;
        weights1[13147] <= 16'b0000000000010111;
        weights1[13148] <= 16'b1111111111111001;
        weights1[13149] <= 16'b0000000000001000;
        weights1[13150] <= 16'b0000000000000010;
        weights1[13151] <= 16'b0000000000001000;
        weights1[13152] <= 16'b1111111111101011;
        weights1[13153] <= 16'b1111111111111000;
        weights1[13154] <= 16'b1111111111110111;
        weights1[13155] <= 16'b1111111111111001;
        weights1[13156] <= 16'b1111111111110100;
        weights1[13157] <= 16'b1111111111111100;
        weights1[13158] <= 16'b1111111111111101;
        weights1[13159] <= 16'b0000000000000010;
        weights1[13160] <= 16'b0000000000000010;
        weights1[13161] <= 16'b1111111111111111;
        weights1[13162] <= 16'b1111111111111111;
        weights1[13163] <= 16'b0000000000000100;
        weights1[13164] <= 16'b1111111111110011;
        weights1[13165] <= 16'b1111111111101111;
        weights1[13166] <= 16'b1111111111101000;
        weights1[13167] <= 16'b0000000000000000;
        weights1[13168] <= 16'b0000000000000010;
        weights1[13169] <= 16'b0000000000010100;
        weights1[13170] <= 16'b1111111111110111;
        weights1[13171] <= 16'b1111111111101000;
        weights1[13172] <= 16'b0000000000000010;
        weights1[13173] <= 16'b0000000000010111;
        weights1[13174] <= 16'b1111111111110110;
        weights1[13175] <= 16'b0000000000000001;
        weights1[13176] <= 16'b1111111111111111;
        weights1[13177] <= 16'b1111111111110101;
        weights1[13178] <= 16'b0000000000000111;
        weights1[13179] <= 16'b0000000000010101;
        weights1[13180] <= 16'b1111111111111001;
        weights1[13181] <= 16'b1111111111111010;
        weights1[13182] <= 16'b0000000000001000;
        weights1[13183] <= 16'b0000000000000100;
        weights1[13184] <= 16'b1111111111111111;
        weights1[13185] <= 16'b1111111111111001;
        weights1[13186] <= 16'b1111111111111010;
        weights1[13187] <= 16'b1111111111111100;
        weights1[13188] <= 16'b1111111111111011;
        weights1[13189] <= 16'b1111111111111111;
        weights1[13190] <= 16'b1111111111110111;
        weights1[13191] <= 16'b0000000000000000;
        weights1[13192] <= 16'b0000000000001001;
        weights1[13193] <= 16'b1111111111100111;
        weights1[13194] <= 16'b1111111111111101;
        weights1[13195] <= 16'b0000000000001001;
        weights1[13196] <= 16'b1111111111110010;
        weights1[13197] <= 16'b1111111111111010;
        weights1[13198] <= 16'b0000000000000000;
        weights1[13199] <= 16'b0000000000010001;
        weights1[13200] <= 16'b0000000000010111;
        weights1[13201] <= 16'b0000000000000010;
        weights1[13202] <= 16'b1111111111101110;
        weights1[13203] <= 16'b1111111111100011;
        weights1[13204] <= 16'b0000000000000110;
        weights1[13205] <= 16'b1111111111100010;
        weights1[13206] <= 16'b1111111111110111;
        weights1[13207] <= 16'b1111111111110011;
        weights1[13208] <= 16'b1111111111100111;
        weights1[13209] <= 16'b1111111111110111;
        weights1[13210] <= 16'b1111111111111001;
        weights1[13211] <= 16'b0000000000001111;
        weights1[13212] <= 16'b1111111111111101;
        weights1[13213] <= 16'b1111111111111000;
        weights1[13214] <= 16'b1111111111101110;
        weights1[13215] <= 16'b1111111111111111;
        weights1[13216] <= 16'b1111111111111011;
        weights1[13217] <= 16'b1111111111111111;
        weights1[13218] <= 16'b0000000000000101;
        weights1[13219] <= 16'b1111111111111100;
        weights1[13220] <= 16'b0000000000000010;
        weights1[13221] <= 16'b0000000000001011;
        weights1[13222] <= 16'b1111111111101011;
        weights1[13223] <= 16'b1111111111101010;
        weights1[13224] <= 16'b1111111111100110;
        weights1[13225] <= 16'b1111111111110111;
        weights1[13226] <= 16'b1111111111110111;
        weights1[13227] <= 16'b1111111111110110;
        weights1[13228] <= 16'b1111111111111011;
        weights1[13229] <= 16'b0000000000011100;
        weights1[13230] <= 16'b1111111111111101;
        weights1[13231] <= 16'b0000000000000010;
        weights1[13232] <= 16'b0000000000011000;
        weights1[13233] <= 16'b1111111111101100;
        weights1[13234] <= 16'b0000000000001101;
        weights1[13235] <= 16'b1111111111111100;
        weights1[13236] <= 16'b1111111111111110;
        weights1[13237] <= 16'b1111111111110110;
        weights1[13238] <= 16'b1111111111101001;
        weights1[13239] <= 16'b1111111111111011;
        weights1[13240] <= 16'b1111111111110101;
        weights1[13241] <= 16'b1111111111111010;
        weights1[13242] <= 16'b1111111111111010;
        weights1[13243] <= 16'b0000000000000010;
        weights1[13244] <= 16'b1111111111111000;
        weights1[13245] <= 16'b1111111111111000;
        weights1[13246] <= 16'b1111111111111100;
        weights1[13247] <= 16'b0000000000000000;
        weights1[13248] <= 16'b0000000000000100;
        weights1[13249] <= 16'b1111111111111110;
        weights1[13250] <= 16'b0000000000000011;
        weights1[13251] <= 16'b0000000000001001;
        weights1[13252] <= 16'b0000000000000011;
        weights1[13253] <= 16'b0000000000001110;
        weights1[13254] <= 16'b0000000000000010;
        weights1[13255] <= 16'b0000000000000101;
        weights1[13256] <= 16'b0000000000000000;
        weights1[13257] <= 16'b1111111111101110;
        weights1[13258] <= 16'b1111111111111010;
        weights1[13259] <= 16'b0000000000100011;
        weights1[13260] <= 16'b1111111111111110;
        weights1[13261] <= 16'b1111111111111010;
        weights1[13262] <= 16'b0000000000000000;
        weights1[13263] <= 16'b1111111111110000;
        weights1[13264] <= 16'b1111111111111110;
        weights1[13265] <= 16'b1111111111110000;
        weights1[13266] <= 16'b1111111111110000;
        weights1[13267] <= 16'b1111111111101100;
        weights1[13268] <= 16'b1111111111101101;
        weights1[13269] <= 16'b1111111111111001;
        weights1[13270] <= 16'b1111111111111100;
        weights1[13271] <= 16'b0000000000000101;
        weights1[13272] <= 16'b1111111111111111;
        weights1[13273] <= 16'b1111111111111101;
        weights1[13274] <= 16'b1111111111111100;
        weights1[13275] <= 16'b1111111111111101;
        weights1[13276] <= 16'b0000000000000100;
        weights1[13277] <= 16'b1111111111111000;
        weights1[13278] <= 16'b1111111111110110;
        weights1[13279] <= 16'b0000000000000010;
        weights1[13280] <= 16'b1111111111111111;
        weights1[13281] <= 16'b1111111111111101;
        weights1[13282] <= 16'b1111111111110100;
        weights1[13283] <= 16'b1111111111101010;
        weights1[13284] <= 16'b1111111111110011;
        weights1[13285] <= 16'b1111111111101110;
        weights1[13286] <= 16'b1111111111111101;
        weights1[13287] <= 16'b1111111111110110;
        weights1[13288] <= 16'b1111111111100010;
        weights1[13289] <= 16'b1111111111110101;
        weights1[13290] <= 16'b1111111111101110;
        weights1[13291] <= 16'b1111111111111100;
        weights1[13292] <= 16'b1111111111111000;
        weights1[13293] <= 16'b1111111111111010;
        weights1[13294] <= 16'b1111111111110110;
        weights1[13295] <= 16'b1111111111110100;
        weights1[13296] <= 16'b1111111111111101;
        weights1[13297] <= 16'b1111111111111101;
        weights1[13298] <= 16'b1111111111111111;
        weights1[13299] <= 16'b0000000000000100;
        weights1[13300] <= 16'b1111111111111110;
        weights1[13301] <= 16'b1111111111111101;
        weights1[13302] <= 16'b1111111111111110;
        weights1[13303] <= 16'b0000000000000011;
        weights1[13304] <= 16'b0000000000000010;
        weights1[13305] <= 16'b1111111111111100;
        weights1[13306] <= 16'b0000000000001011;
        weights1[13307] <= 16'b0000000000001000;
        weights1[13308] <= 16'b0000000000001000;
        weights1[13309] <= 16'b1111111111111010;
        weights1[13310] <= 16'b1111111111110010;
        weights1[13311] <= 16'b1111111111111010;
        weights1[13312] <= 16'b0000000000000111;
        weights1[13313] <= 16'b1111111111111100;
        weights1[13314] <= 16'b1111111111111111;
        weights1[13315] <= 16'b0000000000001000;
        weights1[13316] <= 16'b1111111111110011;
        weights1[13317] <= 16'b1111111111101111;
        weights1[13318] <= 16'b1111111111111111;
        weights1[13319] <= 16'b0000000000000001;
        weights1[13320] <= 16'b1111111111111011;
        weights1[13321] <= 16'b1111111111110001;
        weights1[13322] <= 16'b1111111111111011;
        weights1[13323] <= 16'b1111111111110110;
        weights1[13324] <= 16'b1111111111110110;
        weights1[13325] <= 16'b1111111111111010;
        weights1[13326] <= 16'b1111111111111111;
        weights1[13327] <= 16'b0000000000000001;
        weights1[13328] <= 16'b0000000000000000;
        weights1[13329] <= 16'b0000000000000000;
        weights1[13330] <= 16'b1111111111111110;
        weights1[13331] <= 16'b0000000000000000;
        weights1[13332] <= 16'b1111111111111111;
        weights1[13333] <= 16'b1111111111111111;
        weights1[13334] <= 16'b1111111111111111;
        weights1[13335] <= 16'b0000000000000000;
        weights1[13336] <= 16'b0000000000000010;
        weights1[13337] <= 16'b0000000000000011;
        weights1[13338] <= 16'b1111111111111010;
        weights1[13339] <= 16'b1111111111111110;
        weights1[13340] <= 16'b0000000000000000;
        weights1[13341] <= 16'b1111111111110110;
        weights1[13342] <= 16'b0000000000000101;
        weights1[13343] <= 16'b1111111111110001;
        weights1[13344] <= 16'b1111111111110000;
        weights1[13345] <= 16'b1111111111101111;
        weights1[13346] <= 16'b1111111111110101;
        weights1[13347] <= 16'b1111111111111001;
        weights1[13348] <= 16'b1111111111110001;
        weights1[13349] <= 16'b1111111111101100;
        weights1[13350] <= 16'b1111111111110011;
        weights1[13351] <= 16'b1111111111111001;
        weights1[13352] <= 16'b1111111111111010;
        weights1[13353] <= 16'b0000000000000000;
        weights1[13354] <= 16'b0000000000000000;
        weights1[13355] <= 16'b0000000000000000;
        weights1[13356] <= 16'b0000000000000000;
        weights1[13357] <= 16'b1111111111111111;
        weights1[13358] <= 16'b1111111111111111;
        weights1[13359] <= 16'b1111111111111110;
        weights1[13360] <= 16'b1111111111111100;
        weights1[13361] <= 16'b1111111111111100;
        weights1[13362] <= 16'b1111111111111000;
        weights1[13363] <= 16'b1111111111111000;
        weights1[13364] <= 16'b1111111111110111;
        weights1[13365] <= 16'b0000000000000011;
        weights1[13366] <= 16'b0000000000000010;
        weights1[13367] <= 16'b0000000000000001;
        weights1[13368] <= 16'b0000000000001101;
        weights1[13369] <= 16'b0000000000000011;
        weights1[13370] <= 16'b0000000000010110;
        weights1[13371] <= 16'b1111111111110101;
        weights1[13372] <= 16'b1111111111100001;
        weights1[13373] <= 16'b1111111111111010;
        weights1[13374] <= 16'b0000000000001010;
        weights1[13375] <= 16'b1111111111110001;
        weights1[13376] <= 16'b1111111111111110;
        weights1[13377] <= 16'b1111111111110010;
        weights1[13378] <= 16'b1111111111111010;
        weights1[13379] <= 16'b1111111111111011;
        weights1[13380] <= 16'b1111111111110110;
        weights1[13381] <= 16'b1111111111110110;
        weights1[13382] <= 16'b1111111111111110;
        weights1[13383] <= 16'b1111111111111100;
        weights1[13384] <= 16'b1111111111111110;
        weights1[13385] <= 16'b1111111111111110;
        weights1[13386] <= 16'b1111111111111001;
        weights1[13387] <= 16'b1111111111111001;
        weights1[13388] <= 16'b1111111111110100;
        weights1[13389] <= 16'b1111111111110001;
        weights1[13390] <= 16'b1111111111110110;
        weights1[13391] <= 16'b1111111111101111;
        weights1[13392] <= 16'b1111111111110100;
        weights1[13393] <= 16'b1111111111111100;
        weights1[13394] <= 16'b1111111111111110;
        weights1[13395] <= 16'b0000000000001001;
        weights1[13396] <= 16'b0000000000010010;
        weights1[13397] <= 16'b0000000000011001;
        weights1[13398] <= 16'b0000000000001001;
        weights1[13399] <= 16'b0000000000000000;
        weights1[13400] <= 16'b1111111111100110;
        weights1[13401] <= 16'b1111111111100001;
        weights1[13402] <= 16'b0000000000000001;
        weights1[13403] <= 16'b1111111111111101;
        weights1[13404] <= 16'b1111111111110011;
        weights1[13405] <= 16'b1111111111111010;
        weights1[13406] <= 16'b0000000000001001;
        weights1[13407] <= 16'b1111111111111101;
        weights1[13408] <= 16'b1111111111111001;
        weights1[13409] <= 16'b1111111111111000;
        weights1[13410] <= 16'b1111111111111011;
        weights1[13411] <= 16'b1111111111111100;
        weights1[13412] <= 16'b1111111111111011;
        weights1[13413] <= 16'b1111111111111010;
        weights1[13414] <= 16'b1111111111110110;
        weights1[13415] <= 16'b1111111111101101;
        weights1[13416] <= 16'b1111111111101111;
        weights1[13417] <= 16'b1111111111101010;
        weights1[13418] <= 16'b1111111111100100;
        weights1[13419] <= 16'b1111111111011101;
        weights1[13420] <= 16'b1111111111101000;
        weights1[13421] <= 16'b1111111111100110;
        weights1[13422] <= 16'b1111111111100100;
        weights1[13423] <= 16'b0000000000001001;
        weights1[13424] <= 16'b0000000000001001;
        weights1[13425] <= 16'b1111111111101100;
        weights1[13426] <= 16'b1111111111111011;
        weights1[13427] <= 16'b1111111111111111;
        weights1[13428] <= 16'b1111111111101000;
        weights1[13429] <= 16'b1111111111101111;
        weights1[13430] <= 16'b1111111111111111;
        weights1[13431] <= 16'b0000000000000101;
        weights1[13432] <= 16'b0000000000001111;
        weights1[13433] <= 16'b1111111111111010;
        weights1[13434] <= 16'b1111111111111101;
        weights1[13435] <= 16'b1111111111110001;
        weights1[13436] <= 16'b0000000000000000;
        weights1[13437] <= 16'b1111111111111010;
        weights1[13438] <= 16'b1111111111111000;
        weights1[13439] <= 16'b1111111111111011;
        weights1[13440] <= 16'b1111111111111001;
        weights1[13441] <= 16'b1111111111110111;
        weights1[13442] <= 16'b1111111111110000;
        weights1[13443] <= 16'b1111111111110001;
        weights1[13444] <= 16'b1111111111100110;
        weights1[13445] <= 16'b1111111111100001;
        weights1[13446] <= 16'b1111111111011100;
        weights1[13447] <= 16'b1111111111010110;
        weights1[13448] <= 16'b1111111111011010;
        weights1[13449] <= 16'b1111111110111111;
        weights1[13450] <= 16'b1111111111011100;
        weights1[13451] <= 16'b1111111111101010;
        weights1[13452] <= 16'b0000000000000111;
        weights1[13453] <= 16'b0000000000010010;
        weights1[13454] <= 16'b0000000000010110;
        weights1[13455] <= 16'b0000000000000011;
        weights1[13456] <= 16'b1111111111100000;
        weights1[13457] <= 16'b1111111111110001;
        weights1[13458] <= 16'b1111111111100111;
        weights1[13459] <= 16'b1111111111111010;
        weights1[13460] <= 16'b1111111111110101;
        weights1[13461] <= 16'b0000000000001001;
        weights1[13462] <= 16'b0000000000000110;
        weights1[13463] <= 16'b0000000000000100;
        weights1[13464] <= 16'b0000000000000000;
        weights1[13465] <= 16'b1111111111111101;
        weights1[13466] <= 16'b1111111111111010;
        weights1[13467] <= 16'b1111111111111110;
        weights1[13468] <= 16'b1111111111110110;
        weights1[13469] <= 16'b1111111111110000;
        weights1[13470] <= 16'b1111111111101011;
        weights1[13471] <= 16'b1111111111100010;
        weights1[13472] <= 16'b1111111111001101;
        weights1[13473] <= 16'b1111111111001000;
        weights1[13474] <= 16'b1111111111010000;
        weights1[13475] <= 16'b1111111111000101;
        weights1[13476] <= 16'b1111111111000111;
        weights1[13477] <= 16'b1111111111011000;
        weights1[13478] <= 16'b1111111111000101;
        weights1[13479] <= 16'b1111111111000111;
        weights1[13480] <= 16'b1111111111111010;
        weights1[13481] <= 16'b0000000000000110;
        weights1[13482] <= 16'b0000000000010010;
        weights1[13483] <= 16'b0000000000001011;
        weights1[13484] <= 16'b0000000000001110;
        weights1[13485] <= 16'b1111111111111100;
        weights1[13486] <= 16'b1111111111101101;
        weights1[13487] <= 16'b1111111111110100;
        weights1[13488] <= 16'b1111111111101101;
        weights1[13489] <= 16'b1111111111110111;
        weights1[13490] <= 16'b1111111111110100;
        weights1[13491] <= 16'b0000000000000000;
        weights1[13492] <= 16'b1111111111111011;
        weights1[13493] <= 16'b1111111111110001;
        weights1[13494] <= 16'b1111111111110110;
        weights1[13495] <= 16'b1111111111111110;
        weights1[13496] <= 16'b1111111111111011;
        weights1[13497] <= 16'b1111111111110001;
        weights1[13498] <= 16'b1111111111101010;
        weights1[13499] <= 16'b1111111111011110;
        weights1[13500] <= 16'b1111111111001110;
        weights1[13501] <= 16'b1111111111011110;
        weights1[13502] <= 16'b1111111111000110;
        weights1[13503] <= 16'b1111111111010100;
        weights1[13504] <= 16'b0000000000000001;
        weights1[13505] <= 16'b1111111111110011;
        weights1[13506] <= 16'b1111111111011110;
        weights1[13507] <= 16'b1111111111100010;
        weights1[13508] <= 16'b0000000000001111;
        weights1[13509] <= 16'b0000000000001100;
        weights1[13510] <= 16'b0000000000000100;
        weights1[13511] <= 16'b1111111111111101;
        weights1[13512] <= 16'b1111111111111110;
        weights1[13513] <= 16'b0000000000000001;
        weights1[13514] <= 16'b1111111111100100;
        weights1[13515] <= 16'b1111111111110001;
        weights1[13516] <= 16'b1111111111111110;
        weights1[13517] <= 16'b0000000000001000;
        weights1[13518] <= 16'b1111111111111111;
        weights1[13519] <= 16'b0000000000001101;
        weights1[13520] <= 16'b0000000000000111;
        weights1[13521] <= 16'b1111111111111001;
        weights1[13522] <= 16'b1111111111111100;
        weights1[13523] <= 16'b1111111111111101;
        weights1[13524] <= 16'b1111111111111001;
        weights1[13525] <= 16'b1111111111110011;
        weights1[13526] <= 16'b1111111111111000;
        weights1[13527] <= 16'b1111111111110001;
        weights1[13528] <= 16'b1111111111101011;
        weights1[13529] <= 16'b1111111111110100;
        weights1[13530] <= 16'b1111111111110111;
        weights1[13531] <= 16'b0000000000000011;
        weights1[13532] <= 16'b1111111111101000;
        weights1[13533] <= 16'b0000000000000101;
        weights1[13534] <= 16'b1111111111111010;
        weights1[13535] <= 16'b1111111111001111;
        weights1[13536] <= 16'b1111111111011101;
        weights1[13537] <= 16'b0000000000000010;
        weights1[13538] <= 16'b1111111111111000;
        weights1[13539] <= 16'b1111111111110110;
        weights1[13540] <= 16'b0000000000000010;
        weights1[13541] <= 16'b1111111111111100;
        weights1[13542] <= 16'b1111111111110101;
        weights1[13543] <= 16'b0000000000000000;
        weights1[13544] <= 16'b1111111111101110;
        weights1[13545] <= 16'b0000000000000111;
        weights1[13546] <= 16'b1111111111100111;
        weights1[13547] <= 16'b0000000000000101;
        weights1[13548] <= 16'b1111111111011101;
        weights1[13549] <= 16'b1111111111111011;
        weights1[13550] <= 16'b1111111111101110;
        weights1[13551] <= 16'b1111111111111001;
        weights1[13552] <= 16'b0000000000000010;
        weights1[13553] <= 16'b0000000000000011;
        weights1[13554] <= 16'b1111111111111010;
        weights1[13555] <= 16'b0000000000000011;
        weights1[13556] <= 16'b0000000000000111;
        weights1[13557] <= 16'b0000000000011010;
        weights1[13558] <= 16'b0000000000000100;
        weights1[13559] <= 16'b1111111111110100;
        weights1[13560] <= 16'b1111111111110010;
        weights1[13561] <= 16'b0000000000001000;
        weights1[13562] <= 16'b0000000000010011;
        weights1[13563] <= 16'b1111111111011100;
        weights1[13564] <= 16'b1111111111110101;
        weights1[13565] <= 16'b0000000000000111;
        weights1[13566] <= 16'b0000000000000110;
        weights1[13567] <= 16'b0000000000001010;
        weights1[13568] <= 16'b1111111111110111;
        weights1[13569] <= 16'b1111111111111111;
        weights1[13570] <= 16'b1111111111111110;
        weights1[13571] <= 16'b1111111111110001;
        weights1[13572] <= 16'b1111111111111111;
        weights1[13573] <= 16'b1111111111110000;
        weights1[13574] <= 16'b1111111111110111;
        weights1[13575] <= 16'b0000000000001000;
        weights1[13576] <= 16'b1111111111111111;
        weights1[13577] <= 16'b1111111111111110;
        weights1[13578] <= 16'b1111111111110101;
        weights1[13579] <= 16'b1111111111101110;
        weights1[13580] <= 16'b0000000000001000;
        weights1[13581] <= 16'b0000000000001110;
        weights1[13582] <= 16'b0000000000001111;
        weights1[13583] <= 16'b1111111111110100;
        weights1[13584] <= 16'b0000000000101110;
        weights1[13585] <= 16'b0000000000001011;
        weights1[13586] <= 16'b0000000000000101;
        weights1[13587] <= 16'b0000000000001001;
        weights1[13588] <= 16'b1111111111111110;
        weights1[13589] <= 16'b0000000000001000;
        weights1[13590] <= 16'b0000000000010001;
        weights1[13591] <= 16'b1111111111101111;
        weights1[13592] <= 16'b1111111111110011;
        weights1[13593] <= 16'b0000000000000111;
        weights1[13594] <= 16'b0000000000100100;
        weights1[13595] <= 16'b0000000000000100;
        weights1[13596] <= 16'b1111111111111110;
        weights1[13597] <= 16'b1111111111101111;
        weights1[13598] <= 16'b1111111111111111;
        weights1[13599] <= 16'b1111111111111101;
        weights1[13600] <= 16'b1111111111111110;
        weights1[13601] <= 16'b1111111111110101;
        weights1[13602] <= 16'b0000000000000110;
        weights1[13603] <= 16'b1111111111111010;
        weights1[13604] <= 16'b1111111111100000;
        weights1[13605] <= 16'b1111111111111101;
        weights1[13606] <= 16'b1111111111111101;
        weights1[13607] <= 16'b1111111111110000;
        weights1[13608] <= 16'b0000000000001111;
        weights1[13609] <= 16'b0000000000001110;
        weights1[13610] <= 16'b0000000000010010;
        weights1[13611] <= 16'b0000000000000110;
        weights1[13612] <= 16'b0000000000000001;
        weights1[13613] <= 16'b0000000000011111;
        weights1[13614] <= 16'b0000000000010001;
        weights1[13615] <= 16'b0000000000001101;
        weights1[13616] <= 16'b0000000000011110;
        weights1[13617] <= 16'b1111111111111111;
        weights1[13618] <= 16'b0000000000010000;
        weights1[13619] <= 16'b0000000000000011;
        weights1[13620] <= 16'b1111111111101001;
        weights1[13621] <= 16'b0000000000010100;
        weights1[13622] <= 16'b0000000000001110;
        weights1[13623] <= 16'b1111111111101100;
        weights1[13624] <= 16'b1111111111110101;
        weights1[13625] <= 16'b1111111111101101;
        weights1[13626] <= 16'b1111111111101111;
        weights1[13627] <= 16'b1111111111111000;
        weights1[13628] <= 16'b1111111111101001;
        weights1[13629] <= 16'b0000000000000001;
        weights1[13630] <= 16'b1111111111100110;
        weights1[13631] <= 16'b1111111111111011;
        weights1[13632] <= 16'b1111111111111100;
        weights1[13633] <= 16'b0000000000001010;
        weights1[13634] <= 16'b1111111111110111;
        weights1[13635] <= 16'b1111111111110001;
        weights1[13636] <= 16'b0000000000010010;
        weights1[13637] <= 16'b0000000000010011;
        weights1[13638] <= 16'b0000000000000101;
        weights1[13639] <= 16'b0000000000000100;
        weights1[13640] <= 16'b1111111111111011;
        weights1[13641] <= 16'b0000000000000110;
        weights1[13642] <= 16'b0000000000000000;
        weights1[13643] <= 16'b1111111111110101;
        weights1[13644] <= 16'b0000000000001000;
        weights1[13645] <= 16'b0000000000000110;
        weights1[13646] <= 16'b0000000000011010;
        weights1[13647] <= 16'b0000000000011010;
        weights1[13648] <= 16'b1111111111111011;
        weights1[13649] <= 16'b1111111111110011;
        weights1[13650] <= 16'b1111111111101100;
        weights1[13651] <= 16'b1111111111101110;
        weights1[13652] <= 16'b1111111111100010;
        weights1[13653] <= 16'b1111111111110011;
        weights1[13654] <= 16'b1111111111111010;
        weights1[13655] <= 16'b1111111111111110;
        weights1[13656] <= 16'b1111111111111010;
        weights1[13657] <= 16'b1111111111111010;
        weights1[13658] <= 16'b1111111111110111;
        weights1[13659] <= 16'b1111111111101110;
        weights1[13660] <= 16'b1111111111101111;
        weights1[13661] <= 16'b1111111111111101;
        weights1[13662] <= 16'b1111111111110010;
        weights1[13663] <= 16'b1111111111100010;
        weights1[13664] <= 16'b0000000000001100;
        weights1[13665] <= 16'b0000000000010011;
        weights1[13666] <= 16'b0000000000000110;
        weights1[13667] <= 16'b1111111111111011;
        weights1[13668] <= 16'b1111111111111101;
        weights1[13669] <= 16'b0000000000011001;
        weights1[13670] <= 16'b0000000000010000;
        weights1[13671] <= 16'b0000000000001001;
        weights1[13672] <= 16'b0000000000001100;
        weights1[13673] <= 16'b0000000000011010;
        weights1[13674] <= 16'b0000000000011011;
        weights1[13675] <= 16'b0000000000001110;
        weights1[13676] <= 16'b1111111111100111;
        weights1[13677] <= 16'b1111111110111011;
        weights1[13678] <= 16'b1111111111100101;
        weights1[13679] <= 16'b1111111111011110;
        weights1[13680] <= 16'b1111111111100111;
        weights1[13681] <= 16'b1111111111101100;
        weights1[13682] <= 16'b1111111111110110;
        weights1[13683] <= 16'b1111111111101100;
        weights1[13684] <= 16'b1111111111110111;
        weights1[13685] <= 16'b1111111111100110;
        weights1[13686] <= 16'b1111111111100100;
        weights1[13687] <= 16'b1111111111110100;
        weights1[13688] <= 16'b1111111111110011;
        weights1[13689] <= 16'b1111111111011010;
        weights1[13690] <= 16'b1111111111100011;
        weights1[13691] <= 16'b1111111111100011;
        weights1[13692] <= 16'b0000000000001000;
        weights1[13693] <= 16'b0000000000001011;
        weights1[13694] <= 16'b0000000000000000;
        weights1[13695] <= 16'b1111111111111001;
        weights1[13696] <= 16'b1111111111111111;
        weights1[13697] <= 16'b0000000000000111;
        weights1[13698] <= 16'b0000000000000110;
        weights1[13699] <= 16'b0000000000011101;
        weights1[13700] <= 16'b0000000000001100;
        weights1[13701] <= 16'b0000000000100000;
        weights1[13702] <= 16'b0000000000010000;
        weights1[13703] <= 16'b0000000000000110;
        weights1[13704] <= 16'b1111111110100001;
        weights1[13705] <= 16'b1111111111100101;
        weights1[13706] <= 16'b1111111111001111;
        weights1[13707] <= 16'b1111111111011001;
        weights1[13708] <= 16'b1111111111110100;
        weights1[13709] <= 16'b1111111111101011;
        weights1[13710] <= 16'b1111111111111010;
        weights1[13711] <= 16'b1111111111110010;
        weights1[13712] <= 16'b1111111111111100;
        weights1[13713] <= 16'b1111111111111010;
        weights1[13714] <= 16'b1111111111110111;
        weights1[13715] <= 16'b1111111111101000;
        weights1[13716] <= 16'b1111111111100010;
        weights1[13717] <= 16'b1111111111100101;
        weights1[13718] <= 16'b1111111111011001;
        weights1[13719] <= 16'b1111111111100111;
        weights1[13720] <= 16'b0000000000000111;
        weights1[13721] <= 16'b0000000000001101;
        weights1[13722] <= 16'b0000000000000101;
        weights1[13723] <= 16'b0000000000001101;
        weights1[13724] <= 16'b1111111111111000;
        weights1[13725] <= 16'b0000000000010010;
        weights1[13726] <= 16'b0000000000001011;
        weights1[13727] <= 16'b0000000000100001;
        weights1[13728] <= 16'b0000000000011011;
        weights1[13729] <= 16'b0000000000001001;
        weights1[13730] <= 16'b0000000000001000;
        weights1[13731] <= 16'b1111111110101101;
        weights1[13732] <= 16'b1111111101101101;
        weights1[13733] <= 16'b1111111111000111;
        weights1[13734] <= 16'b1111111111010010;
        weights1[13735] <= 16'b1111111111101101;
        weights1[13736] <= 16'b1111111111110010;
        weights1[13737] <= 16'b1111111111111010;
        weights1[13738] <= 16'b1111111111110010;
        weights1[13739] <= 16'b0000000000000010;
        weights1[13740] <= 16'b1111111111111010;
        weights1[13741] <= 16'b1111111111101111;
        weights1[13742] <= 16'b1111111111100100;
        weights1[13743] <= 16'b1111111111100110;
        weights1[13744] <= 16'b1111111111011110;
        weights1[13745] <= 16'b1111111111101101;
        weights1[13746] <= 16'b1111111111110101;
        weights1[13747] <= 16'b1111111111111000;
        weights1[13748] <= 16'b0000000000000011;
        weights1[13749] <= 16'b0000000000010000;
        weights1[13750] <= 16'b0000000000001110;
        weights1[13751] <= 16'b0000000000100111;
        weights1[13752] <= 16'b1111111111111010;
        weights1[13753] <= 16'b0000000000101100;
        weights1[13754] <= 16'b0000000000100001;
        weights1[13755] <= 16'b0000000000000000;
        weights1[13756] <= 16'b0000000000101101;
        weights1[13757] <= 16'b1111111111111111;
        weights1[13758] <= 16'b1111111110011011;
        weights1[13759] <= 16'b1111111101000000;
        weights1[13760] <= 16'b1111111110000101;
        weights1[13761] <= 16'b1111111111100111;
        weights1[13762] <= 16'b1111111111100101;
        weights1[13763] <= 16'b0000000000000000;
        weights1[13764] <= 16'b1111111111100101;
        weights1[13765] <= 16'b1111111111110100;
        weights1[13766] <= 16'b1111111111111011;
        weights1[13767] <= 16'b1111111111110011;
        weights1[13768] <= 16'b1111111111111110;
        weights1[13769] <= 16'b1111111111101110;
        weights1[13770] <= 16'b0000000000000001;
        weights1[13771] <= 16'b1111111111110000;
        weights1[13772] <= 16'b0000000000001011;
        weights1[13773] <= 16'b1111111111101001;
        weights1[13774] <= 16'b1111111111101100;
        weights1[13775] <= 16'b1111111111111000;
        weights1[13776] <= 16'b0000000000000000;
        weights1[13777] <= 16'b0000000000000111;
        weights1[13778] <= 16'b0000000000010001;
        weights1[13779] <= 16'b0000000000010110;
        weights1[13780] <= 16'b0000000000100000;
        weights1[13781] <= 16'b0000000000010101;
        weights1[13782] <= 16'b0000000000001110;
        weights1[13783] <= 16'b0000000000011100;
        weights1[13784] <= 16'b1111111111101011;
        weights1[13785] <= 16'b1111111110101001;
        weights1[13786] <= 16'b1111111100010000;
        weights1[13787] <= 16'b1111111101011111;
        weights1[13788] <= 16'b1111111111100010;
        weights1[13789] <= 16'b1111111111111110;
        weights1[13790] <= 16'b0000000000000001;
        weights1[13791] <= 16'b0000000000010110;
        weights1[13792] <= 16'b1111111111111011;
        weights1[13793] <= 16'b0000000000001100;
        weights1[13794] <= 16'b0000000000001010;
        weights1[13795] <= 16'b0000000000000100;
        weights1[13796] <= 16'b0000000000000111;
        weights1[13797] <= 16'b0000000000100011;
        weights1[13798] <= 16'b0000000000000010;
        weights1[13799] <= 16'b0000000000001100;
        weights1[13800] <= 16'b1111111111110011;
        weights1[13801] <= 16'b1111111111111000;
        weights1[13802] <= 16'b1111111111110111;
        weights1[13803] <= 16'b0000000000010100;
        weights1[13804] <= 16'b1111111111110000;
        weights1[13805] <= 16'b0000000000001001;
        weights1[13806] <= 16'b1111111111101111;
        weights1[13807] <= 16'b1111111111110000;
        weights1[13808] <= 16'b0000000000011011;
        weights1[13809] <= 16'b0000000000000100;
        weights1[13810] <= 16'b1111111111011101;
        weights1[13811] <= 16'b1111111111001111;
        weights1[13812] <= 16'b1111111101111010;
        weights1[13813] <= 16'b1111111100101001;
        weights1[13814] <= 16'b1111111101001110;
        weights1[13815] <= 16'b1111111111001100;
        weights1[13816] <= 16'b0000000000001101;
        weights1[13817] <= 16'b0000000000001001;
        weights1[13818] <= 16'b1111111111111101;
        weights1[13819] <= 16'b1111111111110001;
        weights1[13820] <= 16'b0000000000000010;
        weights1[13821] <= 16'b0000000000000110;
        weights1[13822] <= 16'b0000000000011001;
        weights1[13823] <= 16'b0000000000000100;
        weights1[13824] <= 16'b1111111111101110;
        weights1[13825] <= 16'b1111111111110000;
        weights1[13826] <= 16'b1111111111111110;
        weights1[13827] <= 16'b1111111111111100;
        weights1[13828] <= 16'b0000000000000000;
        weights1[13829] <= 16'b0000000000011111;
        weights1[13830] <= 16'b0000000000011111;
        weights1[13831] <= 16'b0000000000011010;
        weights1[13832] <= 16'b1111111111101110;
        weights1[13833] <= 16'b1111111111110101;
        weights1[13834] <= 16'b1111111111101100;
        weights1[13835] <= 16'b1111111111010000;
        weights1[13836] <= 16'b1111111111100000;
        weights1[13837] <= 16'b1111111111011011;
        weights1[13838] <= 16'b1111111110110000;
        weights1[13839] <= 16'b1111111110001010;
        weights1[13840] <= 16'b1111111100101101;
        weights1[13841] <= 16'b1111111101010101;
        weights1[13842] <= 16'b1111111111010101;
        weights1[13843] <= 16'b0000000000000011;
        weights1[13844] <= 16'b0000000000001100;
        weights1[13845] <= 16'b0000000000010001;
        weights1[13846] <= 16'b0000000000011101;
        weights1[13847] <= 16'b0000000000010100;
        weights1[13848] <= 16'b1111111111111001;
        weights1[13849] <= 16'b0000000000010111;
        weights1[13850] <= 16'b0000000000001000;
        weights1[13851] <= 16'b0000000000010101;
        weights1[13852] <= 16'b0000000000001100;
        weights1[13853] <= 16'b0000000000000111;
        weights1[13854] <= 16'b0000000000010111;
        weights1[13855] <= 16'b1111111111111110;
        weights1[13856] <= 16'b0000000000000000;
        weights1[13857] <= 16'b0000000000100001;
        weights1[13858] <= 16'b0000000000011001;
        weights1[13859] <= 16'b0000000000101101;
        weights1[13860] <= 16'b1111111111100101;
        weights1[13861] <= 16'b1111111111101001;
        weights1[13862] <= 16'b1111111111010101;
        weights1[13863] <= 16'b1111111111010100;
        weights1[13864] <= 16'b1111111111001010;
        weights1[13865] <= 16'b1111111110101010;
        weights1[13866] <= 16'b1111111110000010;
        weights1[13867] <= 16'b1111111101010101;
        weights1[13868] <= 16'b1111111101101011;
        weights1[13869] <= 16'b1111111111001000;
        weights1[13870] <= 16'b1111111111111111;
        weights1[13871] <= 16'b1111111111110101;
        weights1[13872] <= 16'b1111111111111000;
        weights1[13873] <= 16'b0000000000000110;
        weights1[13874] <= 16'b1111111111111001;
        weights1[13875] <= 16'b0000000000001011;
        weights1[13876] <= 16'b0000000000000000;
        weights1[13877] <= 16'b0000000000001000;
        weights1[13878] <= 16'b0000000000001010;
        weights1[13879] <= 16'b0000000000001000;
        weights1[13880] <= 16'b0000000000011000;
        weights1[13881] <= 16'b0000000000000111;
        weights1[13882] <= 16'b1111111111111001;
        weights1[13883] <= 16'b0000000000010100;
        weights1[13884] <= 16'b0000000000100001;
        weights1[13885] <= 16'b0000000000001001;
        weights1[13886] <= 16'b0000000000011111;
        weights1[13887] <= 16'b0000000000101011;
        weights1[13888] <= 16'b1111111111011011;
        weights1[13889] <= 16'b1111111111010100;
        weights1[13890] <= 16'b1111111111000001;
        weights1[13891] <= 16'b1111111110111111;
        weights1[13892] <= 16'b1111111110100010;
        weights1[13893] <= 16'b1111111101111011;
        weights1[13894] <= 16'b1111111101110000;
        weights1[13895] <= 16'b1111111110001110;
        weights1[13896] <= 16'b1111111111011100;
        weights1[13897] <= 16'b0000000000000101;
        weights1[13898] <= 16'b0000000000001010;
        weights1[13899] <= 16'b0000000000001111;
        weights1[13900] <= 16'b0000000000010101;
        weights1[13901] <= 16'b0000000000000010;
        weights1[13902] <= 16'b0000000000010100;
        weights1[13903] <= 16'b0000000000010110;
        weights1[13904] <= 16'b0000000000000010;
        weights1[13905] <= 16'b0000000000000100;
        weights1[13906] <= 16'b0000000000001000;
        weights1[13907] <= 16'b1111111111111101;
        weights1[13908] <= 16'b0000000000001010;
        weights1[13909] <= 16'b0000000000001010;
        weights1[13910] <= 16'b0000000000000100;
        weights1[13911] <= 16'b0000000000001001;
        weights1[13912] <= 16'b0000000000011010;
        weights1[13913] <= 16'b0000000000000111;
        weights1[13914] <= 16'b0000000000010011;
        weights1[13915] <= 16'b0000000000011011;
        weights1[13916] <= 16'b1111111111011111;
        weights1[13917] <= 16'b1111111111010010;
        weights1[13918] <= 16'b1111111111000000;
        weights1[13919] <= 16'b1111111110110011;
        weights1[13920] <= 16'b1111111110010100;
        weights1[13921] <= 16'b1111111110010010;
        weights1[13922] <= 16'b1111111110100110;
        weights1[13923] <= 16'b1111111111011101;
        weights1[13924] <= 16'b0000000000001010;
        weights1[13925] <= 16'b0000000000010100;
        weights1[13926] <= 16'b0000000000001101;
        weights1[13927] <= 16'b0000000000010110;
        weights1[13928] <= 16'b0000000000001110;
        weights1[13929] <= 16'b0000000000011000;
        weights1[13930] <= 16'b0000000000001000;
        weights1[13931] <= 16'b0000000000010110;
        weights1[13932] <= 16'b0000000000010110;
        weights1[13933] <= 16'b0000000000010011;
        weights1[13934] <= 16'b0000000000000001;
        weights1[13935] <= 16'b0000000000000100;
        weights1[13936] <= 16'b0000000000000101;
        weights1[13937] <= 16'b0000000000000001;
        weights1[13938] <= 16'b0000000000010011;
        weights1[13939] <= 16'b0000000000011000;
        weights1[13940] <= 16'b0000000000001110;
        weights1[13941] <= 16'b0000000000011011;
        weights1[13942] <= 16'b0000000000011011;
        weights1[13943] <= 16'b0000000000101101;
        weights1[13944] <= 16'b1111111111010110;
        weights1[13945] <= 16'b1111111111001110;
        weights1[13946] <= 16'b1111111111001101;
        weights1[13947] <= 16'b1111111110111010;
        weights1[13948] <= 16'b1111111110011100;
        weights1[13949] <= 16'b1111111110110001;
        weights1[13950] <= 16'b1111111111101100;
        weights1[13951] <= 16'b0000000000100010;
        weights1[13952] <= 16'b0000000000010111;
        weights1[13953] <= 16'b0000000000011011;
        weights1[13954] <= 16'b0000000000001011;
        weights1[13955] <= 16'b0000000000001111;
        weights1[13956] <= 16'b0000000000011011;
        weights1[13957] <= 16'b0000000000001111;
        weights1[13958] <= 16'b0000000000011011;
        weights1[13959] <= 16'b0000000000010000;
        weights1[13960] <= 16'b1111111111110101;
        weights1[13961] <= 16'b0000000000000101;
        weights1[13962] <= 16'b1111111111110100;
        weights1[13963] <= 16'b1111111111110001;
        weights1[13964] <= 16'b1111111111111011;
        weights1[13965] <= 16'b0000000000001010;
        weights1[13966] <= 16'b0000000000001110;
        weights1[13967] <= 16'b0000000000011101;
        weights1[13968] <= 16'b0000000000011010;
        weights1[13969] <= 16'b0000000000001111;
        weights1[13970] <= 16'b0000000000001110;
        weights1[13971] <= 16'b0000000000011001;
        weights1[13972] <= 16'b1111111111011100;
        weights1[13973] <= 16'b1111111111001010;
        weights1[13974] <= 16'b1111111111001010;
        weights1[13975] <= 16'b1111111111001010;
        weights1[13976] <= 16'b1111111111010001;
        weights1[13977] <= 16'b1111111111111110;
        weights1[13978] <= 16'b0000000000000111;
        weights1[13979] <= 16'b0000000000011110;
        weights1[13980] <= 16'b1111111111111000;
        weights1[13981] <= 16'b0000000000001011;
        weights1[13982] <= 16'b0000000000011101;
        weights1[13983] <= 16'b0000000000010001;
        weights1[13984] <= 16'b0000000000001000;
        weights1[13985] <= 16'b0000000000000100;
        weights1[13986] <= 16'b0000000000001110;
        weights1[13987] <= 16'b0000000000010111;
        weights1[13988] <= 16'b0000000000001001;
        weights1[13989] <= 16'b0000000000001101;
        weights1[13990] <= 16'b0000000000000011;
        weights1[13991] <= 16'b0000000000001101;
        weights1[13992] <= 16'b0000000000000000;
        weights1[13993] <= 16'b0000000000010111;
        weights1[13994] <= 16'b1111111111111110;
        weights1[13995] <= 16'b0000000000001101;
        weights1[13996] <= 16'b0000000000100011;
        weights1[13997] <= 16'b0000000000010110;
        weights1[13998] <= 16'b0000000000010100;
        weights1[13999] <= 16'b0000000000010110;
        weights1[14000] <= 16'b1111111111100110;
        weights1[14001] <= 16'b1111111111011010;
        weights1[14002] <= 16'b1111111111000011;
        weights1[14003] <= 16'b1111111111011011;
        weights1[14004] <= 16'b1111111111100110;
        weights1[14005] <= 16'b1111111111110001;
        weights1[14006] <= 16'b0000000000101001;
        weights1[14007] <= 16'b0000000000010011;
        weights1[14008] <= 16'b0000000000000110;
        weights1[14009] <= 16'b0000000000010001;
        weights1[14010] <= 16'b1111111111111100;
        weights1[14011] <= 16'b0000000000000110;
        weights1[14012] <= 16'b1111111111110011;
        weights1[14013] <= 16'b1111111111111111;
        weights1[14014] <= 16'b0000000000001100;
        weights1[14015] <= 16'b1111111111110111;
        weights1[14016] <= 16'b1111111111111110;
        weights1[14017] <= 16'b0000000000010010;
        weights1[14018] <= 16'b0000000000010000;
        weights1[14019] <= 16'b0000000000000101;
        weights1[14020] <= 16'b0000000000000110;
        weights1[14021] <= 16'b1111111111111100;
        weights1[14022] <= 16'b0000000000001011;
        weights1[14023] <= 16'b0000000000010010;
        weights1[14024] <= 16'b0000000000010111;
        weights1[14025] <= 16'b0000000000001011;
        weights1[14026] <= 16'b0000000000001100;
        weights1[14027] <= 16'b0000000000010011;
        weights1[14028] <= 16'b1111111111110101;
        weights1[14029] <= 16'b1111111111100110;
        weights1[14030] <= 16'b1111111111011111;
        weights1[14031] <= 16'b1111111111100101;
        weights1[14032] <= 16'b1111111111100111;
        weights1[14033] <= 16'b1111111111111111;
        weights1[14034] <= 16'b0000000000001111;
        weights1[14035] <= 16'b0000000000001010;
        weights1[14036] <= 16'b0000000000001110;
        weights1[14037] <= 16'b0000000000011110;
        weights1[14038] <= 16'b0000000000000001;
        weights1[14039] <= 16'b0000000000011101;
        weights1[14040] <= 16'b0000000000010101;
        weights1[14041] <= 16'b1111111111111101;
        weights1[14042] <= 16'b1111111111111011;
        weights1[14043] <= 16'b1111111111110101;
        weights1[14044] <= 16'b1111111111111111;
        weights1[14045] <= 16'b0000000000000011;
        weights1[14046] <= 16'b0000000000001101;
        weights1[14047] <= 16'b0000000000001010;
        weights1[14048] <= 16'b1111111111111010;
        weights1[14049] <= 16'b0000000000010101;
        weights1[14050] <= 16'b0000000000000000;
        weights1[14051] <= 16'b1111111111111101;
        weights1[14052] <= 16'b0000000000001010;
        weights1[14053] <= 16'b0000000000001111;
        weights1[14054] <= 16'b0000000000000100;
        weights1[14055] <= 16'b0000000000000111;
        weights1[14056] <= 16'b1111111111111110;
        weights1[14057] <= 16'b1111111111111110;
        weights1[14058] <= 16'b1111111111110111;
        weights1[14059] <= 16'b0000000000000001;
        weights1[14060] <= 16'b0000000000010001;
        weights1[14061] <= 16'b1111111111111101;
        weights1[14062] <= 16'b0000000000001000;
        weights1[14063] <= 16'b0000000000001101;
        weights1[14064] <= 16'b0000000000100100;
        weights1[14065] <= 16'b0000000000001100;
        weights1[14066] <= 16'b1111111111111011;
        weights1[14067] <= 16'b0000000000010111;
        weights1[14068] <= 16'b0000000000000011;
        weights1[14069] <= 16'b0000000000001011;
        weights1[14070] <= 16'b1111111111111110;
        weights1[14071] <= 16'b0000000000000011;
        weights1[14072] <= 16'b0000000000001001;
        weights1[14073] <= 16'b0000000000000101;
        weights1[14074] <= 16'b0000000000000000;
        weights1[14075] <= 16'b0000000000001101;
        weights1[14076] <= 16'b0000000000000001;
        weights1[14077] <= 16'b0000000000001100;
        weights1[14078] <= 16'b1111111111111100;
        weights1[14079] <= 16'b0000000000000000;
        weights1[14080] <= 16'b0000000000000100;
        weights1[14081] <= 16'b0000000000000111;
        weights1[14082] <= 16'b0000000000001101;
        weights1[14083] <= 16'b0000000000000101;
        weights1[14084] <= 16'b1111111111111111;
        weights1[14085] <= 16'b0000000000000011;
        weights1[14086] <= 16'b0000000000001101;
        weights1[14087] <= 16'b0000000000010100;
        weights1[14088] <= 16'b0000000000001100;
        weights1[14089] <= 16'b0000000000001110;
        weights1[14090] <= 16'b0000000000010011;
        weights1[14091] <= 16'b0000000000010100;
        weights1[14092] <= 16'b0000000000010000;
        weights1[14093] <= 16'b0000000000010000;
        weights1[14094] <= 16'b0000000000101011;
        weights1[14095] <= 16'b0000000000001000;
        weights1[14096] <= 16'b0000000000000110;
        weights1[14097] <= 16'b1111111111111011;
        weights1[14098] <= 16'b0000000000000001;
        weights1[14099] <= 16'b1111111111110001;
        weights1[14100] <= 16'b1111111111110101;
        weights1[14101] <= 16'b1111111111111000;
        weights1[14102] <= 16'b0000000000000100;
        weights1[14103] <= 16'b1111111111110110;
        weights1[14104] <= 16'b0000000000000111;
        weights1[14105] <= 16'b0000000000000010;
        weights1[14106] <= 16'b1111111111110111;
        weights1[14107] <= 16'b0000000000001001;
        weights1[14108] <= 16'b1111111111111011;
        weights1[14109] <= 16'b1111111111111110;
        weights1[14110] <= 16'b0000000000000010;
        weights1[14111] <= 16'b0000000000000010;
        weights1[14112] <= 16'b0000000000000000;
        weights1[14113] <= 16'b0000000000000000;
        weights1[14114] <= 16'b0000000000000001;
        weights1[14115] <= 16'b0000000000000010;
        weights1[14116] <= 16'b1111111111111110;
        weights1[14117] <= 16'b0000000000000100;
        weights1[14118] <= 16'b0000000000000000;
        weights1[14119] <= 16'b1111111111111101;
        weights1[14120] <= 16'b0000000000001000;
        weights1[14121] <= 16'b1111111111111100;
        weights1[14122] <= 16'b1111111111111111;
        weights1[14123] <= 16'b0000000000010011;
        weights1[14124] <= 16'b0000000000010111;
        weights1[14125] <= 16'b0000000000001010;
        weights1[14126] <= 16'b0000000000001101;
        weights1[14127] <= 16'b0000000000000110;
        weights1[14128] <= 16'b1111111111110110;
        weights1[14129] <= 16'b1111111111111101;
        weights1[14130] <= 16'b1111111111101101;
        weights1[14131] <= 16'b0000000000001000;
        weights1[14132] <= 16'b0000000000001011;
        weights1[14133] <= 16'b0000000000000110;
        weights1[14134] <= 16'b0000000000000100;
        weights1[14135] <= 16'b1111111111110110;
        weights1[14136] <= 16'b1111111111111111;
        weights1[14137] <= 16'b0000000000000010;
        weights1[14138] <= 16'b0000000000000011;
        weights1[14139] <= 16'b1111111111111110;
        weights1[14140] <= 16'b0000000000000000;
        weights1[14141] <= 16'b0000000000000000;
        weights1[14142] <= 16'b0000000000000001;
        weights1[14143] <= 16'b0000000000000101;
        weights1[14144] <= 16'b0000000000000101;
        weights1[14145] <= 16'b0000000000000110;
        weights1[14146] <= 16'b0000000000000010;
        weights1[14147] <= 16'b1111111111110100;
        weights1[14148] <= 16'b0000000000000101;
        weights1[14149] <= 16'b1111111111110011;
        weights1[14150] <= 16'b1111111111110111;
        weights1[14151] <= 16'b1111111111111110;
        weights1[14152] <= 16'b0000000000000011;
        weights1[14153] <= 16'b0000000000000101;
        weights1[14154] <= 16'b1111111111110010;
        weights1[14155] <= 16'b0000000000001011;
        weights1[14156] <= 16'b0000000000001010;
        weights1[14157] <= 16'b0000000000001011;
        weights1[14158] <= 16'b0000000000000110;
        weights1[14159] <= 16'b1111111111111000;
        weights1[14160] <= 16'b1111111111111010;
        weights1[14161] <= 16'b1111111111111111;
        weights1[14162] <= 16'b0000000000000010;
        weights1[14163] <= 16'b1111111111111010;
        weights1[14164] <= 16'b1111111111111101;
        weights1[14165] <= 16'b1111111111111100;
        weights1[14166] <= 16'b1111111111110111;
        weights1[14167] <= 16'b1111111111111111;
        weights1[14168] <= 16'b1111111111111111;
        weights1[14169] <= 16'b0000000000000001;
        weights1[14170] <= 16'b0000000000000011;
        weights1[14171] <= 16'b0000000000001001;
        weights1[14172] <= 16'b0000000000001000;
        weights1[14173] <= 16'b0000000000000101;
        weights1[14174] <= 16'b0000000000001100;
        weights1[14175] <= 16'b1111111111101010;
        weights1[14176] <= 16'b0000000000000000;
        weights1[14177] <= 16'b1111111111101110;
        weights1[14178] <= 16'b1111111111100110;
        weights1[14179] <= 16'b1111111111011101;
        weights1[14180] <= 16'b1111111111011111;
        weights1[14181] <= 16'b1111111111111101;
        weights1[14182] <= 16'b0000000000000101;
        weights1[14183] <= 16'b1111111111110010;
        weights1[14184] <= 16'b1111111111111111;
        weights1[14185] <= 16'b0000000000000011;
        weights1[14186] <= 16'b0000000000000100;
        weights1[14187] <= 16'b0000000000001111;
        weights1[14188] <= 16'b0000000000000111;
        weights1[14189] <= 16'b0000000000000001;
        weights1[14190] <= 16'b0000000000001011;
        weights1[14191] <= 16'b1111111111111010;
        weights1[14192] <= 16'b0000000000001011;
        weights1[14193] <= 16'b0000000000000001;
        weights1[14194] <= 16'b0000000000000001;
        weights1[14195] <= 16'b1111111111111111;
        weights1[14196] <= 16'b0000000000000001;
        weights1[14197] <= 16'b0000000000000011;
        weights1[14198] <= 16'b0000000000000010;
        weights1[14199] <= 16'b0000000000000110;
        weights1[14200] <= 16'b1111111111111111;
        weights1[14201] <= 16'b0000000000010000;
        weights1[14202] <= 16'b0000000000001111;
        weights1[14203] <= 16'b0000000000011000;
        weights1[14204] <= 16'b0000000000011101;
        weights1[14205] <= 16'b0000000000000100;
        weights1[14206] <= 16'b0000000000001100;
        weights1[14207] <= 16'b1111111111111110;
        weights1[14208] <= 16'b0000000000000100;
        weights1[14209] <= 16'b0000000000000100;
        weights1[14210] <= 16'b0000000000001101;
        weights1[14211] <= 16'b0000000000001000;
        weights1[14212] <= 16'b0000000000000111;
        weights1[14213] <= 16'b0000000000001111;
        weights1[14214] <= 16'b1111111111101010;
        weights1[14215] <= 16'b0000000000000010;
        weights1[14216] <= 16'b0000000000000000;
        weights1[14217] <= 16'b0000000000010000;
        weights1[14218] <= 16'b1111111111111110;
        weights1[14219] <= 16'b1111111111110111;
        weights1[14220] <= 16'b0000000000000011;
        weights1[14221] <= 16'b1111111111110001;
        weights1[14222] <= 16'b1111111111111001;
        weights1[14223] <= 16'b0000000000000111;
        weights1[14224] <= 16'b0000000000001000;
        weights1[14225] <= 16'b0000000000001001;
        weights1[14226] <= 16'b0000000000000100;
        weights1[14227] <= 16'b1111111111111001;
        weights1[14228] <= 16'b0000000000011000;
        weights1[14229] <= 16'b0000000000100000;
        weights1[14230] <= 16'b0000000000010110;
        weights1[14231] <= 16'b0000000000100111;
        weights1[14232] <= 16'b0000000000010001;
        weights1[14233] <= 16'b0000000000101110;
        weights1[14234] <= 16'b0000000000100110;
        weights1[14235] <= 16'b0000000000011011;
        weights1[14236] <= 16'b0000000000011001;
        weights1[14237] <= 16'b0000000000000100;
        weights1[14238] <= 16'b1111111111101100;
        weights1[14239] <= 16'b1111111111101110;
        weights1[14240] <= 16'b1111111111101111;
        weights1[14241] <= 16'b1111111111110111;
        weights1[14242] <= 16'b0000000000010000;
        weights1[14243] <= 16'b1111111111111111;
        weights1[14244] <= 16'b1111111111111010;
        weights1[14245] <= 16'b1111111111101111;
        weights1[14246] <= 16'b0000000000001001;
        weights1[14247] <= 16'b0000000000000010;
        weights1[14248] <= 16'b0000000000001110;
        weights1[14249] <= 16'b1111111111110010;
        weights1[14250] <= 16'b0000000000000100;
        weights1[14251] <= 16'b1111111111111111;
        weights1[14252] <= 16'b0000000000001000;
        weights1[14253] <= 16'b0000000000001101;
        weights1[14254] <= 16'b0000000000000101;
        weights1[14255] <= 16'b0000000000100001;
        weights1[14256] <= 16'b0000000000110000;
        weights1[14257] <= 16'b0000000000100011;
        weights1[14258] <= 16'b0000000000010110;
        weights1[14259] <= 16'b0000000000010111;
        weights1[14260] <= 16'b0000000000010001;
        weights1[14261] <= 16'b0000000000010110;
        weights1[14262] <= 16'b1111111111111100;
        weights1[14263] <= 16'b1111111111101011;
        weights1[14264] <= 16'b0000000000000011;
        weights1[14265] <= 16'b1111111111111010;
        weights1[14266] <= 16'b0000000000001010;
        weights1[14267] <= 16'b1111111111111101;
        weights1[14268] <= 16'b0000000000010101;
        weights1[14269] <= 16'b0000000000001010;
        weights1[14270] <= 16'b1111111111110111;
        weights1[14271] <= 16'b1111111111110101;
        weights1[14272] <= 16'b0000000000001101;
        weights1[14273] <= 16'b1111111111111110;
        weights1[14274] <= 16'b0000000000010011;
        weights1[14275] <= 16'b1111111111111110;
        weights1[14276] <= 16'b1111111111110001;
        weights1[14277] <= 16'b1111111111111111;
        weights1[14278] <= 16'b1111111111110110;
        weights1[14279] <= 16'b1111111111110000;
        weights1[14280] <= 16'b0000000000000100;
        weights1[14281] <= 16'b0000000000001110;
        weights1[14282] <= 16'b0000000000011001;
        weights1[14283] <= 16'b0000000000101100;
        weights1[14284] <= 16'b0000000000111100;
        weights1[14285] <= 16'b0000000000010111;
        weights1[14286] <= 16'b0000000000010011;
        weights1[14287] <= 16'b0000000000011001;
        weights1[14288] <= 16'b0000000000001011;
        weights1[14289] <= 16'b0000000000011010;
        weights1[14290] <= 16'b0000000000011100;
        weights1[14291] <= 16'b0000000000010111;
        weights1[14292] <= 16'b0000000000011000;
        weights1[14293] <= 16'b1111111111110101;
        weights1[14294] <= 16'b0000000000100111;
        weights1[14295] <= 16'b1111111111111101;
        weights1[14296] <= 16'b0000000000000101;
        weights1[14297] <= 16'b1111111111110011;
        weights1[14298] <= 16'b0000000000010001;
        weights1[14299] <= 16'b0000000000010000;
        weights1[14300] <= 16'b1111111111111110;
        weights1[14301] <= 16'b1111111111101110;
        weights1[14302] <= 16'b0000000000010000;
        weights1[14303] <= 16'b0000000000000110;
        weights1[14304] <= 16'b1111111111101000;
        weights1[14305] <= 16'b1111111111111110;
        weights1[14306] <= 16'b1111111111111111;
        weights1[14307] <= 16'b1111111111111100;
        weights1[14308] <= 16'b0000000000000100;
        weights1[14309] <= 16'b0000000000010101;
        weights1[14310] <= 16'b0000000000100101;
        weights1[14311] <= 16'b0000000000111000;
        weights1[14312] <= 16'b0000000001000001;
        weights1[14313] <= 16'b0000000000110111;
        weights1[14314] <= 16'b0000000001100111;
        weights1[14315] <= 16'b0000000000110010;
        weights1[14316] <= 16'b0000000000100101;
        weights1[14317] <= 16'b0000000000110000;
        weights1[14318] <= 16'b0000000000111001;
        weights1[14319] <= 16'b0000000000110000;
        weights1[14320] <= 16'b0000000000010001;
        weights1[14321] <= 16'b0000000000100110;
        weights1[14322] <= 16'b0000000000010010;
        weights1[14323] <= 16'b0000000000010001;
        weights1[14324] <= 16'b0000000000001111;
        weights1[14325] <= 16'b0000000000010110;
        weights1[14326] <= 16'b0000000000000110;
        weights1[14327] <= 16'b1111111111111111;
        weights1[14328] <= 16'b0000000000000111;
        weights1[14329] <= 16'b0000000000000111;
        weights1[14330] <= 16'b0000000000000111;
        weights1[14331] <= 16'b1111111111101110;
        weights1[14332] <= 16'b0000000000001100;
        weights1[14333] <= 16'b1111111111110011;
        weights1[14334] <= 16'b0000000000000010;
        weights1[14335] <= 16'b0000000000000000;
        weights1[14336] <= 16'b0000000000000111;
        weights1[14337] <= 16'b0000000000001010;
        weights1[14338] <= 16'b0000000000010111;
        weights1[14339] <= 16'b0000000000101111;
        weights1[14340] <= 16'b0000000001001111;
        weights1[14341] <= 16'b0000000000110111;
        weights1[14342] <= 16'b0000000001010110;
        weights1[14343] <= 16'b0000000001000000;
        weights1[14344] <= 16'b0000000001011111;
        weights1[14345] <= 16'b0000000000111011;
        weights1[14346] <= 16'b0000000001000001;
        weights1[14347] <= 16'b0000000001000001;
        weights1[14348] <= 16'b0000000000101100;
        weights1[14349] <= 16'b0000000000110010;
        weights1[14350] <= 16'b0000000000100110;
        weights1[14351] <= 16'b0000000000010111;
        weights1[14352] <= 16'b0000000000001101;
        weights1[14353] <= 16'b0000000000011010;
        weights1[14354] <= 16'b0000000000001111;
        weights1[14355] <= 16'b0000000000001000;
        weights1[14356] <= 16'b0000000000010110;
        weights1[14357] <= 16'b0000000000000101;
        weights1[14358] <= 16'b0000000000000100;
        weights1[14359] <= 16'b1111111111101001;
        weights1[14360] <= 16'b0000000000001011;
        weights1[14361] <= 16'b0000000000001010;
        weights1[14362] <= 16'b0000000000000101;
        weights1[14363] <= 16'b0000000000001010;
        weights1[14364] <= 16'b0000000000000000;
        weights1[14365] <= 16'b1111111111101111;
        weights1[14366] <= 16'b1111111111111001;
        weights1[14367] <= 16'b0000000000001001;
        weights1[14368] <= 16'b0000000000011011;
        weights1[14369] <= 16'b0000000000001110;
        weights1[14370] <= 16'b0000000000010011;
        weights1[14371] <= 16'b0000000000100001;
        weights1[14372] <= 16'b0000000000110111;
        weights1[14373] <= 16'b0000000000001111;
        weights1[14374] <= 16'b0000000000011011;
        weights1[14375] <= 16'b0000000000101111;
        weights1[14376] <= 16'b0000000000100100;
        weights1[14377] <= 16'b0000000000010000;
        weights1[14378] <= 16'b0000000000001010;
        weights1[14379] <= 16'b0000000000010001;
        weights1[14380] <= 16'b0000000000000001;
        weights1[14381] <= 16'b1111111111110111;
        weights1[14382] <= 16'b0000000000000101;
        weights1[14383] <= 16'b0000000000000010;
        weights1[14384] <= 16'b1111111111111001;
        weights1[14385] <= 16'b0000000000010000;
        weights1[14386] <= 16'b0000000000010010;
        weights1[14387] <= 16'b1111111111111100;
        weights1[14388] <= 16'b0000000000000010;
        weights1[14389] <= 16'b0000000000000110;
        weights1[14390] <= 16'b0000000000001110;
        weights1[14391] <= 16'b0000000000001001;
        weights1[14392] <= 16'b1111111111101011;
        weights1[14393] <= 16'b1111111111001001;
        weights1[14394] <= 16'b1111111110111011;
        weights1[14395] <= 16'b1111111110111000;
        weights1[14396] <= 16'b1111111110101100;
        weights1[14397] <= 16'b1111111110111100;
        weights1[14398] <= 16'b1111111111000010;
        weights1[14399] <= 16'b1111111110111001;
        weights1[14400] <= 16'b1111111110111001;
        weights1[14401] <= 16'b1111111111001001;
        weights1[14402] <= 16'b1111111110111010;
        weights1[14403] <= 16'b1111111110011100;
        weights1[14404] <= 16'b1111111110111100;
        weights1[14405] <= 16'b1111111110110111;
        weights1[14406] <= 16'b1111111110111000;
        weights1[14407] <= 16'b1111111110111100;
        weights1[14408] <= 16'b1111111111110000;
        weights1[14409] <= 16'b1111111111110001;
        weights1[14410] <= 16'b1111111111101101;
        weights1[14411] <= 16'b1111111111110100;
        weights1[14412] <= 16'b1111111111111111;
        weights1[14413] <= 16'b1111111111110110;
        weights1[14414] <= 16'b1111111111110001;
        weights1[14415] <= 16'b0000000000000111;
        weights1[14416] <= 16'b1111111111101100;
        weights1[14417] <= 16'b0000000000010011;
        weights1[14418] <= 16'b1111111111111111;
        weights1[14419] <= 16'b0000000000010000;
        weights1[14420] <= 16'b1111111111000010;
        weights1[14421] <= 16'b1111111110010101;
        weights1[14422] <= 16'b1111111110000110;
        weights1[14423] <= 16'b1111111101111011;
        weights1[14424] <= 16'b1111111101010001;
        weights1[14425] <= 16'b1111111101001000;
        weights1[14426] <= 16'b1111111101001000;
        weights1[14427] <= 16'b1111111100110110;
        weights1[14428] <= 16'b1111111100000011;
        weights1[14429] <= 16'b1111111100001101;
        weights1[14430] <= 16'b1111111100101111;
        weights1[14431] <= 16'b1111111101100001;
        weights1[14432] <= 16'b1111111101111110;
        weights1[14433] <= 16'b1111111110011101;
        weights1[14434] <= 16'b1111111111010001;
        weights1[14435] <= 16'b1111111111001101;
        weights1[14436] <= 16'b1111111111100011;
        weights1[14437] <= 16'b1111111111110010;
        weights1[14438] <= 16'b1111111111100101;
        weights1[14439] <= 16'b1111111111110101;
        weights1[14440] <= 16'b1111111111111011;
        weights1[14441] <= 16'b1111111111100111;
        weights1[14442] <= 16'b1111111111111101;
        weights1[14443] <= 16'b1111111111111110;
        weights1[14444] <= 16'b0000000000000100;
        weights1[14445] <= 16'b0000000000001010;
        weights1[14446] <= 16'b0000000000000100;
        weights1[14447] <= 16'b1111111111110110;
        weights1[14448] <= 16'b1111111110110100;
        weights1[14449] <= 16'b1111111110001011;
        weights1[14450] <= 16'b1111111101110001;
        weights1[14451] <= 16'b1111111101001100;
        weights1[14452] <= 16'b1111111100110000;
        weights1[14453] <= 16'b1111111100001000;
        weights1[14454] <= 16'b1111111011101101;
        weights1[14455] <= 16'b1111111011010010;
        weights1[14456] <= 16'b1111111100000101;
        weights1[14457] <= 16'b1111111101100000;
        weights1[14458] <= 16'b1111111110101001;
        weights1[14459] <= 16'b1111111111000000;
        weights1[14460] <= 16'b1111111111100101;
        weights1[14461] <= 16'b1111111111101100;
        weights1[14462] <= 16'b1111111111111011;
        weights1[14463] <= 16'b1111111111111010;
        weights1[14464] <= 16'b0000000000001110;
        weights1[14465] <= 16'b1111111111110101;
        weights1[14466] <= 16'b0000000000001101;
        weights1[14467] <= 16'b1111111111111110;
        weights1[14468] <= 16'b0000000000001011;
        weights1[14469] <= 16'b0000000000000100;
        weights1[14470] <= 16'b0000000000000011;
        weights1[14471] <= 16'b0000000000000010;
        weights1[14472] <= 16'b1111111111111000;
        weights1[14473] <= 16'b0000000000001101;
        weights1[14474] <= 16'b1111111111110110;
        weights1[14475] <= 16'b1111111111111011;
        weights1[14476] <= 16'b1111111110110000;
        weights1[14477] <= 16'b1111111110010001;
        weights1[14478] <= 16'b1111111110000000;
        weights1[14479] <= 16'b1111111101101001;
        weights1[14480] <= 16'b1111111101011001;
        weights1[14481] <= 16'b1111111101110011;
        weights1[14482] <= 16'b1111111110001010;
        weights1[14483] <= 16'b1111111111001001;
        weights1[14484] <= 16'b0000000000001001;
        weights1[14485] <= 16'b0000000000001101;
        weights1[14486] <= 16'b0000000000011000;
        weights1[14487] <= 16'b0000000000011001;
        weights1[14488] <= 16'b0000000000010100;
        weights1[14489] <= 16'b0000000000010001;
        weights1[14490] <= 16'b0000000000001011;
        weights1[14491] <= 16'b0000000000000110;
        weights1[14492] <= 16'b0000000000001110;
        weights1[14493] <= 16'b1111111111110011;
        weights1[14494] <= 16'b1111111111111100;
        weights1[14495] <= 16'b0000000000000000;
        weights1[14496] <= 16'b1111111111110110;
        weights1[14497] <= 16'b0000000000011001;
        weights1[14498] <= 16'b0000000000000101;
        weights1[14499] <= 16'b0000000000000011;
        weights1[14500] <= 16'b1111111111111010;
        weights1[14501] <= 16'b0000000000001100;
        weights1[14502] <= 16'b1111111111111111;
        weights1[14503] <= 16'b0000000000000011;
        weights1[14504] <= 16'b1111111111000111;
        weights1[14505] <= 16'b1111111110101011;
        weights1[14506] <= 16'b1111111110110011;
        weights1[14507] <= 16'b1111111110111111;
        weights1[14508] <= 16'b1111111111011100;
        weights1[14509] <= 16'b0000000000010011;
        weights1[14510] <= 16'b0000000001000000;
        weights1[14511] <= 16'b0000000001001110;
        weights1[14512] <= 16'b0000000000111000;
        weights1[14513] <= 16'b0000000000111001;
        weights1[14514] <= 16'b0000000000101010;
        weights1[14515] <= 16'b0000000000100110;
        weights1[14516] <= 16'b0000000000011100;
        weights1[14517] <= 16'b0000000000001011;
        weights1[14518] <= 16'b0000000000011010;
        weights1[14519] <= 16'b0000000000000011;
        weights1[14520] <= 16'b0000000000000100;
        weights1[14521] <= 16'b0000000000000011;
        weights1[14522] <= 16'b0000000000001000;
        weights1[14523] <= 16'b0000000000000110;
        weights1[14524] <= 16'b0000000000001001;
        weights1[14525] <= 16'b1111111111111111;
        weights1[14526] <= 16'b0000000000000110;
        weights1[14527] <= 16'b0000000000000011;
        weights1[14528] <= 16'b1111111111111000;
        weights1[14529] <= 16'b1111111111111100;
        weights1[14530] <= 16'b1111111111110111;
        weights1[14531] <= 16'b1111111111111010;
        weights1[14532] <= 16'b1111111111011000;
        weights1[14533] <= 16'b1111111111010111;
        weights1[14534] <= 16'b1111111111100101;
        weights1[14535] <= 16'b1111111111110110;
        weights1[14536] <= 16'b0000000000100001;
        weights1[14537] <= 16'b0000000000111101;
        weights1[14538] <= 16'b0000000000111011;
        weights1[14539] <= 16'b0000000000111111;
        weights1[14540] <= 16'b0000000000100000;
        weights1[14541] <= 16'b0000000000010010;
        weights1[14542] <= 16'b0000000000001001;
        weights1[14543] <= 16'b0000000000011111;
        weights1[14544] <= 16'b0000000000000010;
        weights1[14545] <= 16'b1111111111111111;
        weights1[14546] <= 16'b1111111111111000;
        weights1[14547] <= 16'b0000000000001011;
        weights1[14548] <= 16'b0000000000010010;
        weights1[14549] <= 16'b0000000000001100;
        weights1[14550] <= 16'b0000000000000000;
        weights1[14551] <= 16'b0000000000000100;
        weights1[14552] <= 16'b1111111111110010;
        weights1[14553] <= 16'b1111111111110101;
        weights1[14554] <= 16'b0000000000000001;
        weights1[14555] <= 16'b0000000000000000;
        weights1[14556] <= 16'b0000000000000000;
        weights1[14557] <= 16'b0000000000000010;
        weights1[14558] <= 16'b0000000000000110;
        weights1[14559] <= 16'b0000000000010011;
        weights1[14560] <= 16'b1111111111110110;
        weights1[14561] <= 16'b0000000000000010;
        weights1[14562] <= 16'b0000000000010010;
        weights1[14563] <= 16'b0000000000011010;
        weights1[14564] <= 16'b0000000000111111;
        weights1[14565] <= 16'b0000000000000100;
        weights1[14566] <= 16'b0000000000100100;
        weights1[14567] <= 16'b0000000000011101;
        weights1[14568] <= 16'b0000000000010001;
        weights1[14569] <= 16'b0000000000001100;
        weights1[14570] <= 16'b0000000000000001;
        weights1[14571] <= 16'b1111111111110100;
        weights1[14572] <= 16'b0000000000000100;
        weights1[14573] <= 16'b1111111111111011;
        weights1[14574] <= 16'b0000000000000101;
        weights1[14575] <= 16'b1111111111110111;
        weights1[14576] <= 16'b0000000000000010;
        weights1[14577] <= 16'b1111111111110100;
        weights1[14578] <= 16'b0000000000001010;
        weights1[14579] <= 16'b0000000000001100;
        weights1[14580] <= 16'b0000000000010000;
        weights1[14581] <= 16'b1111111111111101;
        weights1[14582] <= 16'b0000000000001000;
        weights1[14583] <= 16'b0000000000001001;
        weights1[14584] <= 16'b0000000000001100;
        weights1[14585] <= 16'b0000000000010101;
        weights1[14586] <= 16'b0000000000010111;
        weights1[14587] <= 16'b0000000000001000;
        weights1[14588] <= 16'b0000000000001101;
        weights1[14589] <= 16'b0000000000100000;
        weights1[14590] <= 16'b0000000000010011;
        weights1[14591] <= 16'b1111111111111111;
        weights1[14592] <= 16'b0000000000010011;
        weights1[14593] <= 16'b1111111111111101;
        weights1[14594] <= 16'b1111111111110000;
        weights1[14595] <= 16'b1111111111111100;
        weights1[14596] <= 16'b1111111111101111;
        weights1[14597] <= 16'b0000000000000000;
        weights1[14598] <= 16'b1111111111111100;
        weights1[14599] <= 16'b0000000000001101;
        weights1[14600] <= 16'b1111111111110101;
        weights1[14601] <= 16'b0000000000000011;
        weights1[14602] <= 16'b0000000000000001;
        weights1[14603] <= 16'b1111111111110110;
        weights1[14604] <= 16'b0000000000000101;
        weights1[14605] <= 16'b1111111111110111;
        weights1[14606] <= 16'b1111111111111101;
        weights1[14607] <= 16'b1111111111110101;
        weights1[14608] <= 16'b0000000000000111;
        weights1[14609] <= 16'b0000000000001011;
        weights1[14610] <= 16'b0000000000000101;
        weights1[14611] <= 16'b0000000000000110;
        weights1[14612] <= 16'b1111111111111100;
        weights1[14613] <= 16'b0000000000000011;
        weights1[14614] <= 16'b0000000000000000;
        weights1[14615] <= 16'b1111111111111110;
        weights1[14616] <= 16'b0000000000100100;
        weights1[14617] <= 16'b0000000000010000;
        weights1[14618] <= 16'b0000000000011000;
        weights1[14619] <= 16'b0000000000001011;
        weights1[14620] <= 16'b0000000000010111;
        weights1[14621] <= 16'b0000000000000101;
        weights1[14622] <= 16'b0000000000011011;
        weights1[14623] <= 16'b0000000000011110;
        weights1[14624] <= 16'b0000000000000011;
        weights1[14625] <= 16'b0000000000010110;
        weights1[14626] <= 16'b0000000000000001;
        weights1[14627] <= 16'b1111111111110011;
        weights1[14628] <= 16'b0000000000000011;
        weights1[14629] <= 16'b1111111111111010;
        weights1[14630] <= 16'b1111111111111100;
        weights1[14631] <= 16'b1111111111111000;
        weights1[14632] <= 16'b1111111111110011;
        weights1[14633] <= 16'b1111111111110111;
        weights1[14634] <= 16'b1111111111110110;
        weights1[14635] <= 16'b1111111111111111;
        weights1[14636] <= 16'b1111111111111001;
        weights1[14637] <= 16'b1111111111101101;
        weights1[14638] <= 16'b1111111111101010;
        weights1[14639] <= 16'b0000000000000000;
        weights1[14640] <= 16'b1111111111110111;
        weights1[14641] <= 16'b0000000000000110;
        weights1[14642] <= 16'b0000000000000011;
        weights1[14643] <= 16'b1111111111111111;
        weights1[14644] <= 16'b0000000000010110;
        weights1[14645] <= 16'b0000000000001011;
        weights1[14646] <= 16'b0000000000001110;
        weights1[14647] <= 16'b1111111111111110;
        weights1[14648] <= 16'b0000000000000011;
        weights1[14649] <= 16'b1111111111101101;
        weights1[14650] <= 16'b1111111111101110;
        weights1[14651] <= 16'b0000000000001001;
        weights1[14652] <= 16'b1111111111110001;
        weights1[14653] <= 16'b1111111111110001;
        weights1[14654] <= 16'b1111111111111001;
        weights1[14655] <= 16'b0000000000001011;
        weights1[14656] <= 16'b1111111111101111;
        weights1[14657] <= 16'b0000000000001010;
        weights1[14658] <= 16'b0000000000001101;
        weights1[14659] <= 16'b1111111111111101;
        weights1[14660] <= 16'b0000000000001001;
        weights1[14661] <= 16'b1111111111111110;
        weights1[14662] <= 16'b1111111111111000;
        weights1[14663] <= 16'b0000000000000001;
        weights1[14664] <= 16'b1111111111111111;
        weights1[14665] <= 16'b1111111111111110;
        weights1[14666] <= 16'b0000000000000111;
        weights1[14667] <= 16'b0000000000000001;
        weights1[14668] <= 16'b1111111111111010;
        weights1[14669] <= 16'b1111111111110110;
        weights1[14670] <= 16'b1111111111111111;
        weights1[14671] <= 16'b0000000000000001;
        weights1[14672] <= 16'b0000000000001001;
        weights1[14673] <= 16'b0000000000010100;
        weights1[14674] <= 16'b1111111111111001;
        weights1[14675] <= 16'b0000000000010001;
        weights1[14676] <= 16'b0000000000001010;
        weights1[14677] <= 16'b0000000000001111;
        weights1[14678] <= 16'b0000000000001100;
        weights1[14679] <= 16'b1111111111111101;
        weights1[14680] <= 16'b1111111111111110;
        weights1[14681] <= 16'b0000000000001000;
        weights1[14682] <= 16'b0000000000000000;
        weights1[14683] <= 16'b0000000000001010;
        weights1[14684] <= 16'b1111111111111101;
        weights1[14685] <= 16'b1111111111110100;
        weights1[14686] <= 16'b1111111111111100;
        weights1[14687] <= 16'b1111111111110110;
        weights1[14688] <= 16'b0000000000001001;
        weights1[14689] <= 16'b1111111111111111;
        weights1[14690] <= 16'b1111111111110100;
        weights1[14691] <= 16'b1111111111111000;
        weights1[14692] <= 16'b1111111111111000;
        weights1[14693] <= 16'b1111111111101000;
        weights1[14694] <= 16'b1111111111101010;
        weights1[14695] <= 16'b1111111111101001;
        weights1[14696] <= 16'b1111111111101110;
        weights1[14697] <= 16'b1111111111110010;
        weights1[14698] <= 16'b1111111111110011;
        weights1[14699] <= 16'b1111111111111000;
        weights1[14700] <= 16'b0000000000000001;
        weights1[14701] <= 16'b1111111111111010;
        weights1[14702] <= 16'b1111111111110110;
        weights1[14703] <= 16'b0000000000001000;
        weights1[14704] <= 16'b0000000000000011;
        weights1[14705] <= 16'b1111111111110101;
        weights1[14706] <= 16'b1111111111110000;
        weights1[14707] <= 16'b1111111111111111;
        weights1[14708] <= 16'b0000000000010011;
        weights1[14709] <= 16'b0000000000001110;
        weights1[14710] <= 16'b0000000000010100;
        weights1[14711] <= 16'b0000000000001101;
        weights1[14712] <= 16'b0000000000001010;
        weights1[14713] <= 16'b0000000000001001;
        weights1[14714] <= 16'b0000000000000100;
        weights1[14715] <= 16'b1111111111110101;
        weights1[14716] <= 16'b1111111111110100;
        weights1[14717] <= 16'b1111111111111010;
        weights1[14718] <= 16'b1111111111111111;
        weights1[14719] <= 16'b0000000000000011;
        weights1[14720] <= 16'b0000000000010101;
        weights1[14721] <= 16'b0000000000000010;
        weights1[14722] <= 16'b1111111111110011;
        weights1[14723] <= 16'b0000000000001100;
        weights1[14724] <= 16'b1111111111111001;
        weights1[14725] <= 16'b1111111111110101;
        weights1[14726] <= 16'b1111111111101110;
        weights1[14727] <= 16'b0000000000000001;
        weights1[14728] <= 16'b1111111111111001;
        weights1[14729] <= 16'b1111111111101111;
        weights1[14730] <= 16'b1111111111101110;
        weights1[14731] <= 16'b1111111111111011;
        weights1[14732] <= 16'b1111111111110100;
        weights1[14733] <= 16'b0000000000000011;
        weights1[14734] <= 16'b1111111111111101;
        weights1[14735] <= 16'b0000000000000010;
        weights1[14736] <= 16'b1111111111111101;
        weights1[14737] <= 16'b1111111111101001;
        weights1[14738] <= 16'b1111111111110000;
        weights1[14739] <= 16'b1111111111110100;
        weights1[14740] <= 16'b1111111111111110;
        weights1[14741] <= 16'b0000000000000000;
        weights1[14742] <= 16'b1111111111110100;
        weights1[14743] <= 16'b0000000000000111;
        weights1[14744] <= 16'b0000000000000011;
        weights1[14745] <= 16'b1111111111111001;
        weights1[14746] <= 16'b1111111111111100;
        weights1[14747] <= 16'b0000000000001110;
        weights1[14748] <= 16'b0000000000000011;
        weights1[14749] <= 16'b0000000000000011;
        weights1[14750] <= 16'b0000000000000100;
        weights1[14751] <= 16'b1111111111111100;
        weights1[14752] <= 16'b0000000000001001;
        weights1[14753] <= 16'b0000000000001000;
        weights1[14754] <= 16'b1111111111110101;
        weights1[14755] <= 16'b1111111111111110;
        weights1[14756] <= 16'b1111111111110101;
        weights1[14757] <= 16'b1111111111101111;
        weights1[14758] <= 16'b1111111111110001;
        weights1[14759] <= 16'b1111111111101110;
        weights1[14760] <= 16'b1111111111111011;
        weights1[14761] <= 16'b1111111111111001;
        weights1[14762] <= 16'b0000000000000010;
        weights1[14763] <= 16'b1111111111111010;
        weights1[14764] <= 16'b0000000000001010;
        weights1[14765] <= 16'b0000000000001111;
        weights1[14766] <= 16'b1111111111110101;
        weights1[14767] <= 16'b0000000000000100;
        weights1[14768] <= 16'b1111111111111000;
        weights1[14769] <= 16'b1111111111110110;
        weights1[14770] <= 16'b0000000000001100;
        weights1[14771] <= 16'b0000000000000001;
        weights1[14772] <= 16'b1111111111110111;
        weights1[14773] <= 16'b1111111111110010;
        weights1[14774] <= 16'b1111111111101100;
        weights1[14775] <= 16'b1111111111110101;
        weights1[14776] <= 16'b1111111111111010;
        weights1[14777] <= 16'b0000000000001110;
        weights1[14778] <= 16'b1111111111111110;
        weights1[14779] <= 16'b1111111111110011;
        weights1[14780] <= 16'b0000000000000101;
        weights1[14781] <= 16'b1111111111111111;
        weights1[14782] <= 16'b1111111111111100;
        weights1[14783] <= 16'b0000000000000101;
        weights1[14784] <= 16'b1111111111111001;
        weights1[14785] <= 16'b1111111111101011;
        weights1[14786] <= 16'b1111111111110011;
        weights1[14787] <= 16'b1111111111111010;
        weights1[14788] <= 16'b0000000000000000;
        weights1[14789] <= 16'b0000000000001010;
        weights1[14790] <= 16'b1111111111110110;
        weights1[14791] <= 16'b1111111111110111;
        weights1[14792] <= 16'b1111111111110101;
        weights1[14793] <= 16'b1111111111110100;
        weights1[14794] <= 16'b0000000000000100;
        weights1[14795] <= 16'b0000000000001110;
        weights1[14796] <= 16'b1111111111110101;
        weights1[14797] <= 16'b0000000000000001;
        weights1[14798] <= 16'b1111111111101010;
        weights1[14799] <= 16'b0000000000001100;
        weights1[14800] <= 16'b1111111111111000;
        weights1[14801] <= 16'b0000000000000000;
        weights1[14802] <= 16'b0000000000000010;
        weights1[14803] <= 16'b1111111111110110;
        weights1[14804] <= 16'b0000000000001001;
        weights1[14805] <= 16'b0000000000000011;
        weights1[14806] <= 16'b0000000000010010;
        weights1[14807] <= 16'b1111111111111100;
        weights1[14808] <= 16'b0000000000000010;
        weights1[14809] <= 16'b0000000000000100;
        weights1[14810] <= 16'b0000000000000110;
        weights1[14811] <= 16'b0000000000000011;
        weights1[14812] <= 16'b1111111111111110;
        weights1[14813] <= 16'b1111111111101101;
        weights1[14814] <= 16'b1111111111110011;
        weights1[14815] <= 16'b1111111111111001;
        weights1[14816] <= 16'b1111111111111101;
        weights1[14817] <= 16'b0000000000000100;
        weights1[14818] <= 16'b1111111111111101;
        weights1[14819] <= 16'b1111111111111011;
        weights1[14820] <= 16'b1111111111111101;
        weights1[14821] <= 16'b0000000000010101;
        weights1[14822] <= 16'b1111111111111100;
        weights1[14823] <= 16'b1111111111110111;
        weights1[14824] <= 16'b0000000000001011;
        weights1[14825] <= 16'b1111111111111011;
        weights1[14826] <= 16'b0000000000001000;
        weights1[14827] <= 16'b0000000000000101;
        weights1[14828] <= 16'b1111111111111111;
        weights1[14829] <= 16'b0000000000010000;
        weights1[14830] <= 16'b1111111111110001;
        weights1[14831] <= 16'b1111111111110101;
        weights1[14832] <= 16'b1111111111111110;
        weights1[14833] <= 16'b1111111111110111;
        weights1[14834] <= 16'b0000000000001111;
        weights1[14835] <= 16'b0000000000001000;
        weights1[14836] <= 16'b0000000000010001;
        weights1[14837] <= 16'b0000000000001001;
        weights1[14838] <= 16'b0000000000001001;
        weights1[14839] <= 16'b0000000000000001;
        weights1[14840] <= 16'b0000000000000000;
        weights1[14841] <= 16'b0000000000000010;
        weights1[14842] <= 16'b1111111111110101;
        weights1[14843] <= 16'b1111111111110001;
        weights1[14844] <= 16'b1111111111110010;
        weights1[14845] <= 16'b1111111111101110;
        weights1[14846] <= 16'b1111111111110001;
        weights1[14847] <= 16'b1111111111110111;
        weights1[14848] <= 16'b1111111111110010;
        weights1[14849] <= 16'b1111111111101110;
        weights1[14850] <= 16'b1111111111110110;
        weights1[14851] <= 16'b1111111111111000;
        weights1[14852] <= 16'b1111111111110110;
        weights1[14853] <= 16'b1111111111111010;
        weights1[14854] <= 16'b1111111111101101;
        weights1[14855] <= 16'b1111111111110100;
        weights1[14856] <= 16'b0000000000000001;
        weights1[14857] <= 16'b0000000000000010;
        weights1[14858] <= 16'b0000000000000110;
        weights1[14859] <= 16'b0000000000001011;
        weights1[14860] <= 16'b0000000000000100;
        weights1[14861] <= 16'b0000000000001001;
        weights1[14862] <= 16'b1111111111111101;
        weights1[14863] <= 16'b0000000000000001;
        weights1[14864] <= 16'b0000000000000110;
        weights1[14865] <= 16'b0000000000000110;
        weights1[14866] <= 16'b0000000000000100;
        weights1[14867] <= 16'b0000000000000000;
        weights1[14868] <= 16'b1111111111111110;
        weights1[14869] <= 16'b0000000000000000;
        weights1[14870] <= 16'b1111111111111001;
        weights1[14871] <= 16'b1111111111110111;
        weights1[14872] <= 16'b1111111111111001;
        weights1[14873] <= 16'b0000000000000100;
        weights1[14874] <= 16'b1111111111111100;
        weights1[14875] <= 16'b1111111111110001;
        weights1[14876] <= 16'b1111111111110110;
        weights1[14877] <= 16'b0000000000000110;
        weights1[14878] <= 16'b0000000000001100;
        weights1[14879] <= 16'b0000000000000111;
        weights1[14880] <= 16'b0000000000000001;
        weights1[14881] <= 16'b1111111111110110;
        weights1[14882] <= 16'b1111111111111100;
        weights1[14883] <= 16'b0000000000001010;
        weights1[14884] <= 16'b0000000000001101;
        weights1[14885] <= 16'b0000000000001001;
        weights1[14886] <= 16'b0000000000001001;
        weights1[14887] <= 16'b0000000000000111;
        weights1[14888] <= 16'b0000000000001000;
        weights1[14889] <= 16'b0000000000000111;
        weights1[14890] <= 16'b1111111111111011;
        weights1[14891] <= 16'b0000000000000110;
        weights1[14892] <= 16'b0000000000001010;
        weights1[14893] <= 16'b0000000000001011;
        weights1[14894] <= 16'b0000000000000010;
        weights1[14895] <= 16'b1111111111111111;
        weights1[14896] <= 16'b0000000000000000;
        weights1[14897] <= 16'b0000000000000000;
        weights1[14898] <= 16'b1111111111111111;
        weights1[14899] <= 16'b1111111111111111;
        weights1[14900] <= 16'b0000000000000000;
        weights1[14901] <= 16'b1111111111111101;
        weights1[14902] <= 16'b1111111111111100;
        weights1[14903] <= 16'b1111111111111110;
        weights1[14904] <= 16'b0000000000000010;
        weights1[14905] <= 16'b0000000000000001;
        weights1[14906] <= 16'b0000000000000111;
        weights1[14907] <= 16'b0000000000011101;
        weights1[14908] <= 16'b0000000000110001;
        weights1[14909] <= 16'b0000000000011101;
        weights1[14910] <= 16'b0000000000100001;
        weights1[14911] <= 16'b0000000000011011;
        weights1[14912] <= 16'b0000000000000110;
        weights1[14913] <= 16'b0000000000010010;
        weights1[14914] <= 16'b0000000000000101;
        weights1[14915] <= 16'b1111111111111001;
        weights1[14916] <= 16'b1111111111110000;
        weights1[14917] <= 16'b1111111111110101;
        weights1[14918] <= 16'b1111111111110010;
        weights1[14919] <= 16'b1111111111101101;
        weights1[14920] <= 16'b1111111111111000;
        weights1[14921] <= 16'b1111111111111100;
        weights1[14922] <= 16'b1111111111111010;
        weights1[14923] <= 16'b1111111111111101;
        weights1[14924] <= 16'b0000000000000000;
        weights1[14925] <= 16'b1111111111111111;
        weights1[14926] <= 16'b1111111111111101;
        weights1[14927] <= 16'b1111111111111110;
        weights1[14928] <= 16'b1111111111111011;
        weights1[14929] <= 16'b1111111111101111;
        weights1[14930] <= 16'b1111111111100111;
        weights1[14931] <= 16'b1111111111100110;
        weights1[14932] <= 16'b1111111111101001;
        weights1[14933] <= 16'b1111111111110101;
        weights1[14934] <= 16'b0000000000001011;
        weights1[14935] <= 16'b0000000000011111;
        weights1[14936] <= 16'b0000000000101011;
        weights1[14937] <= 16'b0000000000100111;
        weights1[14938] <= 16'b0000000000101111;
        weights1[14939] <= 16'b0000000000100011;
        weights1[14940] <= 16'b0000000000010010;
        weights1[14941] <= 16'b0000000000010111;
        weights1[14942] <= 16'b0000000000000101;
        weights1[14943] <= 16'b1111111111111101;
        weights1[14944] <= 16'b1111111111111101;
        weights1[14945] <= 16'b1111111111111010;
        weights1[14946] <= 16'b1111111111111000;
        weights1[14947] <= 16'b1111111111110110;
        weights1[14948] <= 16'b1111111111110001;
        weights1[14949] <= 16'b1111111111110010;
        weights1[14950] <= 16'b1111111111110111;
        weights1[14951] <= 16'b1111111111111011;
        weights1[14952] <= 16'b0000000000000000;
        weights1[14953] <= 16'b1111111111111111;
        weights1[14954] <= 16'b1111111111111010;
        weights1[14955] <= 16'b1111111111110100;
        weights1[14956] <= 16'b1111111111101001;
        weights1[14957] <= 16'b1111111111100010;
        weights1[14958] <= 16'b1111111111011010;
        weights1[14959] <= 16'b1111111111001110;
        weights1[14960] <= 16'b1111111111010000;
        weights1[14961] <= 16'b1111111111010101;
        weights1[14962] <= 16'b1111111111100000;
        weights1[14963] <= 16'b1111111111110011;
        weights1[14964] <= 16'b0000000000000100;
        weights1[14965] <= 16'b0000000000011101;
        weights1[14966] <= 16'b0000000000100111;
        weights1[14967] <= 16'b0000000000101001;
        weights1[14968] <= 16'b0000000000100110;
        weights1[14969] <= 16'b0000000000100001;
        weights1[14970] <= 16'b0000000000011111;
        weights1[14971] <= 16'b0000000000010000;
        weights1[14972] <= 16'b0000000000000011;
        weights1[14973] <= 16'b0000000000001011;
        weights1[14974] <= 16'b1111111111111100;
        weights1[14975] <= 16'b1111111111110000;
        weights1[14976] <= 16'b1111111111110100;
        weights1[14977] <= 16'b1111111111110001;
        weights1[14978] <= 16'b1111111111110101;
        weights1[14979] <= 16'b1111111111111001;
        weights1[14980] <= 16'b1111111111111101;
        weights1[14981] <= 16'b1111111111111101;
        weights1[14982] <= 16'b1111111111110110;
        weights1[14983] <= 16'b1111111111101000;
        weights1[14984] <= 16'b1111111111010111;
        weights1[14985] <= 16'b1111111111001001;
        weights1[14986] <= 16'b1111111111000000;
        weights1[14987] <= 16'b1111111110110010;
        weights1[14988] <= 16'b1111111111000101;
        weights1[14989] <= 16'b1111111110111000;
        weights1[14990] <= 16'b1111111111000001;
        weights1[14991] <= 16'b1111111111000101;
        weights1[14992] <= 16'b1111111111011000;
        weights1[14993] <= 16'b1111111111101000;
        weights1[14994] <= 16'b1111111111101000;
        weights1[14995] <= 16'b0000000000000010;
        weights1[14996] <= 16'b0000000000001010;
        weights1[14997] <= 16'b0000000000010110;
        weights1[14998] <= 16'b0000000000011001;
        weights1[14999] <= 16'b0000000000010011;
        weights1[15000] <= 16'b0000000000000110;
        weights1[15001] <= 16'b0000000000000110;
        weights1[15002] <= 16'b0000000000000111;
        weights1[15003] <= 16'b0000000000000001;
        weights1[15004] <= 16'b1111111111111100;
        weights1[15005] <= 16'b1111111111100110;
        weights1[15006] <= 16'b1111111111101001;
        weights1[15007] <= 16'b1111111111110110;
        weights1[15008] <= 16'b1111111111111110;
        weights1[15009] <= 16'b1111111111110110;
        weights1[15010] <= 16'b1111111111101001;
        weights1[15011] <= 16'b1111111111011110;
        weights1[15012] <= 16'b1111111111000111;
        weights1[15013] <= 16'b1111111110111011;
        weights1[15014] <= 16'b1111111110110000;
        weights1[15015] <= 16'b1111111110110001;
        weights1[15016] <= 16'b1111111110101100;
        weights1[15017] <= 16'b1111111110011001;
        weights1[15018] <= 16'b1111111110010110;
        weights1[15019] <= 16'b1111111110010010;
        weights1[15020] <= 16'b1111111110100000;
        weights1[15021] <= 16'b1111111110111111;
        weights1[15022] <= 16'b1111111111001001;
        weights1[15023] <= 16'b1111111111010011;
        weights1[15024] <= 16'b1111111111001010;
        weights1[15025] <= 16'b1111111111010111;
        weights1[15026] <= 16'b1111111111111000;
        weights1[15027] <= 16'b0000000000000010;
        weights1[15028] <= 16'b0000000000001000;
        weights1[15029] <= 16'b0000000000010001;
        weights1[15030] <= 16'b0000000000010101;
        weights1[15031] <= 16'b0000000000001100;
        weights1[15032] <= 16'b1111111111110011;
        weights1[15033] <= 16'b1111111111110000;
        weights1[15034] <= 16'b1111111111110010;
        weights1[15035] <= 16'b1111111111110101;
        weights1[15036] <= 16'b1111111111111100;
        weights1[15037] <= 16'b1111111111110101;
        weights1[15038] <= 16'b1111111111100111;
        weights1[15039] <= 16'b1111111111010001;
        weights1[15040] <= 16'b1111111110111111;
        weights1[15041] <= 16'b1111111111000010;
        weights1[15042] <= 16'b1111111111001101;
        weights1[15043] <= 16'b1111111110111011;
        weights1[15044] <= 16'b1111111110011111;
        weights1[15045] <= 16'b1111111110001101;
        weights1[15046] <= 16'b1111111101111001;
        weights1[15047] <= 16'b1111111110001011;
        weights1[15048] <= 16'b1111111101111111;
        weights1[15049] <= 16'b1111111110100010;
        weights1[15050] <= 16'b1111111111010010;
        weights1[15051] <= 16'b1111111111110101;
        weights1[15052] <= 16'b1111111111111011;
        weights1[15053] <= 16'b1111111111101110;
        weights1[15054] <= 16'b1111111111110111;
        weights1[15055] <= 16'b0000000000001000;
        weights1[15056] <= 16'b0000000000000000;
        weights1[15057] <= 16'b1111111111111010;
        weights1[15058] <= 16'b1111111111111101;
        weights1[15059] <= 16'b0000000000001011;
        weights1[15060] <= 16'b1111111111111010;
        weights1[15061] <= 16'b1111111111110011;
        weights1[15062] <= 16'b1111111111101000;
        weights1[15063] <= 16'b1111111111101100;
        weights1[15064] <= 16'b1111111111111100;
        weights1[15065] <= 16'b1111111111110100;
        weights1[15066] <= 16'b1111111111110000;
        weights1[15067] <= 16'b1111111111100000;
        weights1[15068] <= 16'b1111111111101110;
        weights1[15069] <= 16'b1111111111101110;
        weights1[15070] <= 16'b1111111111011010;
        weights1[15071] <= 16'b1111111111001000;
        weights1[15072] <= 16'b1111111111101010;
        weights1[15073] <= 16'b1111111111100101;
        weights1[15074] <= 16'b1111111111000010;
        weights1[15075] <= 16'b1111111111010111;
        weights1[15076] <= 16'b1111111111010000;
        weights1[15077] <= 16'b1111111111011010;
        weights1[15078] <= 16'b1111111111010101;
        weights1[15079] <= 16'b1111111111001111;
        weights1[15080] <= 16'b1111111111101110;
        weights1[15081] <= 16'b0000000000000000;
        weights1[15082] <= 16'b1111111111111000;
        weights1[15083] <= 16'b0000000000000110;
        weights1[15084] <= 16'b1111111111101010;
        weights1[15085] <= 16'b0000000000010110;
        weights1[15086] <= 16'b1111111111101110;
        weights1[15087] <= 16'b1111111111111011;
        weights1[15088] <= 16'b0000000000000101;
        weights1[15089] <= 16'b1111111111110101;
        weights1[15090] <= 16'b1111111111110100;
        weights1[15091] <= 16'b1111111111111000;
        weights1[15092] <= 16'b1111111111111110;
        weights1[15093] <= 16'b1111111111111111;
        weights1[15094] <= 16'b1111111111111100;
        weights1[15095] <= 16'b1111111111111000;
        weights1[15096] <= 16'b0000000000001100;
        weights1[15097] <= 16'b0000000000100100;
        weights1[15098] <= 16'b0000000000110011;
        weights1[15099] <= 16'b0000000000100000;
        weights1[15100] <= 16'b0000000000000010;
        weights1[15101] <= 16'b0000000000010111;
        weights1[15102] <= 16'b0000000000010111;
        weights1[15103] <= 16'b1111111111100100;
        weights1[15104] <= 16'b1111111111101100;
        weights1[15105] <= 16'b1111111111111110;
        weights1[15106] <= 16'b1111111111110011;
        weights1[15107] <= 16'b1111111111110001;
        weights1[15108] <= 16'b1111111111101001;
        weights1[15109] <= 16'b0000000000000011;
        weights1[15110] <= 16'b0000000000000110;
        weights1[15111] <= 16'b1111111111111001;
        weights1[15112] <= 16'b0000000000001110;
        weights1[15113] <= 16'b0000000000000111;
        weights1[15114] <= 16'b0000000000001001;
        weights1[15115] <= 16'b1111111111110010;
        weights1[15116] <= 16'b1111111111101011;
        weights1[15117] <= 16'b1111111111111010;
        weights1[15118] <= 16'b1111111111111100;
        weights1[15119] <= 16'b1111111111111010;
        weights1[15120] <= 16'b0000000000000110;
        weights1[15121] <= 16'b0000000000001010;
        weights1[15122] <= 16'b0000000000000110;
        weights1[15123] <= 16'b0000000000010111;
        weights1[15124] <= 16'b0000000001001010;
        weights1[15125] <= 16'b0000000000100110;
        weights1[15126] <= 16'b0000000000100101;
        weights1[15127] <= 16'b0000000000110101;
        weights1[15128] <= 16'b0000000001001001;
        weights1[15129] <= 16'b0000000000001101;
        weights1[15130] <= 16'b0000000000100110;
        weights1[15131] <= 16'b0000000000010001;
        weights1[15132] <= 16'b0000000000000110;
        weights1[15133] <= 16'b1111111111111100;
        weights1[15134] <= 16'b0000000000000000;
        weights1[15135] <= 16'b1111111111111100;
        weights1[15136] <= 16'b0000000000000010;
        weights1[15137] <= 16'b1111111111111111;
        weights1[15138] <= 16'b0000000000000000;
        weights1[15139] <= 16'b0000000000000000;
        weights1[15140] <= 16'b1111111111111010;
        weights1[15141] <= 16'b1111111111111100;
        weights1[15142] <= 16'b1111111111111111;
        weights1[15143] <= 16'b0000000000010000;
        weights1[15144] <= 16'b1111111111101001;
        weights1[15145] <= 16'b1111111111110110;
        weights1[15146] <= 16'b1111111111111111;
        weights1[15147] <= 16'b1111111111110000;
        weights1[15148] <= 16'b0000000000001100;
        weights1[15149] <= 16'b0000000000001010;
        weights1[15150] <= 16'b0000000000011001;
        weights1[15151] <= 16'b0000000000010110;
        weights1[15152] <= 16'b0000000000100000;
        weights1[15153] <= 16'b0000000000110110;
        weights1[15154] <= 16'b0000000000010011;
        weights1[15155] <= 16'b0000000000100100;
        weights1[15156] <= 16'b0000000000000000;
        weights1[15157] <= 16'b0000000000100101;
        weights1[15158] <= 16'b0000000000011101;
        weights1[15159] <= 16'b0000000000011000;
        weights1[15160] <= 16'b0000000000010100;
        weights1[15161] <= 16'b0000000000011101;
        weights1[15162] <= 16'b0000000000100010;
        weights1[15163] <= 16'b0000000000001010;
        weights1[15164] <= 16'b1111111111110001;
        weights1[15165] <= 16'b0000000000001001;
        weights1[15166] <= 16'b1111111111101001;
        weights1[15167] <= 16'b1111111111101110;
        weights1[15168] <= 16'b0000000000001110;
        weights1[15169] <= 16'b1111111111111100;
        weights1[15170] <= 16'b1111111111111101;
        weights1[15171] <= 16'b1111111111110101;
        weights1[15172] <= 16'b0000000000000010;
        weights1[15173] <= 16'b1111111111110111;
        weights1[15174] <= 16'b0000000000001000;
        weights1[15175] <= 16'b1111111111101000;
        weights1[15176] <= 16'b0000000000010011;
        weights1[15177] <= 16'b0000000000010111;
        weights1[15178] <= 16'b0000000000011011;
        weights1[15179] <= 16'b0000000000000100;
        weights1[15180] <= 16'b0000000000011111;
        weights1[15181] <= 16'b0000000000100000;
        weights1[15182] <= 16'b0000000000010111;
        weights1[15183] <= 16'b0000000000100110;
        weights1[15184] <= 16'b0000000000011001;
        weights1[15185] <= 16'b0000000000111010;
        weights1[15186] <= 16'b0000000000100110;
        weights1[15187] <= 16'b0000000000110001;
        weights1[15188] <= 16'b0000000000110101;
        weights1[15189] <= 16'b0000000000011011;
        weights1[15190] <= 16'b0000000000100010;
        weights1[15191] <= 16'b0000000000011000;
        weights1[15192] <= 16'b0000000000000110;
        weights1[15193] <= 16'b0000000000001111;
        weights1[15194] <= 16'b0000000000001000;
        weights1[15195] <= 16'b0000000000001001;
        weights1[15196] <= 16'b0000000000000001;
        weights1[15197] <= 16'b1111111111110101;
        weights1[15198] <= 16'b1111111111110111;
        weights1[15199] <= 16'b1111111111101001;
        weights1[15200] <= 16'b1111111111111100;
        weights1[15201] <= 16'b1111111111111100;
        weights1[15202] <= 16'b1111111111111011;
        weights1[15203] <= 16'b1111111111110110;
        weights1[15204] <= 16'b0000000000011010;
        weights1[15205] <= 16'b0000000000100010;
        weights1[15206] <= 16'b0000000000010010;
        weights1[15207] <= 16'b0000000000001011;
        weights1[15208] <= 16'b0000000000011111;
        weights1[15209] <= 16'b0000000000000111;
        weights1[15210] <= 16'b0000000000001101;
        weights1[15211] <= 16'b0000000000111000;
        weights1[15212] <= 16'b1111111111110110;
        weights1[15213] <= 16'b0000000000011011;
        weights1[15214] <= 16'b0000000000111111;
        weights1[15215] <= 16'b0000000000011111;
        weights1[15216] <= 16'b0000000000011101;
        weights1[15217] <= 16'b0000000000000001;
        weights1[15218] <= 16'b0000000000000011;
        weights1[15219] <= 16'b0000000000000011;
        weights1[15220] <= 16'b0000000000001100;
        weights1[15221] <= 16'b1111111111111010;
        weights1[15222] <= 16'b0000000000000011;
        weights1[15223] <= 16'b1111111111110111;
        weights1[15224] <= 16'b0000000000000011;
        weights1[15225] <= 16'b1111111111111011;
        weights1[15226] <= 16'b0000000000010000;
        weights1[15227] <= 16'b0000000000000000;
        weights1[15228] <= 16'b1111111111111101;
        weights1[15229] <= 16'b1111111111111111;
        weights1[15230] <= 16'b1111111111111110;
        weights1[15231] <= 16'b1111111111100100;
        weights1[15232] <= 16'b0000000000001111;
        weights1[15233] <= 16'b0000000000001111;
        weights1[15234] <= 16'b0000000000010001;
        weights1[15235] <= 16'b0000000000010101;
        weights1[15236] <= 16'b0000000000100101;
        weights1[15237] <= 16'b0000000000010001;
        weights1[15238] <= 16'b0000000000010101;
        weights1[15239] <= 16'b0000000000101111;
        weights1[15240] <= 16'b0000000000010110;
        weights1[15241] <= 16'b0000000000010110;
        weights1[15242] <= 16'b0000000000000010;
        weights1[15243] <= 16'b1111111111101100;
        weights1[15244] <= 16'b1111111111111010;
        weights1[15245] <= 16'b1111111111100110;
        weights1[15246] <= 16'b1111111111101111;
        weights1[15247] <= 16'b1111111111110001;
        weights1[15248] <= 16'b1111111111011111;
        weights1[15249] <= 16'b0000000000001101;
        weights1[15250] <= 16'b1111111111111011;
        weights1[15251] <= 16'b0000000000011011;
        weights1[15252] <= 16'b1111111111111100;
        weights1[15253] <= 16'b0000000000000001;
        weights1[15254] <= 16'b0000000000010000;
        weights1[15255] <= 16'b1111111111101110;
        weights1[15256] <= 16'b1111111111110111;
        weights1[15257] <= 16'b0000000000010011;
        weights1[15258] <= 16'b0000000000001010;
        weights1[15259] <= 16'b1111111111110111;
        weights1[15260] <= 16'b0000000000001010;
        weights1[15261] <= 16'b1111111111111001;
        weights1[15262] <= 16'b0000000000010010;
        weights1[15263] <= 16'b0000000000010111;
        weights1[15264] <= 16'b0000000000001011;
        weights1[15265] <= 16'b0000000000001111;
        weights1[15266] <= 16'b0000000000011010;
        weights1[15267] <= 16'b0000000000001011;
        weights1[15268] <= 16'b0000000000000111;
        weights1[15269] <= 16'b1111111111010001;
        weights1[15270] <= 16'b1111111110111011;
        weights1[15271] <= 16'b1111111110101001;
        weights1[15272] <= 16'b1111111110100000;
        weights1[15273] <= 16'b1111111111000010;
        weights1[15274] <= 16'b1111111111010100;
        weights1[15275] <= 16'b1111111111100100;
        weights1[15276] <= 16'b1111111111110101;
        weights1[15277] <= 16'b1111111111111110;
        weights1[15278] <= 16'b1111111111111111;
        weights1[15279] <= 16'b1111111111101011;
        weights1[15280] <= 16'b1111111111111010;
        weights1[15281] <= 16'b1111111111111000;
        weights1[15282] <= 16'b0000000000000010;
        weights1[15283] <= 16'b0000000000001000;
        weights1[15284] <= 16'b0000000000001000;
        weights1[15285] <= 16'b1111111111110001;
        weights1[15286] <= 16'b0000000000010011;
        weights1[15287] <= 16'b1111111111101010;
        weights1[15288] <= 16'b1111111111101011;
        weights1[15289] <= 16'b1111111111011000;
        weights1[15290] <= 16'b1111111111101101;
        weights1[15291] <= 16'b1111111111111000;
        weights1[15292] <= 16'b1111111111111111;
        weights1[15293] <= 16'b0000000000000001;
        weights1[15294] <= 16'b1111111111000110;
        weights1[15295] <= 16'b1111111110110011;
        weights1[15296] <= 16'b1111111101111101;
        weights1[15297] <= 16'b1111111100011110;
        weights1[15298] <= 16'b1111111101111100;
        weights1[15299] <= 16'b1111111110011110;
        weights1[15300] <= 16'b1111111111011001;
        weights1[15301] <= 16'b1111111111001101;
        weights1[15302] <= 16'b1111111111100101;
        weights1[15303] <= 16'b1111111111111000;
        weights1[15304] <= 16'b1111111111111000;
        weights1[15305] <= 16'b1111111111111110;
        weights1[15306] <= 16'b1111111111101110;
        weights1[15307] <= 16'b0000000000000010;
        weights1[15308] <= 16'b1111111111111000;
        weights1[15309] <= 16'b1111111111111111;
        weights1[15310] <= 16'b1111111111110110;
        weights1[15311] <= 16'b0000000000011000;
        weights1[15312] <= 16'b1111111111101001;
        weights1[15313] <= 16'b1111111111111100;
        weights1[15314] <= 16'b1111111111111111;
        weights1[15315] <= 16'b1111111111110111;
        weights1[15316] <= 16'b1111111111011001;
        weights1[15317] <= 16'b1111111110111101;
        weights1[15318] <= 16'b1111111111000010;
        weights1[15319] <= 16'b1111111110111111;
        weights1[15320] <= 16'b1111111110100100;
        weights1[15321] <= 16'b1111111110011001;
        weights1[15322] <= 16'b1111111101100100;
        weights1[15323] <= 16'b1111111100000110;
        weights1[15324] <= 16'b1111111100010011;
        weights1[15325] <= 16'b1111111110000111;
        weights1[15326] <= 16'b1111111111011101;
        weights1[15327] <= 16'b0000000000000000;
        weights1[15328] <= 16'b0000000000000000;
        weights1[15329] <= 16'b0000000000000110;
        weights1[15330] <= 16'b0000000000001110;
        weights1[15331] <= 16'b0000000000000111;
        weights1[15332] <= 16'b0000000000001101;
        weights1[15333] <= 16'b0000000000010001;
        weights1[15334] <= 16'b0000000000000101;
        weights1[15335] <= 16'b0000000000000000;
        weights1[15336] <= 16'b0000000000011010;
        weights1[15337] <= 16'b0000000000010001;
        weights1[15338] <= 16'b0000000000000100;
        weights1[15339] <= 16'b0000000000001111;
        weights1[15340] <= 16'b0000000000001001;
        weights1[15341] <= 16'b0000000000000010;
        weights1[15342] <= 16'b0000000000000011;
        weights1[15343] <= 16'b0000000000000101;
        weights1[15344] <= 16'b1111111111000001;
        weights1[15345] <= 16'b1111111110110100;
        weights1[15346] <= 16'b1111111110101011;
        weights1[15347] <= 16'b1111111110001111;
        weights1[15348] <= 16'b1111111101010110;
        weights1[15349] <= 16'b1111111100111001;
        weights1[15350] <= 16'b1111111100100010;
        weights1[15351] <= 16'b1111111101010101;
        weights1[15352] <= 16'b1111111111110010;
        weights1[15353] <= 16'b0000000000010100;
        weights1[15354] <= 16'b0000000000001101;
        weights1[15355] <= 16'b0000000000001110;
        weights1[15356] <= 16'b0000000000100000;
        weights1[15357] <= 16'b0000000000001010;
        weights1[15358] <= 16'b0000000000000001;
        weights1[15359] <= 16'b0000000000000011;
        weights1[15360] <= 16'b0000000000010011;
        weights1[15361] <= 16'b0000000000010001;
        weights1[15362] <= 16'b0000000000010000;
        weights1[15363] <= 16'b0000000000000010;
        weights1[15364] <= 16'b0000000000000011;
        weights1[15365] <= 16'b0000000000000000;
        weights1[15366] <= 16'b0000000000001010;
        weights1[15367] <= 16'b0000000000000011;
        weights1[15368] <= 16'b1111111111111111;
        weights1[15369] <= 16'b0000000000011000;
        weights1[15370] <= 16'b1111111111111001;
        weights1[15371] <= 16'b0000000000000101;
        weights1[15372] <= 16'b1111111110111110;
        weights1[15373] <= 16'b1111111110110100;
        weights1[15374] <= 16'b1111111110100001;
        weights1[15375] <= 16'b1111111110001100;
        weights1[15376] <= 16'b1111111110000010;
        weights1[15377] <= 16'b1111111110010110;
        weights1[15378] <= 16'b1111111110101001;
        weights1[15379] <= 16'b0000000000001011;
        weights1[15380] <= 16'b0000000000000111;
        weights1[15381] <= 16'b0000000000011001;
        weights1[15382] <= 16'b0000000000010100;
        weights1[15383] <= 16'b0000000000011011;
        weights1[15384] <= 16'b0000000000001101;
        weights1[15385] <= 16'b0000000000001110;
        weights1[15386] <= 16'b0000000000001101;
        weights1[15387] <= 16'b0000000000000000;
        weights1[15388] <= 16'b1111111111111000;
        weights1[15389] <= 16'b0000000000000000;
        weights1[15390] <= 16'b0000000000001100;
        weights1[15391] <= 16'b0000000000000000;
        weights1[15392] <= 16'b0000000000011111;
        weights1[15393] <= 16'b1111111111111111;
        weights1[15394] <= 16'b1111111111110110;
        weights1[15395] <= 16'b0000000000001000;
        weights1[15396] <= 16'b0000000000000101;
        weights1[15397] <= 16'b1111111111111010;
        weights1[15398] <= 16'b1111111111110001;
        weights1[15399] <= 16'b1111111111110100;
        weights1[15400] <= 16'b1111111111000101;
        weights1[15401] <= 16'b1111111110111100;
        weights1[15402] <= 16'b1111111110101001;
        weights1[15403] <= 16'b1111111110101001;
        weights1[15404] <= 16'b1111111111001100;
        weights1[15405] <= 16'b1111111111110010;
        weights1[15406] <= 16'b0000000000000100;
        weights1[15407] <= 16'b0000000000101010;
        weights1[15408] <= 16'b0000000000110000;
        weights1[15409] <= 16'b0000000000001100;
        weights1[15410] <= 16'b0000000000011001;
        weights1[15411] <= 16'b0000000000010001;
        weights1[15412] <= 16'b1111111111111011;
        weights1[15413] <= 16'b0000000000000010;
        weights1[15414] <= 16'b0000000000000100;
        weights1[15415] <= 16'b0000000000001110;
        weights1[15416] <= 16'b0000000000000010;
        weights1[15417] <= 16'b1111111111111010;
        weights1[15418] <= 16'b1111111111111111;
        weights1[15419] <= 16'b0000000000000100;
        weights1[15420] <= 16'b0000000000000010;
        weights1[15421] <= 16'b0000000000000011;
        weights1[15422] <= 16'b0000000000001111;
        weights1[15423] <= 16'b1111111111110110;
        weights1[15424] <= 16'b1111111111110000;
        weights1[15425] <= 16'b1111111111111011;
        weights1[15426] <= 16'b0000000000001001;
        weights1[15427] <= 16'b0000000000100000;
        weights1[15428] <= 16'b1111111111010111;
        weights1[15429] <= 16'b1111111111010001;
        weights1[15430] <= 16'b1111111111001110;
        weights1[15431] <= 16'b1111111111001111;
        weights1[15432] <= 16'b1111111111101111;
        weights1[15433] <= 16'b0000000000100000;
        weights1[15434] <= 16'b0000000000000101;
        weights1[15435] <= 16'b0000000000010001;
        weights1[15436] <= 16'b0000000000000011;
        weights1[15437] <= 16'b0000000000000000;
        weights1[15438] <= 16'b1111111111111100;
        weights1[15439] <= 16'b1111111111111100;
        weights1[15440] <= 16'b0000000000000111;
        weights1[15441] <= 16'b1111111111111001;
        weights1[15442] <= 16'b0000000000000111;
        weights1[15443] <= 16'b0000000000000011;
        weights1[15444] <= 16'b0000000000001011;
        weights1[15445] <= 16'b1111111111111101;
        weights1[15446] <= 16'b1111111111101011;
        weights1[15447] <= 16'b0000000000000101;
        weights1[15448] <= 16'b0000000000000000;
        weights1[15449] <= 16'b0000000000000010;
        weights1[15450] <= 16'b0000000000000011;
        weights1[15451] <= 16'b0000000000010100;
        weights1[15452] <= 16'b1111111111111010;
        weights1[15453] <= 16'b1111111111111111;
        weights1[15454] <= 16'b1111111111111111;
        weights1[15455] <= 16'b0000000000010110;
        weights1[15456] <= 16'b1111111111101111;
        weights1[15457] <= 16'b1111111111101011;
        weights1[15458] <= 16'b1111111111111001;
        weights1[15459] <= 16'b1111111111111011;
        weights1[15460] <= 16'b0000000000100001;
        weights1[15461] <= 16'b1111111111111001;
        weights1[15462] <= 16'b1111111111101010;
        weights1[15463] <= 16'b1111111111111100;
        weights1[15464] <= 16'b0000000000001000;
        weights1[15465] <= 16'b0000000000010101;
        weights1[15466] <= 16'b1111111111101101;
        weights1[15467] <= 16'b0000000000001100;
        weights1[15468] <= 16'b1111111111111001;
        weights1[15469] <= 16'b1111111111111101;
        weights1[15470] <= 16'b0000000000000010;
        weights1[15471] <= 16'b1111111111111001;
        weights1[15472] <= 16'b0000000000000001;
        weights1[15473] <= 16'b1111111111111101;
        weights1[15474] <= 16'b0000000000001110;
        weights1[15475] <= 16'b0000000000000110;
        weights1[15476] <= 16'b1111111111111110;
        weights1[15477] <= 16'b1111111111110011;
        weights1[15478] <= 16'b0000000000000110;
        weights1[15479] <= 16'b0000000000000101;
        weights1[15480] <= 16'b1111111111111111;
        weights1[15481] <= 16'b1111111111111001;
        weights1[15482] <= 16'b1111111111111111;
        weights1[15483] <= 16'b0000000000000001;
        weights1[15484] <= 16'b1111111111111010;
        weights1[15485] <= 16'b1111111111111100;
        weights1[15486] <= 16'b0000000000001111;
        weights1[15487] <= 16'b0000000000001011;
        weights1[15488] <= 16'b0000000000000011;
        weights1[15489] <= 16'b1111111111111101;
        weights1[15490] <= 16'b1111111111111011;
        weights1[15491] <= 16'b0000000000000100;
        weights1[15492] <= 16'b1111111111111010;
        weights1[15493] <= 16'b1111111111110110;
        weights1[15494] <= 16'b0000000000010000;
        weights1[15495] <= 16'b1111111111101000;
        weights1[15496] <= 16'b0000000000010000;
        weights1[15497] <= 16'b0000000000000001;
        weights1[15498] <= 16'b0000000000000001;
        weights1[15499] <= 16'b1111111111111011;
        weights1[15500] <= 16'b1111111111111101;
        weights1[15501] <= 16'b1111111111110001;
        weights1[15502] <= 16'b1111111111111001;
        weights1[15503] <= 16'b1111111111111000;
        weights1[15504] <= 16'b1111111111111100;
        weights1[15505] <= 16'b1111111111111000;
        weights1[15506] <= 16'b0000000000000000;
        weights1[15507] <= 16'b0000000000001000;
        weights1[15508] <= 16'b1111111111111010;
        weights1[15509] <= 16'b0000000000000101;
        weights1[15510] <= 16'b1111111111111011;
        weights1[15511] <= 16'b1111111111111110;
        weights1[15512] <= 16'b0000000000001001;
        weights1[15513] <= 16'b1111111111111111;
        weights1[15514] <= 16'b0000000000001110;
        weights1[15515] <= 16'b0000000000010001;
        weights1[15516] <= 16'b0000000000001010;
        weights1[15517] <= 16'b1111111111111011;
        weights1[15518] <= 16'b0000000000011100;
        weights1[15519] <= 16'b1111111111111011;
        weights1[15520] <= 16'b1111111111111111;
        weights1[15521] <= 16'b1111111111111111;
        weights1[15522] <= 16'b0000000000011011;
        weights1[15523] <= 16'b1111111111110011;
        weights1[15524] <= 16'b0000000000000110;
        weights1[15525] <= 16'b1111111111111010;
        weights1[15526] <= 16'b1111111111111000;
        weights1[15527] <= 16'b1111111111110000;
        weights1[15528] <= 16'b1111111111110001;
        weights1[15529] <= 16'b0000000000001010;
        weights1[15530] <= 16'b1111111111101100;
        weights1[15531] <= 16'b0000000000001001;
        weights1[15532] <= 16'b0000000000001001;
        weights1[15533] <= 16'b1111111111111100;
        weights1[15534] <= 16'b0000000000000101;
        weights1[15535] <= 16'b0000000000000001;
        weights1[15536] <= 16'b1111111111111101;
        weights1[15537] <= 16'b1111111111111110;
        weights1[15538] <= 16'b0000000000000001;
        weights1[15539] <= 16'b0000000000000011;
        weights1[15540] <= 16'b0000000000000011;
        weights1[15541] <= 16'b0000000000000001;
        weights1[15542] <= 16'b0000000000010001;
        weights1[15543] <= 16'b0000000000001100;
        weights1[15544] <= 16'b1111111111111110;
        weights1[15545] <= 16'b0000000000011010;
        weights1[15546] <= 16'b0000000000010010;
        weights1[15547] <= 16'b0000000000011100;
        weights1[15548] <= 16'b1111111111111100;
        weights1[15549] <= 16'b0000000000000101;
        weights1[15550] <= 16'b1111111111111110;
        weights1[15551] <= 16'b0000000000001011;
        weights1[15552] <= 16'b0000000000000000;
        weights1[15553] <= 16'b1111111111110111;
        weights1[15554] <= 16'b0000000000000010;
        weights1[15555] <= 16'b0000000000010000;
        weights1[15556] <= 16'b0000000000000110;
        weights1[15557] <= 16'b1111111111110110;
        weights1[15558] <= 16'b0000000000010100;
        weights1[15559] <= 16'b1111111111101111;
        weights1[15560] <= 16'b0000000000000111;
        weights1[15561] <= 16'b1111111111110100;
        weights1[15562] <= 16'b0000000000000001;
        weights1[15563] <= 16'b0000000000000111;
        weights1[15564] <= 16'b0000000000000001;
        weights1[15565] <= 16'b1111111111111011;
        weights1[15566] <= 16'b1111111111111101;
        weights1[15567] <= 16'b0000000000000111;
        weights1[15568] <= 16'b0000000000000001;
        weights1[15569] <= 16'b0000000000000011;
        weights1[15570] <= 16'b0000000000001110;
        weights1[15571] <= 16'b0000000000000101;
        weights1[15572] <= 16'b0000000000000001;
        weights1[15573] <= 16'b0000000000001001;
        weights1[15574] <= 16'b1111111111101110;
        weights1[15575] <= 16'b0000000000001100;
        weights1[15576] <= 16'b1111111111011010;
        weights1[15577] <= 16'b0000000000011100;
        weights1[15578] <= 16'b1111111111111111;
        weights1[15579] <= 16'b0000000000010110;
        weights1[15580] <= 16'b0000000000000110;
        weights1[15581] <= 16'b1111111111110110;
        weights1[15582] <= 16'b0000000000010110;
        weights1[15583] <= 16'b0000000000000001;
        weights1[15584] <= 16'b1111111111111111;
        weights1[15585] <= 16'b0000000000001110;
        weights1[15586] <= 16'b0000000000001010;
        weights1[15587] <= 16'b1111111111111111;
        weights1[15588] <= 16'b0000000000000010;
        weights1[15589] <= 16'b0000000000001011;
        weights1[15590] <= 16'b1111111111111010;
        weights1[15591] <= 16'b1111111111110010;
        weights1[15592] <= 16'b1111111111110111;
        weights1[15593] <= 16'b0000000000000000;
        weights1[15594] <= 16'b1111111111110001;
        weights1[15595] <= 16'b0000000000000001;
        weights1[15596] <= 16'b1111111111111111;
        weights1[15597] <= 16'b0000000000000011;
        weights1[15598] <= 16'b0000000000001100;
        weights1[15599] <= 16'b1111111111111000;
        weights1[15600] <= 16'b0000000000000110;
        weights1[15601] <= 16'b1111111111110011;
        weights1[15602] <= 16'b1111111111110011;
        weights1[15603] <= 16'b0000000000000101;
        weights1[15604] <= 16'b0000000000010010;
        weights1[15605] <= 16'b0000000000001011;
        weights1[15606] <= 16'b1111111111010110;
        weights1[15607] <= 16'b1111111111111000;
        weights1[15608] <= 16'b0000000000000111;
        weights1[15609] <= 16'b0000000000001100;
        weights1[15610] <= 16'b0000000000001100;
        weights1[15611] <= 16'b1111111111110010;
        weights1[15612] <= 16'b0000000000000010;
        weights1[15613] <= 16'b1111111111111000;
        weights1[15614] <= 16'b0000000000000101;
        weights1[15615] <= 16'b1111111111111100;
        weights1[15616] <= 16'b0000000000010010;
        weights1[15617] <= 16'b1111111111111111;
        weights1[15618] <= 16'b0000000000000000;
        weights1[15619] <= 16'b1111111111111001;
        weights1[15620] <= 16'b1111111111101101;
        weights1[15621] <= 16'b1111111111110110;
        weights1[15622] <= 16'b1111111111110000;
        weights1[15623] <= 16'b0000000000000011;
        weights1[15624] <= 16'b0000000000000010;
        weights1[15625] <= 16'b1111111111111110;
        weights1[15626] <= 16'b0000000000001000;
        weights1[15627] <= 16'b1111111111111100;
        weights1[15628] <= 16'b1111111111111011;
        weights1[15629] <= 16'b1111111111011110;
        weights1[15630] <= 16'b1111111111110100;
        weights1[15631] <= 16'b0000000000001011;
        weights1[15632] <= 16'b0000000000000000;
        weights1[15633] <= 16'b0000000000000101;
        weights1[15634] <= 16'b0000000000010001;
        weights1[15635] <= 16'b0000000000000011;
        weights1[15636] <= 16'b0000000000001000;
        weights1[15637] <= 16'b1111111111110111;
        weights1[15638] <= 16'b0000000000000001;
        weights1[15639] <= 16'b1111111111111101;
        weights1[15640] <= 16'b1111111111111000;
        weights1[15641] <= 16'b1111111111111110;
        weights1[15642] <= 16'b1111111111101011;
        weights1[15643] <= 16'b0000000000000011;
        weights1[15644] <= 16'b1111111111111000;
        weights1[15645] <= 16'b0000000000001001;
        weights1[15646] <= 16'b0000000000000101;
        weights1[15647] <= 16'b1111111111111110;
        weights1[15648] <= 16'b1111111111110101;
        weights1[15649] <= 16'b1111111111111101;
        weights1[15650] <= 16'b0000000000000001;
        weights1[15651] <= 16'b0000000000000001;
        weights1[15652] <= 16'b0000000000000010;
        weights1[15653] <= 16'b1111111111111111;
        weights1[15654] <= 16'b0000000000001010;
        weights1[15655] <= 16'b0000000000010001;
        weights1[15656] <= 16'b0000000000001110;
        weights1[15657] <= 16'b0000000000000011;
        weights1[15658] <= 16'b0000000000001111;
        weights1[15659] <= 16'b0000000000001101;
        weights1[15660] <= 16'b0000000000000111;
        weights1[15661] <= 16'b1111111111111011;
        weights1[15662] <= 16'b0000000000001000;
        weights1[15663] <= 16'b0000000000001010;
        weights1[15664] <= 16'b1111111111111001;
        weights1[15665] <= 16'b0000000000001001;
        weights1[15666] <= 16'b0000000000000010;
        weights1[15667] <= 16'b1111111111111011;
        weights1[15668] <= 16'b1111111111111111;
        weights1[15669] <= 16'b0000000000010100;
        weights1[15670] <= 16'b1111111111110011;
        weights1[15671] <= 16'b1111111111110111;
        weights1[15672] <= 16'b1111111111111001;
        weights1[15673] <= 16'b1111111111111001;
        weights1[15674] <= 16'b1111111111110000;
        weights1[15675] <= 16'b1111111111111110;
        weights1[15676] <= 16'b1111111111111011;
        weights1[15677] <= 16'b1111111111111110;
        weights1[15678] <= 16'b0000000000000011;
        weights1[15679] <= 16'b0000000000000011;
        weights1[15680] <= 16'b0000000000000000;
        weights1[15681] <= 16'b0000000000000000;
        weights1[15682] <= 16'b0000000000000000;
        weights1[15683] <= 16'b0000000000000000;
        weights1[15684] <= 16'b0000000000000000;
        weights1[15685] <= 16'b1111111111111111;
        weights1[15686] <= 16'b1111111111111101;
        weights1[15687] <= 16'b1111111111111101;
        weights1[15688] <= 16'b1111111111111101;
        weights1[15689] <= 16'b1111111111111010;
        weights1[15690] <= 16'b1111111111111011;
        weights1[15691] <= 16'b1111111111110101;
        weights1[15692] <= 16'b1111111111101110;
        weights1[15693] <= 16'b1111111111110010;
        weights1[15694] <= 16'b1111111111110100;
        weights1[15695] <= 16'b1111111111110110;
        weights1[15696] <= 16'b1111111111110110;
        weights1[15697] <= 16'b1111111111110011;
        weights1[15698] <= 16'b1111111111110110;
        weights1[15699] <= 16'b1111111111110110;
        weights1[15700] <= 16'b1111111111111011;
        weights1[15701] <= 16'b1111111111111011;
        weights1[15702] <= 16'b1111111111111101;
        weights1[15703] <= 16'b1111111111111111;
        weights1[15704] <= 16'b1111111111111110;
        weights1[15705] <= 16'b0000000000000000;
        weights1[15706] <= 16'b0000000000000000;
        weights1[15707] <= 16'b0000000000000000;
        weights1[15708] <= 16'b0000000000000000;
        weights1[15709] <= 16'b0000000000000000;
        weights1[15710] <= 16'b0000000000000000;
        weights1[15711] <= 16'b1111111111111110;
        weights1[15712] <= 16'b1111111111111110;
        weights1[15713] <= 16'b1111111111111010;
        weights1[15714] <= 16'b1111111111111000;
        weights1[15715] <= 16'b1111111111111001;
        weights1[15716] <= 16'b1111111111111000;
        weights1[15717] <= 16'b1111111111110101;
        weights1[15718] <= 16'b1111111111101101;
        weights1[15719] <= 16'b1111111111110000;
        weights1[15720] <= 16'b1111111111101110;
        weights1[15721] <= 16'b1111111111101110;
        weights1[15722] <= 16'b1111111111101101;
        weights1[15723] <= 16'b1111111111110001;
        weights1[15724] <= 16'b1111111111101100;
        weights1[15725] <= 16'b1111111111101110;
        weights1[15726] <= 16'b1111111111101101;
        weights1[15727] <= 16'b1111111111101111;
        weights1[15728] <= 16'b1111111111101110;
        weights1[15729] <= 16'b1111111111100101;
        weights1[15730] <= 16'b1111111111101100;
        weights1[15731] <= 16'b1111111111110111;
        weights1[15732] <= 16'b1111111111111110;
        weights1[15733] <= 16'b1111111111111111;
        weights1[15734] <= 16'b0000000000000001;
        weights1[15735] <= 16'b0000000000000000;
        weights1[15736] <= 16'b0000000000000000;
        weights1[15737] <= 16'b0000000000000000;
        weights1[15738] <= 16'b0000000000000000;
        weights1[15739] <= 16'b1111111111111101;
        weights1[15740] <= 16'b1111111111111010;
        weights1[15741] <= 16'b1111111111110101;
        weights1[15742] <= 16'b1111111111110101;
        weights1[15743] <= 16'b1111111111110010;
        weights1[15744] <= 16'b1111111111101110;
        weights1[15745] <= 16'b1111111111101110;
        weights1[15746] <= 16'b1111111111100011;
        weights1[15747] <= 16'b1111111111100101;
        weights1[15748] <= 16'b1111111111100101;
        weights1[15749] <= 16'b1111111111100100;
        weights1[15750] <= 16'b1111111111100100;
        weights1[15751] <= 16'b1111111111100111;
        weights1[15752] <= 16'b1111111111011110;
        weights1[15753] <= 16'b1111111111100010;
        weights1[15754] <= 16'b1111111111011111;
        weights1[15755] <= 16'b1111111111100111;
        weights1[15756] <= 16'b1111111111100101;
        weights1[15757] <= 16'b1111111111100101;
        weights1[15758] <= 16'b1111111111100000;
        weights1[15759] <= 16'b1111111111101111;
        weights1[15760] <= 16'b1111111111110101;
        weights1[15761] <= 16'b1111111111111011;
        weights1[15762] <= 16'b1111111111111100;
        weights1[15763] <= 16'b1111111111111110;
        weights1[15764] <= 16'b0000000000000000;
        weights1[15765] <= 16'b0000000000000000;
        weights1[15766] <= 16'b1111111111111100;
        weights1[15767] <= 16'b1111111111111001;
        weights1[15768] <= 16'b1111111111110100;
        weights1[15769] <= 16'b1111111111110000;
        weights1[15770] <= 16'b1111111111100011;
        weights1[15771] <= 16'b1111111111100011;
        weights1[15772] <= 16'b1111111111011111;
        weights1[15773] <= 16'b1111111111011000;
        weights1[15774] <= 16'b1111111111011000;
        weights1[15775] <= 16'b1111111111100001;
        weights1[15776] <= 16'b1111111111011100;
        weights1[15777] <= 16'b1111111111011001;
        weights1[15778] <= 16'b1111111111011101;
        weights1[15779] <= 16'b1111111111011100;
        weights1[15780] <= 16'b1111111111011100;
        weights1[15781] <= 16'b1111111111011010;
        weights1[15782] <= 16'b1111111111100101;
        weights1[15783] <= 16'b1111111111100010;
        weights1[15784] <= 16'b1111111111011110;
        weights1[15785] <= 16'b1111111111011000;
        weights1[15786] <= 16'b1111111111100110;
        weights1[15787] <= 16'b1111111111101011;
        weights1[15788] <= 16'b1111111111110000;
        weights1[15789] <= 16'b1111111111110101;
        weights1[15790] <= 16'b1111111111111001;
        weights1[15791] <= 16'b1111111111111110;
        weights1[15792] <= 16'b0000000000000000;
        weights1[15793] <= 16'b1111111111111110;
        weights1[15794] <= 16'b1111111111110101;
        weights1[15795] <= 16'b1111111111101110;
        weights1[15796] <= 16'b1111111111101000;
        weights1[15797] <= 16'b1111111111100001;
        weights1[15798] <= 16'b1111111111100000;
        weights1[15799] <= 16'b1111111111011100;
        weights1[15800] <= 16'b1111111111011011;
        weights1[15801] <= 16'b1111111111001101;
        weights1[15802] <= 16'b1111111111010101;
        weights1[15803] <= 16'b1111111111010111;
        weights1[15804] <= 16'b1111111111010110;
        weights1[15805] <= 16'b1111111111010100;
        weights1[15806] <= 16'b1111111111001111;
        weights1[15807] <= 16'b1111111111010011;
        weights1[15808] <= 16'b1111111111010101;
        weights1[15809] <= 16'b1111111111010111;
        weights1[15810] <= 16'b1111111111011101;
        weights1[15811] <= 16'b1111111111100011;
        weights1[15812] <= 16'b1111111111011000;
        weights1[15813] <= 16'b1111111111010011;
        weights1[15814] <= 16'b1111111111011011;
        weights1[15815] <= 16'b1111111111101000;
        weights1[15816] <= 16'b1111111111101100;
        weights1[15817] <= 16'b1111111111101101;
        weights1[15818] <= 16'b1111111111110001;
        weights1[15819] <= 16'b1111111111110110;
        weights1[15820] <= 16'b0000000000000001;
        weights1[15821] <= 16'b1111111111111001;
        weights1[15822] <= 16'b1111111111101011;
        weights1[15823] <= 16'b1111111111011101;
        weights1[15824] <= 16'b1111111111010011;
        weights1[15825] <= 16'b1111111111001100;
        weights1[15826] <= 16'b1111111111001010;
        weights1[15827] <= 16'b1111111111000110;
        weights1[15828] <= 16'b1111111111000000;
        weights1[15829] <= 16'b1111111110110001;
        weights1[15830] <= 16'b1111111111000001;
        weights1[15831] <= 16'b1111111111001101;
        weights1[15832] <= 16'b1111111111000111;
        weights1[15833] <= 16'b1111111111001100;
        weights1[15834] <= 16'b1111111111001111;
        weights1[15835] <= 16'b1111111111001110;
        weights1[15836] <= 16'b1111111111000100;
        weights1[15837] <= 16'b1111111111001010;
        weights1[15838] <= 16'b1111111111010011;
        weights1[15839] <= 16'b1111111111010011;
        weights1[15840] <= 16'b1111111111001001;
        weights1[15841] <= 16'b1111111111001000;
        weights1[15842] <= 16'b1111111111011000;
        weights1[15843] <= 16'b1111111111011101;
        weights1[15844] <= 16'b1111111111011111;
        weights1[15845] <= 16'b1111111111101001;
        weights1[15846] <= 16'b1111111111101011;
        weights1[15847] <= 16'b1111111111110001;
        weights1[15848] <= 16'b1111111111111110;
        weights1[15849] <= 16'b1111111111110110;
        weights1[15850] <= 16'b1111111111101101;
        weights1[15851] <= 16'b1111111111010101;
        weights1[15852] <= 16'b1111111111000010;
        weights1[15853] <= 16'b1111111110110101;
        weights1[15854] <= 16'b1111111110101001;
        weights1[15855] <= 16'b1111111110011101;
        weights1[15856] <= 16'b1111111110100110;
        weights1[15857] <= 16'b1111111110010100;
        weights1[15858] <= 16'b1111111110011000;
        weights1[15859] <= 16'b1111111110100000;
        weights1[15860] <= 16'b1111111110101011;
        weights1[15861] <= 16'b1111111110011101;
        weights1[15862] <= 16'b1111111110101010;
        weights1[15863] <= 16'b1111111110011011;
        weights1[15864] <= 16'b1111111110111000;
        weights1[15865] <= 16'b1111111110110001;
        weights1[15866] <= 16'b1111111110101110;
        weights1[15867] <= 16'b1111111110111010;
        weights1[15868] <= 16'b1111111110111011;
        weights1[15869] <= 16'b1111111110111111;
        weights1[15870] <= 16'b1111111111001101;
        weights1[15871] <= 16'b1111111111011011;
        weights1[15872] <= 16'b1111111111011110;
        weights1[15873] <= 16'b1111111111011110;
        weights1[15874] <= 16'b1111111111100110;
        weights1[15875] <= 16'b1111111111110000;
        weights1[15876] <= 16'b1111111111111101;
        weights1[15877] <= 16'b1111111111110100;
        weights1[15878] <= 16'b1111111111100110;
        weights1[15879] <= 16'b1111111111000111;
        weights1[15880] <= 16'b1111111110110011;
        weights1[15881] <= 16'b1111111110011111;
        weights1[15882] <= 16'b1111111110000000;
        weights1[15883] <= 16'b1111111110000111;
        weights1[15884] <= 16'b1111111110100110;
        weights1[15885] <= 16'b1111111110010000;
        weights1[15886] <= 16'b1111111110001010;
        weights1[15887] <= 16'b1111111110010000;
        weights1[15888] <= 16'b1111111110010111;
        weights1[15889] <= 16'b1111111110010011;
        weights1[15890] <= 16'b1111111110011111;
        weights1[15891] <= 16'b1111111110100101;
        weights1[15892] <= 16'b1111111110111011;
        weights1[15893] <= 16'b1111111110010111;
        weights1[15894] <= 16'b1111111110010101;
        weights1[15895] <= 16'b1111111110100101;
        weights1[15896] <= 16'b1111111110010101;
        weights1[15897] <= 16'b1111111110101100;
        weights1[15898] <= 16'b1111111110111100;
        weights1[15899] <= 16'b1111111111001011;
        weights1[15900] <= 16'b1111111111001101;
        weights1[15901] <= 16'b1111111111011101;
        weights1[15902] <= 16'b1111111111011101;
        weights1[15903] <= 16'b1111111111101101;
        weights1[15904] <= 16'b1111111111111100;
        weights1[15905] <= 16'b1111111111110101;
        weights1[15906] <= 16'b1111111111100100;
        weights1[15907] <= 16'b1111111111001101;
        weights1[15908] <= 16'b1111111110111100;
        weights1[15909] <= 16'b1111111110101010;
        weights1[15910] <= 16'b1111111110111010;
        weights1[15911] <= 16'b1111111111001101;
        weights1[15912] <= 16'b1111111110110000;
        weights1[15913] <= 16'b1111111110101110;
        weights1[15914] <= 16'b1111111110111010;
        weights1[15915] <= 16'b1111111111000100;
        weights1[15916] <= 16'b1111111111001000;
        weights1[15917] <= 16'b1111111111011010;
        weights1[15918] <= 16'b1111111111001010;
        weights1[15919] <= 16'b1111111111010110;
        weights1[15920] <= 16'b1111111110111110;
        weights1[15921] <= 16'b1111111110111111;
        weights1[15922] <= 16'b1111111111000110;
        weights1[15923] <= 16'b1111111111010011;
        weights1[15924] <= 16'b1111111111001111;
        weights1[15925] <= 16'b1111111111100010;
        weights1[15926] <= 16'b1111111110111111;
        weights1[15927] <= 16'b1111111110111101;
        weights1[15928] <= 16'b1111111111000110;
        weights1[15929] <= 16'b1111111111100001;
        weights1[15930] <= 16'b1111111111110000;
        weights1[15931] <= 16'b1111111111111000;
        weights1[15932] <= 16'b0000000000000111;
        weights1[15933] <= 16'b1111111111111100;
        weights1[15934] <= 16'b1111111111101010;
        weights1[15935] <= 16'b1111111111101000;
        weights1[15936] <= 16'b1111111111101100;
        weights1[15937] <= 16'b1111111111101101;
        weights1[15938] <= 16'b1111111111110001;
        weights1[15939] <= 16'b1111111111110011;
        weights1[15940] <= 16'b1111111111111011;
        weights1[15941] <= 16'b1111111111011100;
        weights1[15942] <= 16'b1111111111001111;
        weights1[15943] <= 16'b1111111111011001;
        weights1[15944] <= 16'b1111111111011100;
        weights1[15945] <= 16'b1111111111011111;
        weights1[15946] <= 16'b1111111111001100;
        weights1[15947] <= 16'b1111111111100000;
        weights1[15948] <= 16'b1111111111010111;
        weights1[15949] <= 16'b1111111111101010;
        weights1[15950] <= 16'b1111111111010011;
        weights1[15951] <= 16'b1111111111011100;
        weights1[15952] <= 16'b1111111111100010;
        weights1[15953] <= 16'b1111111111110111;
        weights1[15954] <= 16'b1111111111010110;
        weights1[15955] <= 16'b1111111111101110;
        weights1[15956] <= 16'b1111111111101111;
        weights1[15957] <= 16'b1111111111111000;
        weights1[15958] <= 16'b1111111111111000;
        weights1[15959] <= 16'b0000000000001110;
        weights1[15960] <= 16'b0000000000001010;
        weights1[15961] <= 16'b0000000000000110;
        weights1[15962] <= 16'b1111111111110010;
        weights1[15963] <= 16'b1111111111111011;
        weights1[15964] <= 16'b1111111111111101;
        weights1[15965] <= 16'b0000000000000000;
        weights1[15966] <= 16'b0000000000000011;
        weights1[15967] <= 16'b0000000000100100;
        weights1[15968] <= 16'b0000000000000100;
        weights1[15969] <= 16'b0000000000100000;
        weights1[15970] <= 16'b0000000000000000;
        weights1[15971] <= 16'b1111111111110100;
        weights1[15972] <= 16'b1111111111010111;
        weights1[15973] <= 16'b1111111111010101;
        weights1[15974] <= 16'b1111111111011010;
        weights1[15975] <= 16'b1111111111100011;
        weights1[15976] <= 16'b1111111111100101;
        weights1[15977] <= 16'b1111111111111101;
        weights1[15978] <= 16'b1111111111101000;
        weights1[15979] <= 16'b1111111111100101;
        weights1[15980] <= 16'b0000000000000000;
        weights1[15981] <= 16'b1111111111110000;
        weights1[15982] <= 16'b0000000000011001;
        weights1[15983] <= 16'b1111111111110010;
        weights1[15984] <= 16'b1111111111110000;
        weights1[15985] <= 16'b0000000000010001;
        weights1[15986] <= 16'b1111111111111101;
        weights1[15987] <= 16'b1111111111111100;
        weights1[15988] <= 16'b0000000000000101;
        weights1[15989] <= 16'b0000000000000010;
        weights1[15990] <= 16'b0000000000001001;
        weights1[15991] <= 16'b0000000000001000;
        weights1[15992] <= 16'b0000000000100001;
        weights1[15993] <= 16'b0000000000010100;
        weights1[15994] <= 16'b0000000000011011;
        weights1[15995] <= 16'b0000000000011101;
        weights1[15996] <= 16'b0000000000100001;
        weights1[15997] <= 16'b0000000000001100;
        weights1[15998] <= 16'b0000000000001001;
        weights1[15999] <= 16'b0000000000010101;
        weights1[16000] <= 16'b0000000000100001;
        weights1[16001] <= 16'b0000000000010011;
        weights1[16002] <= 16'b1111111111111110;
        weights1[16003] <= 16'b1111111111111110;
        weights1[16004] <= 16'b1111111111111011;
        weights1[16005] <= 16'b1111111111110001;
        weights1[16006] <= 16'b0000000000000011;
        weights1[16007] <= 16'b1111111111111111;
        weights1[16008] <= 16'b0000000000000010;
        weights1[16009] <= 16'b0000000000000001;
        weights1[16010] <= 16'b0000000000000010;
        weights1[16011] <= 16'b1111111111100110;
        weights1[16012] <= 16'b1111111111111011;
        weights1[16013] <= 16'b0000000000000001;
        weights1[16014] <= 16'b1111111111111010;
        weights1[16015] <= 16'b1111111111111110;
        weights1[16016] <= 16'b0000000000001011;
        weights1[16017] <= 16'b0000000000001000;
        weights1[16018] <= 16'b0000000000000000;
        weights1[16019] <= 16'b0000000000010011;
        weights1[16020] <= 16'b0000000000000011;
        weights1[16021] <= 16'b0000000000001101;
        weights1[16022] <= 16'b1111111111110110;
        weights1[16023] <= 16'b0000000000011100;
        weights1[16024] <= 16'b0000000000101111;
        weights1[16025] <= 16'b0000000000011110;
        weights1[16026] <= 16'b0000000000101000;
        weights1[16027] <= 16'b0000000000100011;
        weights1[16028] <= 16'b0000000000100101;
        weights1[16029] <= 16'b0000000000101010;
        weights1[16030] <= 16'b0000000000010111;
        weights1[16031] <= 16'b0000000000011001;
        weights1[16032] <= 16'b0000000000001010;
        weights1[16033] <= 16'b0000000000011110;
        weights1[16034] <= 16'b0000000000001001;
        weights1[16035] <= 16'b0000000000001110;
        weights1[16036] <= 16'b1111111111111111;
        weights1[16037] <= 16'b1111111111111111;
        weights1[16038] <= 16'b1111111111111101;
        weights1[16039] <= 16'b0000000000001010;
        weights1[16040] <= 16'b1111111111111101;
        weights1[16041] <= 16'b0000000000000001;
        weights1[16042] <= 16'b0000000000000100;
        weights1[16043] <= 16'b0000000000000110;
        weights1[16044] <= 16'b0000000000010001;
        weights1[16045] <= 16'b0000000000010110;
        weights1[16046] <= 16'b0000000000011010;
        weights1[16047] <= 16'b0000000000011011;
        weights1[16048] <= 16'b0000000000010101;
        weights1[16049] <= 16'b0000000000010011;
        weights1[16050] <= 16'b0000000000000011;
        weights1[16051] <= 16'b0000000000011010;
        weights1[16052] <= 16'b0000000000011000;
        weights1[16053] <= 16'b0000000000100001;
        weights1[16054] <= 16'b0000000000100101;
        weights1[16055] <= 16'b0000000000110000;
        weights1[16056] <= 16'b0000000000101110;
        weights1[16057] <= 16'b0000000000011011;
        weights1[16058] <= 16'b0000000000100010;
        weights1[16059] <= 16'b0000000000011000;
        weights1[16060] <= 16'b0000000000011000;
        weights1[16061] <= 16'b0000000000010110;
        weights1[16062] <= 16'b0000000000010110;
        weights1[16063] <= 16'b0000000000001010;
        weights1[16064] <= 16'b0000000000010111;
        weights1[16065] <= 16'b0000000000010001;
        weights1[16066] <= 16'b0000000000011101;
        weights1[16067] <= 16'b1111111111111010;
        weights1[16068] <= 16'b0000000000001101;
        weights1[16069] <= 16'b0000000000010110;
        weights1[16070] <= 16'b0000000000010011;
        weights1[16071] <= 16'b0000000000010111;
        weights1[16072] <= 16'b0000000000011100;
        weights1[16073] <= 16'b0000000000101100;
        weights1[16074] <= 16'b0000000000010001;
        weights1[16075] <= 16'b0000000000010111;
        weights1[16076] <= 16'b0000000000000011;
        weights1[16077] <= 16'b0000000000001010;
        weights1[16078] <= 16'b0000000000010110;
        weights1[16079] <= 16'b0000000000000111;
        weights1[16080] <= 16'b0000000000011011;
        weights1[16081] <= 16'b0000000000001100;
        weights1[16082] <= 16'b0000000000001110;
        weights1[16083] <= 16'b0000000000100000;
        weights1[16084] <= 16'b0000000000001000;
        weights1[16085] <= 16'b0000000000101001;
        weights1[16086] <= 16'b0000000000011011;
        weights1[16087] <= 16'b0000000000011100;
        weights1[16088] <= 16'b0000000000010110;
        weights1[16089] <= 16'b0000000000000100;
        weights1[16090] <= 16'b0000000000011010;
        weights1[16091] <= 16'b0000000000000110;
        weights1[16092] <= 16'b0000000000000000;
        weights1[16093] <= 16'b0000000000001011;
        weights1[16094] <= 16'b0000000000000110;
        weights1[16095] <= 16'b0000000000010111;
        weights1[16096] <= 16'b0000000000000111;
        weights1[16097] <= 16'b1111111111111100;
        weights1[16098] <= 16'b0000000000001110;
        weights1[16099] <= 16'b0000000000011000;
        weights1[16100] <= 16'b0000000000011100;
        weights1[16101] <= 16'b0000000000011110;
        weights1[16102] <= 16'b0000000000000111;
        weights1[16103] <= 16'b0000000000001110;
        weights1[16104] <= 16'b0000000000001000;
        weights1[16105] <= 16'b0000000000001001;
        weights1[16106] <= 16'b0000000000010110;
        weights1[16107] <= 16'b1111111111111100;
        weights1[16108] <= 16'b0000000000010001;
        weights1[16109] <= 16'b0000000000000011;
        weights1[16110] <= 16'b0000000000000100;
        weights1[16111] <= 16'b0000000000001001;
        weights1[16112] <= 16'b0000000000001011;
        weights1[16113] <= 16'b0000000000000100;
        weights1[16114] <= 16'b0000000000001100;
        weights1[16115] <= 16'b0000000000010010;
        weights1[16116] <= 16'b0000000000001000;
        weights1[16117] <= 16'b0000000000000100;
        weights1[16118] <= 16'b0000000000010001;
        weights1[16119] <= 16'b0000000000001001;
        weights1[16120] <= 16'b0000000000010100;
        weights1[16121] <= 16'b0000000000000010;
        weights1[16122] <= 16'b0000000000001111;
        weights1[16123] <= 16'b0000000000000011;
        weights1[16124] <= 16'b0000000000001011;
        weights1[16125] <= 16'b1111111111111111;
        weights1[16126] <= 16'b0000000000001110;
        weights1[16127] <= 16'b0000000000001110;
        weights1[16128] <= 16'b0000000000100000;
        weights1[16129] <= 16'b0000000000100100;
        weights1[16130] <= 16'b0000000000001000;
        weights1[16131] <= 16'b0000000000001011;
        weights1[16132] <= 16'b0000000000000111;
        weights1[16133] <= 16'b1111111111110101;
        weights1[16134] <= 16'b0000000000010000;
        weights1[16135] <= 16'b0000000000010011;
        weights1[16136] <= 16'b1111111111110110;
        weights1[16137] <= 16'b0000000000000101;
        weights1[16138] <= 16'b1111111111101001;
        weights1[16139] <= 16'b1111111111110110;
        weights1[16140] <= 16'b1111111111111001;
        weights1[16141] <= 16'b1111111111111101;
        weights1[16142] <= 16'b0000000000000000;
        weights1[16143] <= 16'b0000000000001011;
        weights1[16144] <= 16'b1111111111110000;
        weights1[16145] <= 16'b1111111111111111;
        weights1[16146] <= 16'b1111111111111111;
        weights1[16147] <= 16'b1111111111110001;
        weights1[16148] <= 16'b1111111111111111;
        weights1[16149] <= 16'b0000000000000101;
        weights1[16150] <= 16'b1111111111111100;
        weights1[16151] <= 16'b0000000000010000;
        weights1[16152] <= 16'b0000000000010111;
        weights1[16153] <= 16'b0000000000011000;
        weights1[16154] <= 16'b0000000000011110;
        weights1[16155] <= 16'b0000000000001100;
        weights1[16156] <= 16'b0000000000000111;
        weights1[16157] <= 16'b0000000000011000;
        weights1[16158] <= 16'b0000000000001001;
        weights1[16159] <= 16'b0000000000001010;
        weights1[16160] <= 16'b0000000000000101;
        weights1[16161] <= 16'b0000000000011011;
        weights1[16162] <= 16'b0000000000001111;
        weights1[16163] <= 16'b0000000000000001;
        weights1[16164] <= 16'b0000000000000001;
        weights1[16165] <= 16'b1111111111111010;
        weights1[16166] <= 16'b1111111111111101;
        weights1[16167] <= 16'b1111111111100101;
        weights1[16168] <= 16'b0000000000000010;
        weights1[16169] <= 16'b1111111111110111;
        weights1[16170] <= 16'b1111111111101010;
        weights1[16171] <= 16'b1111111111100101;
        weights1[16172] <= 16'b1111111111101010;
        weights1[16173] <= 16'b1111111111101110;
        weights1[16174] <= 16'b0000000000000100;
        weights1[16175] <= 16'b1111111111110010;
        weights1[16176] <= 16'b0000000000001001;
        weights1[16177] <= 16'b0000000000011001;
        weights1[16178] <= 16'b0000000000010111;
        weights1[16179] <= 16'b0000000000000011;
        weights1[16180] <= 16'b0000000000011011;
        weights1[16181] <= 16'b0000000000010000;
        weights1[16182] <= 16'b0000000000100010;
        weights1[16183] <= 16'b0000000000000010;
        weights1[16184] <= 16'b1111111111110101;
        weights1[16185] <= 16'b0000000000001110;
        weights1[16186] <= 16'b0000000000011001;
        weights1[16187] <= 16'b0000000000001000;
        weights1[16188] <= 16'b0000000000011001;
        weights1[16189] <= 16'b0000000000000110;
        weights1[16190] <= 16'b1111111111110101;
        weights1[16191] <= 16'b0000000000001100;
        weights1[16192] <= 16'b0000000000000001;
        weights1[16193] <= 16'b1111111111111111;
        weights1[16194] <= 16'b1111111111110100;
        weights1[16195] <= 16'b1111111111100100;
        weights1[16196] <= 16'b0000000000001001;
        weights1[16197] <= 16'b1111111111110001;
        weights1[16198] <= 16'b1111111111100100;
        weights1[16199] <= 16'b1111111111111110;
        weights1[16200] <= 16'b1111111111110111;
        weights1[16201] <= 16'b1111111111111001;
        weights1[16202] <= 16'b0000000000000101;
        weights1[16203] <= 16'b0000000000000111;
        weights1[16204] <= 16'b0000000000000101;
        weights1[16205] <= 16'b0000000000001100;
        weights1[16206] <= 16'b0000000000010100;
        weights1[16207] <= 16'b0000000000010011;
        weights1[16208] <= 16'b0000000000001010;
        weights1[16209] <= 16'b0000000000010111;
        weights1[16210] <= 16'b0000000000010101;
        weights1[16211] <= 16'b0000000000000000;
        weights1[16212] <= 16'b1111111111110010;
        weights1[16213] <= 16'b0000000000000111;
        weights1[16214] <= 16'b0000000000001110;
        weights1[16215] <= 16'b0000000000001010;
        weights1[16216] <= 16'b0000000000001100;
        weights1[16217] <= 16'b0000000000000100;
        weights1[16218] <= 16'b0000000000000011;
        weights1[16219] <= 16'b1111111111111111;
        weights1[16220] <= 16'b1111111111110111;
        weights1[16221] <= 16'b1111111111111111;
        weights1[16222] <= 16'b0000000000000111;
        weights1[16223] <= 16'b0000000000010001;
        weights1[16224] <= 16'b0000000000001001;
        weights1[16225] <= 16'b0000000000001100;
        weights1[16226] <= 16'b1111111111111111;
        weights1[16227] <= 16'b0000000000000110;
        weights1[16228] <= 16'b1111111111111111;
        weights1[16229] <= 16'b0000000000000000;
        weights1[16230] <= 16'b0000000000010001;
        weights1[16231] <= 16'b0000000000000111;
        weights1[16232] <= 16'b0000000000000111;
        weights1[16233] <= 16'b0000000000000011;
        weights1[16234] <= 16'b0000000000001001;
        weights1[16235] <= 16'b1111111111111000;
        weights1[16236] <= 16'b0000000000000110;
        weights1[16237] <= 16'b0000000000000001;
        weights1[16238] <= 16'b0000000000000111;
        weights1[16239] <= 16'b0000000000000101;
        weights1[16240] <= 16'b1111111111101111;
        weights1[16241] <= 16'b0000000000000000;
        weights1[16242] <= 16'b0000000000000110;
        weights1[16243] <= 16'b1111111111111010;
        weights1[16244] <= 16'b1111111111111100;
        weights1[16245] <= 16'b0000000000001010;
        weights1[16246] <= 16'b1111111111111011;
        weights1[16247] <= 16'b0000000000000100;
        weights1[16248] <= 16'b0000000000001111;
        weights1[16249] <= 16'b0000000000000110;
        weights1[16250] <= 16'b0000000000000011;
        weights1[16251] <= 16'b0000000000000110;
        weights1[16252] <= 16'b0000000000010101;
        weights1[16253] <= 16'b0000000000010001;
        weights1[16254] <= 16'b0000000000000101;
        weights1[16255] <= 16'b0000000000001000;
        weights1[16256] <= 16'b0000000000010001;
        weights1[16257] <= 16'b0000000000000011;
        weights1[16258] <= 16'b0000000000010001;
        weights1[16259] <= 16'b1111111111111011;
        weights1[16260] <= 16'b0000000000010010;
        weights1[16261] <= 16'b0000000000011000;
        weights1[16262] <= 16'b0000000000001000;
        weights1[16263] <= 16'b0000000000001010;
        weights1[16264] <= 16'b1111111111110111;
        weights1[16265] <= 16'b1111111111110101;
        weights1[16266] <= 16'b1111111111111100;
        weights1[16267] <= 16'b0000000000000101;
        weights1[16268] <= 16'b1111111111110001;
        weights1[16269] <= 16'b1111111111101111;
        weights1[16270] <= 16'b1111111111101100;
        weights1[16271] <= 16'b1111111111111001;
        weights1[16272] <= 16'b1111111111101011;
        weights1[16273] <= 16'b0000000000001111;
        weights1[16274] <= 16'b0000000000000011;
        weights1[16275] <= 16'b0000000000000011;
        weights1[16276] <= 16'b0000000000000110;
        weights1[16277] <= 16'b0000000000000101;
        weights1[16278] <= 16'b0000000000010110;
        weights1[16279] <= 16'b0000000000000010;
        weights1[16280] <= 16'b1111111111111101;
        weights1[16281] <= 16'b0000000000001010;
        weights1[16282] <= 16'b0000000000001100;
        weights1[16283] <= 16'b0000000000010110;
        weights1[16284] <= 16'b0000000000001000;
        weights1[16285] <= 16'b0000000000000011;
        weights1[16286] <= 16'b0000000000010110;
        weights1[16287] <= 16'b1111111111111000;
        weights1[16288] <= 16'b0000000000000001;
        weights1[16289] <= 16'b0000000000000000;
        weights1[16290] <= 16'b1111111111110111;
        weights1[16291] <= 16'b0000000000000001;
        weights1[16292] <= 16'b1111111111111110;
        weights1[16293] <= 16'b1111111111111010;
        weights1[16294] <= 16'b1111111111110111;
        weights1[16295] <= 16'b0000000000000001;
        weights1[16296] <= 16'b1111111111111000;
        weights1[16297] <= 16'b1111111111110000;
        weights1[16298] <= 16'b1111111111101001;
        weights1[16299] <= 16'b1111111111110110;
        weights1[16300] <= 16'b1111111111110001;
        weights1[16301] <= 16'b1111111111101111;
        weights1[16302] <= 16'b1111111111110101;
        weights1[16303] <= 16'b1111111111110101;
        weights1[16304] <= 16'b1111111111111001;
        weights1[16305] <= 16'b1111111111110110;
        weights1[16306] <= 16'b1111111111101111;
        weights1[16307] <= 16'b1111111111101001;
        weights1[16308] <= 16'b0000000000000110;
        weights1[16309] <= 16'b0000000000001100;
        weights1[16310] <= 16'b1111111111110111;
        weights1[16311] <= 16'b1111111111111101;
        weights1[16312] <= 16'b1111111111111000;
        weights1[16313] <= 16'b0000000000000111;
        weights1[16314] <= 16'b0000000000001001;
        weights1[16315] <= 16'b1111111111111111;
        weights1[16316] <= 16'b0000000000000001;
        weights1[16317] <= 16'b0000000000001001;
        weights1[16318] <= 16'b0000000000000100;
        weights1[16319] <= 16'b1111111111110000;
        weights1[16320] <= 16'b1111111111111000;
        weights1[16321] <= 16'b1111111111110111;
        weights1[16322] <= 16'b1111111111110011;
        weights1[16323] <= 16'b1111111111111000;
        weights1[16324] <= 16'b1111111111110101;
        weights1[16325] <= 16'b1111111111100111;
        weights1[16326] <= 16'b1111111111100100;
        weights1[16327] <= 16'b1111111111100111;
        weights1[16328] <= 16'b1111111111110001;
        weights1[16329] <= 16'b1111111111110010;
        weights1[16330] <= 16'b1111111111100000;
        weights1[16331] <= 16'b1111111111101010;
        weights1[16332] <= 16'b1111111111110101;
        weights1[16333] <= 16'b1111111111110100;
        weights1[16334] <= 16'b1111111111111011;
        weights1[16335] <= 16'b1111111111110000;
        weights1[16336] <= 16'b1111111111101111;
        weights1[16337] <= 16'b1111111111111100;
        weights1[16338] <= 16'b1111111111111101;
        weights1[16339] <= 16'b1111111111111001;
        weights1[16340] <= 16'b0000000000000001;
        weights1[16341] <= 16'b1111111111111010;
        weights1[16342] <= 16'b0000000000000000;
        weights1[16343] <= 16'b1111111111101111;
        weights1[16344] <= 16'b1111111111111001;
        weights1[16345] <= 16'b1111111111101101;
        weights1[16346] <= 16'b1111111111101010;
        weights1[16347] <= 16'b1111111111101011;
        weights1[16348] <= 16'b1111111111111110;
        weights1[16349] <= 16'b0000000000000001;
        weights1[16350] <= 16'b1111111111110111;
        weights1[16351] <= 16'b0000000000000011;
        weights1[16352] <= 16'b1111111111110110;
        weights1[16353] <= 16'b1111111111100111;
        weights1[16354] <= 16'b1111111111110001;
        weights1[16355] <= 16'b1111111111111000;
        weights1[16356] <= 16'b1111111111011110;
        weights1[16357] <= 16'b1111111111100001;
        weights1[16358] <= 16'b1111111111101101;
        weights1[16359] <= 16'b1111111111100101;
        weights1[16360] <= 16'b1111111111110001;
        weights1[16361] <= 16'b0000000000001010;
        weights1[16362] <= 16'b1111111111110110;
        weights1[16363] <= 16'b1111111111111001;
        weights1[16364] <= 16'b0000000000000001;
        weights1[16365] <= 16'b1111111111111110;
        weights1[16366] <= 16'b1111111111110101;
        weights1[16367] <= 16'b1111111111101011;
        weights1[16368] <= 16'b1111111111111100;
        weights1[16369] <= 16'b1111111111111111;
        weights1[16370] <= 16'b1111111111111000;
        weights1[16371] <= 16'b1111111111111001;
        weights1[16372] <= 16'b1111111111110010;
        weights1[16373] <= 16'b1111111111110010;
        weights1[16374] <= 16'b1111111111111000;
        weights1[16375] <= 16'b1111111111101110;
        weights1[16376] <= 16'b0000000000001001;
        weights1[16377] <= 16'b0000000000001010;
        weights1[16378] <= 16'b1111111111111111;
        weights1[16379] <= 16'b0000000000000110;
        weights1[16380] <= 16'b0000000000000011;
        weights1[16381] <= 16'b1111111111110011;
        weights1[16382] <= 16'b1111111111110110;
        weights1[16383] <= 16'b1111111111111001;
        weights1[16384] <= 16'b1111111111110111;
        weights1[16385] <= 16'b1111111111100010;
        weights1[16386] <= 16'b1111111111100111;
        weights1[16387] <= 16'b1111111111101001;
        weights1[16388] <= 16'b1111111111011011;
        weights1[16389] <= 16'b1111111111100000;
        weights1[16390] <= 16'b1111111111101101;
        weights1[16391] <= 16'b1111111111101000;
        weights1[16392] <= 16'b1111111111100001;
        weights1[16393] <= 16'b1111111111101100;
        weights1[16394] <= 16'b1111111111110101;
        weights1[16395] <= 16'b1111111111101011;
        weights1[16396] <= 16'b1111111111101010;
        weights1[16397] <= 16'b1111111111111000;
        weights1[16398] <= 16'b1111111111011101;
        weights1[16399] <= 16'b1111111111011011;
        weights1[16400] <= 16'b1111111111110010;
        weights1[16401] <= 16'b1111111111111000;
        weights1[16402] <= 16'b1111111111111001;
        weights1[16403] <= 16'b1111111111110000;
        weights1[16404] <= 16'b0000000000010010;
        weights1[16405] <= 16'b0000000000010000;
        weights1[16406] <= 16'b0000000000000000;
        weights1[16407] <= 16'b0000000000001010;
        weights1[16408] <= 16'b0000000000000100;
        weights1[16409] <= 16'b0000000000000001;
        weights1[16410] <= 16'b0000000000000111;
        weights1[16411] <= 16'b0000000000001011;
        weights1[16412] <= 16'b1111111111111110;
        weights1[16413] <= 16'b1111111111111110;
        weights1[16414] <= 16'b1111111111111011;
        weights1[16415] <= 16'b1111111111111111;
        weights1[16416] <= 16'b1111111111110011;
        weights1[16417] <= 16'b1111111111110100;
        weights1[16418] <= 16'b1111111111101100;
        weights1[16419] <= 16'b1111111111101100;
        weights1[16420] <= 16'b1111111111101100;
        weights1[16421] <= 16'b1111111111010101;
        weights1[16422] <= 16'b1111111111100111;
        weights1[16423] <= 16'b1111111111101010;
        weights1[16424] <= 16'b1111111111010110;
        weights1[16425] <= 16'b1111111111101110;
        weights1[16426] <= 16'b1111111111110110;
        weights1[16427] <= 16'b1111111111100110;
        weights1[16428] <= 16'b1111111111101101;
        weights1[16429] <= 16'b0000000000000100;
        weights1[16430] <= 16'b0000000000001001;
        weights1[16431] <= 16'b0000000000010011;
        weights1[16432] <= 16'b0000000000010110;
        weights1[16433] <= 16'b0000000000011000;
        weights1[16434] <= 16'b0000000000001110;
        weights1[16435] <= 16'b0000000000001010;
        weights1[16436] <= 16'b0000000000000100;
        weights1[16437] <= 16'b0000000000000100;
        weights1[16438] <= 16'b0000000000000110;
        weights1[16439] <= 16'b0000000000000100;
        weights1[16440] <= 16'b0000000000001000;
        weights1[16441] <= 16'b0000000000010010;
        weights1[16442] <= 16'b0000000000011100;
        weights1[16443] <= 16'b0000000000010010;
        weights1[16444] <= 16'b0000000000010101;
        weights1[16445] <= 16'b0000000000001110;
        weights1[16446] <= 16'b0000000000001100;
        weights1[16447] <= 16'b0000000000001111;
        weights1[16448] <= 16'b0000000000010010;
        weights1[16449] <= 16'b0000000000011011;
        weights1[16450] <= 16'b0000000000010001;
        weights1[16451] <= 16'b0000000000001101;
        weights1[16452] <= 16'b0000000000011101;
        weights1[16453] <= 16'b0000000000011001;
        weights1[16454] <= 16'b0000000000011011;
        weights1[16455] <= 16'b0000000000010101;
        weights1[16456] <= 16'b0000000000100010;
        weights1[16457] <= 16'b0000000000100001;
        weights1[16458] <= 16'b0000000000010101;
        weights1[16459] <= 16'b0000000000011000;
        weights1[16460] <= 16'b0000000000011110;
        weights1[16461] <= 16'b0000000000011011;
        weights1[16462] <= 16'b0000000000010111;
        weights1[16463] <= 16'b0000000000000110;
        weights1[16464] <= 16'b0000000000000000;
        weights1[16465] <= 16'b1111111111111111;
        weights1[16466] <= 16'b1111111111111111;
        weights1[16467] <= 16'b1111111111111111;
        weights1[16468] <= 16'b1111111111111111;
        weights1[16469] <= 16'b1111111111111111;
        weights1[16470] <= 16'b1111111111110111;
        weights1[16471] <= 16'b1111111111111000;
        weights1[16472] <= 16'b1111111111101100;
        weights1[16473] <= 16'b1111111111101010;
        weights1[16474] <= 16'b1111111111100101;
        weights1[16475] <= 16'b1111111111100000;
        weights1[16476] <= 16'b1111111111100011;
        weights1[16477] <= 16'b1111111111101100;
        weights1[16478] <= 16'b1111111111111010;
        weights1[16479] <= 16'b1111111111111110;
        weights1[16480] <= 16'b0000000000001001;
        weights1[16481] <= 16'b0000000000001010;
        weights1[16482] <= 16'b0000000000000100;
        weights1[16483] <= 16'b1111111111111110;
        weights1[16484] <= 16'b0000000000000110;
        weights1[16485] <= 16'b0000000000000100;
        weights1[16486] <= 16'b0000000000001100;
        weights1[16487] <= 16'b0000000000001010;
        weights1[16488] <= 16'b0000000000000100;
        weights1[16489] <= 16'b0000000000000010;
        weights1[16490] <= 16'b1111111111111110;
        weights1[16491] <= 16'b0000000000000011;
        weights1[16492] <= 16'b0000000000000000;
        weights1[16493] <= 16'b1111111111111111;
        weights1[16494] <= 16'b0000000000000000;
        weights1[16495] <= 16'b0000000000000000;
        weights1[16496] <= 16'b1111111111111110;
        weights1[16497] <= 16'b1111111111111010;
        weights1[16498] <= 16'b1111111111110000;
        weights1[16499] <= 16'b1111111111110011;
        weights1[16500] <= 16'b1111111111110000;
        weights1[16501] <= 16'b1111111111101001;
        weights1[16502] <= 16'b1111111111100010;
        weights1[16503] <= 16'b1111111111011011;
        weights1[16504] <= 16'b1111111111010100;
        weights1[16505] <= 16'b1111111111010101;
        weights1[16506] <= 16'b1111111111111001;
        weights1[16507] <= 16'b0000000000001011;
        weights1[16508] <= 16'b0000000000000011;
        weights1[16509] <= 16'b0000000000000011;
        weights1[16510] <= 16'b1111111111111001;
        weights1[16511] <= 16'b1111111111111101;
        weights1[16512] <= 16'b0000000000000111;
        weights1[16513] <= 16'b0000000000001100;
        weights1[16514] <= 16'b0000000000010011;
        weights1[16515] <= 16'b1111111111111111;
        weights1[16516] <= 16'b0000000000000010;
        weights1[16517] <= 16'b1111111111111101;
        weights1[16518] <= 16'b1111111111111111;
        weights1[16519] <= 16'b1111111111111110;
        weights1[16520] <= 16'b1111111111111111;
        weights1[16521] <= 16'b0000000000000001;
        weights1[16522] <= 16'b1111111111111111;
        weights1[16523] <= 16'b1111111111111101;
        weights1[16524] <= 16'b1111111111110011;
        weights1[16525] <= 16'b1111111111110010;
        weights1[16526] <= 16'b1111111111101101;
        weights1[16527] <= 16'b1111111111111000;
        weights1[16528] <= 16'b1111111111110001;
        weights1[16529] <= 16'b1111111111101010;
        weights1[16530] <= 16'b1111111111010101;
        weights1[16531] <= 16'b1111111111001110;
        weights1[16532] <= 16'b1111111111011011;
        weights1[16533] <= 16'b1111111111101101;
        weights1[16534] <= 16'b1111111111111010;
        weights1[16535] <= 16'b0000000000001110;
        weights1[16536] <= 16'b0000000000001111;
        weights1[16537] <= 16'b1111111111110000;
        weights1[16538] <= 16'b0000000000000110;
        weights1[16539] <= 16'b1111111111111101;
        weights1[16540] <= 16'b1111111111111110;
        weights1[16541] <= 16'b0000000000000100;
        weights1[16542] <= 16'b0000000000000000;
        weights1[16543] <= 16'b1111111111111101;
        weights1[16544] <= 16'b1111111111111111;
        weights1[16545] <= 16'b1111111111111110;
        weights1[16546] <= 16'b1111111111111011;
        weights1[16547] <= 16'b1111111111111101;
        weights1[16548] <= 16'b1111111111111111;
        weights1[16549] <= 16'b1111111111111111;
        weights1[16550] <= 16'b1111111111111011;
        weights1[16551] <= 16'b1111111111110001;
        weights1[16552] <= 16'b1111111111101110;
        weights1[16553] <= 16'b1111111111101111;
        weights1[16554] <= 16'b1111111111111001;
        weights1[16555] <= 16'b1111111111110101;
        weights1[16556] <= 16'b1111111111101011;
        weights1[16557] <= 16'b1111111111111011;
        weights1[16558] <= 16'b1111111111110001;
        weights1[16559] <= 16'b1111111111110101;
        weights1[16560] <= 16'b1111111111100000;
        weights1[16561] <= 16'b1111111111110100;
        weights1[16562] <= 16'b1111111111100011;
        weights1[16563] <= 16'b1111111111110010;
        weights1[16564] <= 16'b0000000000000010;
        weights1[16565] <= 16'b1111111111101011;
        weights1[16566] <= 16'b1111111111110011;
        weights1[16567] <= 16'b1111111111111001;
        weights1[16568] <= 16'b1111111111101111;
        weights1[16569] <= 16'b1111111111110000;
        weights1[16570] <= 16'b1111111111110010;
        weights1[16571] <= 16'b0000000000000011;
        weights1[16572] <= 16'b1111111111111010;
        weights1[16573] <= 16'b1111111111110000;
        weights1[16574] <= 16'b1111111111110000;
        weights1[16575] <= 16'b0000000000000000;
        weights1[16576] <= 16'b0000000000000000;
        weights1[16577] <= 16'b0000000000000010;
        weights1[16578] <= 16'b1111111111111100;
        weights1[16579] <= 16'b1111111111110000;
        weights1[16580] <= 16'b1111111111101101;
        weights1[16581] <= 16'b1111111111111000;
        weights1[16582] <= 16'b0000000000001011;
        weights1[16583] <= 16'b0000000000000111;
        weights1[16584] <= 16'b0000000000010100;
        weights1[16585] <= 16'b0000000000000000;
        weights1[16586] <= 16'b1111111111101000;
        weights1[16587] <= 16'b1111111111110100;
        weights1[16588] <= 16'b1111111111111111;
        weights1[16589] <= 16'b1111111111110101;
        weights1[16590] <= 16'b0000000000011000;
        weights1[16591] <= 16'b0000000000000111;
        weights1[16592] <= 16'b0000000000001110;
        weights1[16593] <= 16'b0000000000001100;
        weights1[16594] <= 16'b0000000000001111;
        weights1[16595] <= 16'b0000000000000010;
        weights1[16596] <= 16'b0000000000000110;
        weights1[16597] <= 16'b0000000000000000;
        weights1[16598] <= 16'b1111111111101110;
        weights1[16599] <= 16'b0000000000000101;
        weights1[16600] <= 16'b1111111111111101;
        weights1[16601] <= 16'b1111111111100001;
        weights1[16602] <= 16'b1111111111111001;
        weights1[16603] <= 16'b1111111111110111;
        weights1[16604] <= 16'b0000000000000001;
        weights1[16605] <= 16'b1111111111111011;
        weights1[16606] <= 16'b1111111111110110;
        weights1[16607] <= 16'b1111111111101100;
        weights1[16608] <= 16'b1111111111110111;
        weights1[16609] <= 16'b1111111111110101;
        weights1[16610] <= 16'b0000000000010110;
        weights1[16611] <= 16'b0000000000001011;
        weights1[16612] <= 16'b0000000000100100;
        weights1[16613] <= 16'b0000000000011111;
        weights1[16614] <= 16'b1111111111111100;
        weights1[16615] <= 16'b0000000000010001;
        weights1[16616] <= 16'b1111111111111100;
        weights1[16617] <= 16'b1111111111110011;
        weights1[16618] <= 16'b0000000000010001;
        weights1[16619] <= 16'b1111111111110100;
        weights1[16620] <= 16'b1111111111111010;
        weights1[16621] <= 16'b0000000000000011;
        weights1[16622] <= 16'b0000000000000111;
        weights1[16623] <= 16'b1111111111110001;
        weights1[16624] <= 16'b1111111111111011;
        weights1[16625] <= 16'b0000000000001111;
        weights1[16626] <= 16'b0000000000000001;
        weights1[16627] <= 16'b0000000000010001;
        weights1[16628] <= 16'b0000000000001000;
        weights1[16629] <= 16'b1111111111110011;
        weights1[16630] <= 16'b1111111111111000;
        weights1[16631] <= 16'b1111111111101111;
        weights1[16632] <= 16'b0000000000000010;
        weights1[16633] <= 16'b0000000000000010;
        weights1[16634] <= 16'b0000000000000001;
        weights1[16635] <= 16'b1111111111110000;
        weights1[16636] <= 16'b1111111111111101;
        weights1[16637] <= 16'b0000000000001010;
        weights1[16638] <= 16'b1111111111111001;
        weights1[16639] <= 16'b0000000000010000;
        weights1[16640] <= 16'b0000000000010100;
        weights1[16641] <= 16'b0000000000101111;
        weights1[16642] <= 16'b0000000000000100;
        weights1[16643] <= 16'b1111111111110001;
        weights1[16644] <= 16'b0000000000001001;
        weights1[16645] <= 16'b1111111111111001;
        weights1[16646] <= 16'b1111111111111000;
        weights1[16647] <= 16'b0000000000001101;
        weights1[16648] <= 16'b0000000000001110;
        weights1[16649] <= 16'b0000000000010001;
        weights1[16650] <= 16'b1111111111111101;
        weights1[16651] <= 16'b0000000000000011;
        weights1[16652] <= 16'b1111111111111110;
        weights1[16653] <= 16'b1111111111111100;
        weights1[16654] <= 16'b0000000000010010;
        weights1[16655] <= 16'b1111111111111000;
        weights1[16656] <= 16'b1111111111111100;
        weights1[16657] <= 16'b0000000000000001;
        weights1[16658] <= 16'b0000000000001001;
        weights1[16659] <= 16'b0000000000000100;
        weights1[16660] <= 16'b0000000000000001;
        weights1[16661] <= 16'b0000000000000011;
        weights1[16662] <= 16'b0000000000000101;
        weights1[16663] <= 16'b1111111111111111;
        weights1[16664] <= 16'b1111111111111010;
        weights1[16665] <= 16'b1111111111111110;
        weights1[16666] <= 16'b0000000000000111;
        weights1[16667] <= 16'b0000000000000010;
        weights1[16668] <= 16'b1111111111111010;
        weights1[16669] <= 16'b0000000000011010;
        weights1[16670] <= 16'b0000000000011101;
        weights1[16671] <= 16'b0000000000010100;
        weights1[16672] <= 16'b1111111111111100;
        weights1[16673] <= 16'b0000000000010001;
        weights1[16674] <= 16'b1111111111100100;
        weights1[16675] <= 16'b0000000000001000;
        weights1[16676] <= 16'b1111111111111111;
        weights1[16677] <= 16'b1111111111111000;
        weights1[16678] <= 16'b0000000000010100;
        weights1[16679] <= 16'b0000000000100010;
        weights1[16680] <= 16'b0000000000000001;
        weights1[16681] <= 16'b1111111111101110;
        weights1[16682] <= 16'b0000000000001101;
        weights1[16683] <= 16'b1111111111111000;
        weights1[16684] <= 16'b0000000000010011;
        weights1[16685] <= 16'b0000000000001110;
        weights1[16686] <= 16'b0000000000000001;
        weights1[16687] <= 16'b0000000000000100;
        weights1[16688] <= 16'b0000000000000010;
        weights1[16689] <= 16'b0000000000000011;
        weights1[16690] <= 16'b1111111111111110;
        weights1[16691] <= 16'b1111111111111111;
        weights1[16692] <= 16'b1111111111111010;
        weights1[16693] <= 16'b0000000000011010;
        weights1[16694] <= 16'b1111111111110100;
        weights1[16695] <= 16'b1111111111101100;
        weights1[16696] <= 16'b0000000000001000;
        weights1[16697] <= 16'b0000000000011110;
        weights1[16698] <= 16'b0000000000011010;
        weights1[16699] <= 16'b0000000000010000;
        weights1[16700] <= 16'b0000000000010000;
        weights1[16701] <= 16'b0000000000000011;
        weights1[16702] <= 16'b0000000000000011;
        weights1[16703] <= 16'b1111111111111111;
        weights1[16704] <= 16'b0000000000000001;
        weights1[16705] <= 16'b0000000000001101;
        weights1[16706] <= 16'b0000000000000101;
        weights1[16707] <= 16'b0000000000000100;
        weights1[16708] <= 16'b0000000000001001;
        weights1[16709] <= 16'b1111111111111110;
        weights1[16710] <= 16'b0000000000000110;
        weights1[16711] <= 16'b0000000000000010;
        weights1[16712] <= 16'b1111111111110000;
        weights1[16713] <= 16'b1111111111111001;
        weights1[16714] <= 16'b0000000000001000;
        weights1[16715] <= 16'b0000000000000101;
        weights1[16716] <= 16'b1111111111111111;
        weights1[16717] <= 16'b0000000000000010;
        weights1[16718] <= 16'b0000000000001110;
        weights1[16719] <= 16'b1111111111111101;
        weights1[16720] <= 16'b0000000000000110;
        weights1[16721] <= 16'b0000000000010011;
        weights1[16722] <= 16'b0000000000011011;
        weights1[16723] <= 16'b0000000000100010;
        weights1[16724] <= 16'b0000000000011001;
        weights1[16725] <= 16'b0000000000000111;
        weights1[16726] <= 16'b0000000000000000;
        weights1[16727] <= 16'b0000000000101000;
        weights1[16728] <= 16'b0000000000010101;
        weights1[16729] <= 16'b0000000000000011;
        weights1[16730] <= 16'b1111111110011011;
        weights1[16731] <= 16'b1111111111101000;
        weights1[16732] <= 16'b1111111111111010;
        weights1[16733] <= 16'b1111111111111101;
        weights1[16734] <= 16'b0000000000001001;
        weights1[16735] <= 16'b0000000000000101;
        weights1[16736] <= 16'b1111111111111101;
        weights1[16737] <= 16'b1111111111111111;
        weights1[16738] <= 16'b1111111111111001;
        weights1[16739] <= 16'b1111111111110011;
        weights1[16740] <= 16'b1111111111111110;
        weights1[16741] <= 16'b1111111111111110;
        weights1[16742] <= 16'b1111111111110110;
        weights1[16743] <= 16'b1111111111110101;
        weights1[16744] <= 16'b0000000000000000;
        weights1[16745] <= 16'b0000000000000100;
        weights1[16746] <= 16'b0000000000001001;
        weights1[16747] <= 16'b0000000000001000;
        weights1[16748] <= 16'b1111111111110000;
        weights1[16749] <= 16'b0000000000000010;
        weights1[16750] <= 16'b0000000000000011;
        weights1[16751] <= 16'b1111111111101111;
        weights1[16752] <= 16'b0000000000100011;
        weights1[16753] <= 16'b0000000000010010;
        weights1[16754] <= 16'b0000000000011100;
        weights1[16755] <= 16'b1111111111101001;
        weights1[16756] <= 16'b0000000000001001;
        weights1[16757] <= 16'b1111111110001100;
        weights1[16758] <= 16'b1111111101100111;
        weights1[16759] <= 16'b1111111111010000;
        weights1[16760] <= 16'b1111111111111001;
        weights1[16761] <= 16'b0000000000001101;
        weights1[16762] <= 16'b1111111111111111;
        weights1[16763] <= 16'b1111111111110000;
        weights1[16764] <= 16'b1111111111110110;
        weights1[16765] <= 16'b1111111111111010;
        weights1[16766] <= 16'b0000000000000001;
        weights1[16767] <= 16'b1111111111110011;
        weights1[16768] <= 16'b1111111111111100;
        weights1[16769] <= 16'b1111111111110111;
        weights1[16770] <= 16'b1111111111101111;
        weights1[16771] <= 16'b1111111111101110;
        weights1[16772] <= 16'b0000000000000000;
        weights1[16773] <= 16'b0000000000001001;
        weights1[16774] <= 16'b0000000000001001;
        weights1[16775] <= 16'b1111111111110110;
        weights1[16776] <= 16'b1111111111110111;
        weights1[16777] <= 16'b1111111111110110;
        weights1[16778] <= 16'b0000000000101100;
        weights1[16779] <= 16'b0000000000000111;
        weights1[16780] <= 16'b0000000000001000;
        weights1[16781] <= 16'b0000000000001111;
        weights1[16782] <= 16'b0000000000010001;
        weights1[16783] <= 16'b0000000000001110;
        weights1[16784] <= 16'b1111111110011110;
        weights1[16785] <= 16'b1111111101000110;
        weights1[16786] <= 16'b1111111111001011;
        weights1[16787] <= 16'b1111111111101010;
        weights1[16788] <= 16'b1111111111110110;
        weights1[16789] <= 16'b0000000000000011;
        weights1[16790] <= 16'b1111111111111110;
        weights1[16791] <= 16'b0000000000001011;
        weights1[16792] <= 16'b1111111111110111;
        weights1[16793] <= 16'b1111111111111001;
        weights1[16794] <= 16'b1111111111111100;
        weights1[16795] <= 16'b0000000000000101;
        weights1[16796] <= 16'b0000000000001000;
        weights1[16797] <= 16'b1111111111110000;
        weights1[16798] <= 16'b1111111111110010;
        weights1[16799] <= 16'b1111111111101010;
        weights1[16800] <= 16'b0000000000000010;
        weights1[16801] <= 16'b0000000000000000;
        weights1[16802] <= 16'b1111111111110111;
        weights1[16803] <= 16'b0000000000000011;
        weights1[16804] <= 16'b1111111111111100;
        weights1[16805] <= 16'b1111111111111110;
        weights1[16806] <= 16'b0000000000000011;
        weights1[16807] <= 16'b0000000000001011;
        weights1[16808] <= 16'b0000000000011010;
        weights1[16809] <= 16'b0000000000001100;
        weights1[16810] <= 16'b1111111111100111;
        weights1[16811] <= 16'b1111111111001111;
        weights1[16812] <= 16'b1111111100110101;
        weights1[16813] <= 16'b1111111110000100;
        weights1[16814] <= 16'b0000000000010000;
        weights1[16815] <= 16'b1111111111111001;
        weights1[16816] <= 16'b0000000000001001;
        weights1[16817] <= 16'b0000000000001010;
        weights1[16818] <= 16'b1111111111110110;
        weights1[16819] <= 16'b0000000000000000;
        weights1[16820] <= 16'b1111111111110111;
        weights1[16821] <= 16'b1111111111110011;
        weights1[16822] <= 16'b1111111111110011;
        weights1[16823] <= 16'b0000000000000011;
        weights1[16824] <= 16'b1111111111101110;
        weights1[16825] <= 16'b1111111111100110;
        weights1[16826] <= 16'b1111111111101110;
        weights1[16827] <= 16'b1111111111101010;
        weights1[16828] <= 16'b1111111111111110;
        weights1[16829] <= 16'b1111111111110110;
        weights1[16830] <= 16'b1111111111111100;
        weights1[16831] <= 16'b1111111111110100;
        weights1[16832] <= 16'b1111111111110011;
        weights1[16833] <= 16'b1111111111110101;
        weights1[16834] <= 16'b0000000000000011;
        weights1[16835] <= 16'b1111111111101001;
        weights1[16836] <= 16'b1111111111110010;
        weights1[16837] <= 16'b1111111111001100;
        weights1[16838] <= 16'b1111111110100001;
        weights1[16839] <= 16'b1111111100101011;
        weights1[16840] <= 16'b1111111101111100;
        weights1[16841] <= 16'b0000000000000010;
        weights1[16842] <= 16'b1111111111011101;
        weights1[16843] <= 16'b1111111111111111;
        weights1[16844] <= 16'b0000000000000011;
        weights1[16845] <= 16'b0000000000001010;
        weights1[16846] <= 16'b1111111111110001;
        weights1[16847] <= 16'b1111111111101000;
        weights1[16848] <= 16'b1111111111110010;
        weights1[16849] <= 16'b1111111111110000;
        weights1[16850] <= 16'b1111111111010110;
        weights1[16851] <= 16'b1111111111011100;
        weights1[16852] <= 16'b1111111111100100;
        weights1[16853] <= 16'b1111111111101101;
        weights1[16854] <= 16'b1111111111101100;
        weights1[16855] <= 16'b1111111111101111;
        weights1[16856] <= 16'b1111111111110101;
        weights1[16857] <= 16'b1111111111110100;
        weights1[16858] <= 16'b1111111111100110;
        weights1[16859] <= 16'b1111111111101100;
        weights1[16860] <= 16'b1111111111010110;
        weights1[16861] <= 16'b1111111111011111;
        weights1[16862] <= 16'b1111111111001101;
        weights1[16863] <= 16'b1111111111001001;
        weights1[16864] <= 16'b1111111101111101;
        weights1[16865] <= 16'b1111111101110000;
        weights1[16866] <= 16'b1111111100110001;
        weights1[16867] <= 16'b1111111110110110;
        weights1[16868] <= 16'b1111111111101000;
        weights1[16869] <= 16'b1111111111110011;
        weights1[16870] <= 16'b1111111111111000;
        weights1[16871] <= 16'b1111111111110110;
        weights1[16872] <= 16'b0000000000000100;
        weights1[16873] <= 16'b0000000000010001;
        weights1[16874] <= 16'b0000000000001101;
        weights1[16875] <= 16'b0000000000000011;
        weights1[16876] <= 16'b1111111111101100;
        weights1[16877] <= 16'b1111111111100110;
        weights1[16878] <= 16'b1111111111101000;
        weights1[16879] <= 16'b1111111111010110;
        weights1[16880] <= 16'b1111111111100100;
        weights1[16881] <= 16'b1111111111100001;
        weights1[16882] <= 16'b1111111111100011;
        weights1[16883] <= 16'b1111111111101100;
        weights1[16884] <= 16'b1111111111101010;
        weights1[16885] <= 16'b1111111111100110;
        weights1[16886] <= 16'b1111111111100010;
        weights1[16887] <= 16'b1111111111001111;
        weights1[16888] <= 16'b1111111110111110;
        weights1[16889] <= 16'b1111111110110011;
        weights1[16890] <= 16'b1111111110010001;
        weights1[16891] <= 16'b1111111101101001;
        weights1[16892] <= 16'b1111111101001110;
        weights1[16893] <= 16'b1111111101010011;
        weights1[16894] <= 16'b1111111111000101;
        weights1[16895] <= 16'b1111111111100101;
        weights1[16896] <= 16'b1111111111110111;
        weights1[16897] <= 16'b1111111111111100;
        weights1[16898] <= 16'b0000000000000001;
        weights1[16899] <= 16'b0000000000000001;
        weights1[16900] <= 16'b0000000000000010;
        weights1[16901] <= 16'b0000000000000100;
        weights1[16902] <= 16'b0000000000010010;
        weights1[16903] <= 16'b0000000000010111;
        weights1[16904] <= 16'b1111111111110001;
        weights1[16905] <= 16'b1111111111101110;
        weights1[16906] <= 16'b1111111111100001;
        weights1[16907] <= 16'b1111111111110100;
        weights1[16908] <= 16'b1111111111101100;
        weights1[16909] <= 16'b1111111111011111;
        weights1[16910] <= 16'b1111111111101010;
        weights1[16911] <= 16'b1111111111101010;
        weights1[16912] <= 16'b1111111111101101;
        weights1[16913] <= 16'b1111111111011101;
        weights1[16914] <= 16'b1111111111010101;
        weights1[16915] <= 16'b1111111111001101;
        weights1[16916] <= 16'b1111111110110001;
        weights1[16917] <= 16'b1111111110100010;
        weights1[16918] <= 16'b1111111101111110;
        weights1[16919] <= 16'b1111111101111000;
        weights1[16920] <= 16'b1111111110010010;
        weights1[16921] <= 16'b1111111111111000;
        weights1[16922] <= 16'b0000000000000001;
        weights1[16923] <= 16'b0000000000001010;
        weights1[16924] <= 16'b0000000000000001;
        weights1[16925] <= 16'b0000000000001001;
        weights1[16926] <= 16'b1111111111111100;
        weights1[16927] <= 16'b0000000000000111;
        weights1[16928] <= 16'b0000000000001111;
        weights1[16929] <= 16'b0000000000011010;
        weights1[16930] <= 16'b0000000000000101;
        weights1[16931] <= 16'b1111111111100111;
        weights1[16932] <= 16'b1111111111011100;
        weights1[16933] <= 16'b1111111111100100;
        weights1[16934] <= 16'b1111111111110010;
        weights1[16935] <= 16'b0000000000000111;
        weights1[16936] <= 16'b0000000000000101;
        weights1[16937] <= 16'b1111111111111100;
        weights1[16938] <= 16'b1111111111110111;
        weights1[16939] <= 16'b1111111111111111;
        weights1[16940] <= 16'b1111111111101001;
        weights1[16941] <= 16'b1111111111011000;
        weights1[16942] <= 16'b1111111111001110;
        weights1[16943] <= 16'b1111111111001010;
        weights1[16944] <= 16'b1111111110110000;
        weights1[16945] <= 16'b1111111110110101;
        weights1[16946] <= 16'b1111111110111011;
        weights1[16947] <= 16'b1111111111010111;
        weights1[16948] <= 16'b0000000000010111;
        weights1[16949] <= 16'b0000000000101010;
        weights1[16950] <= 16'b0000000000000001;
        weights1[16951] <= 16'b0000000000100001;
        weights1[16952] <= 16'b1111111111111100;
        weights1[16953] <= 16'b0000000000000111;
        weights1[16954] <= 16'b1111111111111100;
        weights1[16955] <= 16'b0000000000010101;
        weights1[16956] <= 16'b1111111111111101;
        weights1[16957] <= 16'b1111111111110110;
        weights1[16958] <= 16'b0000000000000011;
        weights1[16959] <= 16'b1111111111101001;
        weights1[16960] <= 16'b1111111111101101;
        weights1[16961] <= 16'b1111111111101100;
        weights1[16962] <= 16'b0000000000000110;
        weights1[16963] <= 16'b0000000000011100;
        weights1[16964] <= 16'b0000000000011110;
        weights1[16965] <= 16'b0000000000000110;
        weights1[16966] <= 16'b0000000000010100;
        weights1[16967] <= 16'b0000000000000110;
        weights1[16968] <= 16'b1111111111100110;
        weights1[16969] <= 16'b1111111111011001;
        weights1[16970] <= 16'b1111111111001110;
        weights1[16971] <= 16'b1111111111001101;
        weights1[16972] <= 16'b1111111111010010;
        weights1[16973] <= 16'b1111111111000100;
        weights1[16974] <= 16'b1111111111101111;
        weights1[16975] <= 16'b0000000000100011;
        weights1[16976] <= 16'b0000000000010101;
        weights1[16977] <= 16'b0000000000000010;
        weights1[16978] <= 16'b0000000000000010;
        weights1[16979] <= 16'b1111111111111011;
        weights1[16980] <= 16'b0000000000000000;
        weights1[16981] <= 16'b0000000000000000;
        weights1[16982] <= 16'b0000000000001101;
        weights1[16983] <= 16'b0000000000000100;
        weights1[16984] <= 16'b0000000000000011;
        weights1[16985] <= 16'b0000000000000011;
        weights1[16986] <= 16'b1111111111111011;
        weights1[16987] <= 16'b1111111111110000;
        weights1[16988] <= 16'b0000000000000001;
        weights1[16989] <= 16'b0000000000011111;
        weights1[16990] <= 16'b1111111111111110;
        weights1[16991] <= 16'b1111111111110001;
        weights1[16992] <= 16'b0000000000001111;
        weights1[16993] <= 16'b0000000000010110;
        weights1[16994] <= 16'b0000000000001111;
        weights1[16995] <= 16'b0000000000001011;
        weights1[16996] <= 16'b1111111111101010;
        weights1[16997] <= 16'b1111111111011010;
        weights1[16998] <= 16'b1111111111010100;
        weights1[16999] <= 16'b1111111111010111;
        weights1[17000] <= 16'b1111111111011011;
        weights1[17001] <= 16'b1111111111101110;
        weights1[17002] <= 16'b1111111111110011;
        weights1[17003] <= 16'b0000000000001100;
        weights1[17004] <= 16'b1111111111110110;
        weights1[17005] <= 16'b0000000000011001;
        weights1[17006] <= 16'b1111111111111000;
        weights1[17007] <= 16'b0000000000011011;
        weights1[17008] <= 16'b0000000000001000;
        weights1[17009] <= 16'b0000000000000001;
        weights1[17010] <= 16'b0000000000000100;
        weights1[17011] <= 16'b1111111111110010;
        weights1[17012] <= 16'b0000000000000111;
        weights1[17013] <= 16'b1111111111101111;
        weights1[17014] <= 16'b1111111111101001;
        weights1[17015] <= 16'b0000000000001010;
        weights1[17016] <= 16'b0000000000001000;
        weights1[17017] <= 16'b1111111111110100;
        weights1[17018] <= 16'b0000000000010101;
        weights1[17019] <= 16'b0000000000001010;
        weights1[17020] <= 16'b0000000000010111;
        weights1[17021] <= 16'b0000000000010100;
        weights1[17022] <= 16'b0000000000010011;
        weights1[17023] <= 16'b0000000000000000;
        weights1[17024] <= 16'b1111111111110010;
        weights1[17025] <= 16'b1111111111100100;
        weights1[17026] <= 16'b1111111111100000;
        weights1[17027] <= 16'b1111111111010100;
        weights1[17028] <= 16'b1111111111011010;
        weights1[17029] <= 16'b1111111111101101;
        weights1[17030] <= 16'b0000000000000010;
        weights1[17031] <= 16'b1111111111111110;
        weights1[17032] <= 16'b0000000000011100;
        weights1[17033] <= 16'b0000000000001011;
        weights1[17034] <= 16'b0000000000010010;
        weights1[17035] <= 16'b0000000000010110;
        weights1[17036] <= 16'b0000000000010110;
        weights1[17037] <= 16'b0000000000000000;
        weights1[17038] <= 16'b1111111111110101;
        weights1[17039] <= 16'b1111111111111101;
        weights1[17040] <= 16'b1111111111101111;
        weights1[17041] <= 16'b1111111111101001;
        weights1[17042] <= 16'b1111111111111010;
        weights1[17043] <= 16'b1111111111110111;
        weights1[17044] <= 16'b1111111111111011;
        weights1[17045] <= 16'b0000000000001101;
        weights1[17046] <= 16'b1111111111111111;
        weights1[17047] <= 16'b0000000000000101;
        weights1[17048] <= 16'b0000000000010001;
        weights1[17049] <= 16'b0000000000001001;
        weights1[17050] <= 16'b0000000000000101;
        weights1[17051] <= 16'b0000000000000100;
        weights1[17052] <= 16'b1111111111110110;
        weights1[17053] <= 16'b1111111111101010;
        weights1[17054] <= 16'b1111111111110010;
        weights1[17055] <= 16'b1111111111110101;
        weights1[17056] <= 16'b1111111111111111;
        weights1[17057] <= 16'b0000000000011001;
        weights1[17058] <= 16'b1111111111101111;
        weights1[17059] <= 16'b0000000000001011;
        weights1[17060] <= 16'b0000000000010001;
        weights1[17061] <= 16'b0000000000010101;
        weights1[17062] <= 16'b0000000000010011;
        weights1[17063] <= 16'b0000000000010001;
        weights1[17064] <= 16'b1111111111111111;
        weights1[17065] <= 16'b0000000000000000;
        weights1[17066] <= 16'b1111111111011101;
        weights1[17067] <= 16'b1111111111101110;
        weights1[17068] <= 16'b1111111111100110;
        weights1[17069] <= 16'b1111111111110010;
        weights1[17070] <= 16'b1111111111110010;
        weights1[17071] <= 16'b1111111111111110;
        weights1[17072] <= 16'b1111111111101111;
        weights1[17073] <= 16'b0000000000010110;
        weights1[17074] <= 16'b0000000000001100;
        weights1[17075] <= 16'b0000000000001110;
        weights1[17076] <= 16'b0000000000000100;
        weights1[17077] <= 16'b0000000000001100;
        weights1[17078] <= 16'b0000000000000001;
        weights1[17079] <= 16'b0000000000000101;
        weights1[17080] <= 16'b1111111111111011;
        weights1[17081] <= 16'b1111111111111110;
        weights1[17082] <= 16'b0000000000000111;
        weights1[17083] <= 16'b0000000000011011;
        weights1[17084] <= 16'b0000000000000010;
        weights1[17085] <= 16'b0000000000010101;
        weights1[17086] <= 16'b1111111111111010;
        weights1[17087] <= 16'b0000000000001111;
        weights1[17088] <= 16'b0000000000001000;
        weights1[17089] <= 16'b0000000000000111;
        weights1[17090] <= 16'b1111111111110110;
        weights1[17091] <= 16'b1111111111111110;
        weights1[17092] <= 16'b1111111111111110;
        weights1[17093] <= 16'b1111111111110010;
        weights1[17094] <= 16'b0000000000010010;
        weights1[17095] <= 16'b1111111111100000;
        weights1[17096] <= 16'b1111111111110101;
        weights1[17097] <= 16'b0000000000001000;
        weights1[17098] <= 16'b1111111111110001;
        weights1[17099] <= 16'b0000000000000000;
        weights1[17100] <= 16'b1111111111110011;
        weights1[17101] <= 16'b0000000000000000;
        weights1[17102] <= 16'b0000000000000010;
        weights1[17103] <= 16'b0000000000000100;
        weights1[17104] <= 16'b1111111111111011;
        weights1[17105] <= 16'b1111111111110111;
        weights1[17106] <= 16'b0000000000000100;
        weights1[17107] <= 16'b0000000000000011;
        weights1[17108] <= 16'b0000000000000101;
        weights1[17109] <= 16'b0000000000000110;
        weights1[17110] <= 16'b0000000000100101;
        weights1[17111] <= 16'b0000000000000101;
        weights1[17112] <= 16'b1111111111111000;
        weights1[17113] <= 16'b0000000000001101;
        weights1[17114] <= 16'b0000000000010000;
        weights1[17115] <= 16'b0000000000011000;
        weights1[17116] <= 16'b0000000000001011;
        weights1[17117] <= 16'b1111111111110000;
        weights1[17118] <= 16'b0000000000011011;
        weights1[17119] <= 16'b1111111111101010;
        weights1[17120] <= 16'b1111111111110110;
        weights1[17121] <= 16'b0000000000001100;
        weights1[17122] <= 16'b1111111111011101;
        weights1[17123] <= 16'b1111111111110000;
        weights1[17124] <= 16'b1111111111101011;
        weights1[17125] <= 16'b1111111111011111;
        weights1[17126] <= 16'b1111111111110101;
        weights1[17127] <= 16'b1111111111110001;
        weights1[17128] <= 16'b1111111111111100;
        weights1[17129] <= 16'b1111111111111111;
        weights1[17130] <= 16'b1111111111111111;
        weights1[17131] <= 16'b1111111111111100;
        weights1[17132] <= 16'b0000000000000001;
        weights1[17133] <= 16'b1111111111111001;
        weights1[17134] <= 16'b1111111111111011;
        weights1[17135] <= 16'b0000000000000000;
        weights1[17136] <= 16'b0000000000000111;
        weights1[17137] <= 16'b0000000000001000;
        weights1[17138] <= 16'b0000000000011000;
        weights1[17139] <= 16'b0000000000001110;
        weights1[17140] <= 16'b0000000000011001;
        weights1[17141] <= 16'b0000000000011110;
        weights1[17142] <= 16'b1111111111111111;
        weights1[17143] <= 16'b1111111111111111;
        weights1[17144] <= 16'b1111111111111010;
        weights1[17145] <= 16'b0000000000001101;
        weights1[17146] <= 16'b1111111111101011;
        weights1[17147] <= 16'b1111111111011111;
        weights1[17148] <= 16'b0000000000010001;
        weights1[17149] <= 16'b0000000000001010;
        weights1[17150] <= 16'b1111111111110111;
        weights1[17151] <= 16'b0000000000001101;
        weights1[17152] <= 16'b1111111111101110;
        weights1[17153] <= 16'b1111111111101111;
        weights1[17154] <= 16'b1111111111010111;
        weights1[17155] <= 16'b1111111111100100;
        weights1[17156] <= 16'b1111111111110001;
        weights1[17157] <= 16'b1111111111110111;
        weights1[17158] <= 16'b1111111111111001;
        weights1[17159] <= 16'b1111111111101111;
        weights1[17160] <= 16'b1111111111111011;
        weights1[17161] <= 16'b1111111111111010;
        weights1[17162] <= 16'b1111111111111000;
        weights1[17163] <= 16'b1111111111111111;
        weights1[17164] <= 16'b0000000000000111;
        weights1[17165] <= 16'b0000000000010001;
        weights1[17166] <= 16'b0000000000001110;
        weights1[17167] <= 16'b0000000000010001;
        weights1[17168] <= 16'b0000000000100100;
        weights1[17169] <= 16'b0000000000010010;
        weights1[17170] <= 16'b0000000000000010;
        weights1[17171] <= 16'b0000000000001010;
        weights1[17172] <= 16'b0000000000000111;
        weights1[17173] <= 16'b0000000000001101;
        weights1[17174] <= 16'b1111111111101111;
        weights1[17175] <= 16'b0000000000010010;
        weights1[17176] <= 16'b1111111111111110;
        weights1[17177] <= 16'b0000000000001100;
        weights1[17178] <= 16'b1111111111101000;
        weights1[17179] <= 16'b0000000000001110;
        weights1[17180] <= 16'b1111111111100101;
        weights1[17181] <= 16'b1111111111110111;
        weights1[17182] <= 16'b1111111111110011;
        weights1[17183] <= 16'b1111111111010110;
        weights1[17184] <= 16'b1111111111100000;
        weights1[17185] <= 16'b1111111111110010;
        weights1[17186] <= 16'b1111111111101101;
        weights1[17187] <= 16'b1111111111101110;
        weights1[17188] <= 16'b1111111111101011;
        weights1[17189] <= 16'b1111111111110101;
        weights1[17190] <= 16'b1111111111111000;
        weights1[17191] <= 16'b1111111111111111;
        weights1[17192] <= 16'b0000000000000101;
        weights1[17193] <= 16'b0000000000001110;
        weights1[17194] <= 16'b0000000000000110;
        weights1[17195] <= 16'b0000000000001001;
        weights1[17196] <= 16'b0000000000010101;
        weights1[17197] <= 16'b0000000000000011;
        weights1[17198] <= 16'b1111111111110101;
        weights1[17199] <= 16'b0000000000000111;
        weights1[17200] <= 16'b1111111111110011;
        weights1[17201] <= 16'b1111111111111001;
        weights1[17202] <= 16'b1111111111111100;
        weights1[17203] <= 16'b1111111111111001;
        weights1[17204] <= 16'b1111111111111100;
        weights1[17205] <= 16'b0000000000001111;
        weights1[17206] <= 16'b1111111111111001;
        weights1[17207] <= 16'b1111111111110111;
        weights1[17208] <= 16'b0000000000001110;
        weights1[17209] <= 16'b1111111111111111;
        weights1[17210] <= 16'b1111111111111000;
        weights1[17211] <= 16'b1111111111111100;
        weights1[17212] <= 16'b1111111111101111;
        weights1[17213] <= 16'b1111111111101110;
        weights1[17214] <= 16'b1111111111110100;
        weights1[17215] <= 16'b1111111111101101;
        weights1[17216] <= 16'b1111111111110100;
        weights1[17217] <= 16'b1111111111111110;
        weights1[17218] <= 16'b1111111111111111;
        weights1[17219] <= 16'b0000000000000000;
        weights1[17220] <= 16'b0000000000000011;
        weights1[17221] <= 16'b0000000000001001;
        weights1[17222] <= 16'b0000000000001110;
        weights1[17223] <= 16'b0000000000010001;
        weights1[17224] <= 16'b0000000000010001;
        weights1[17225] <= 16'b0000000000001100;
        weights1[17226] <= 16'b0000000000000000;
        weights1[17227] <= 16'b1111111111100100;
        weights1[17228] <= 16'b1111111111100011;
        weights1[17229] <= 16'b1111111111110100;
        weights1[17230] <= 16'b1111111111100101;
        weights1[17231] <= 16'b1111111111011100;
        weights1[17232] <= 16'b1111111111101011;
        weights1[17233] <= 16'b1111111111111101;
        weights1[17234] <= 16'b1111111111110100;
        weights1[17235] <= 16'b1111111111101010;
        weights1[17236] <= 16'b1111111111110010;
        weights1[17237] <= 16'b1111111111101111;
        weights1[17238] <= 16'b0000000000000011;
        weights1[17239] <= 16'b1111111111111101;
        weights1[17240] <= 16'b0000000000000011;
        weights1[17241] <= 16'b1111111111111101;
        weights1[17242] <= 16'b1111111111110100;
        weights1[17243] <= 16'b1111111111110111;
        weights1[17244] <= 16'b1111111111111011;
        weights1[17245] <= 16'b0000000000000010;
        weights1[17246] <= 16'b0000000000000000;
        weights1[17247] <= 16'b0000000000000001;
        weights1[17248] <= 16'b0000000000000000;
        weights1[17249] <= 16'b0000000000000001;
        weights1[17250] <= 16'b0000000000000000;
        weights1[17251] <= 16'b0000000000000001;
        weights1[17252] <= 16'b0000000000001101;
        weights1[17253] <= 16'b0000000000011101;
        weights1[17254] <= 16'b0000000000100011;
        weights1[17255] <= 16'b0000000000101110;
        weights1[17256] <= 16'b0000000000101011;
        weights1[17257] <= 16'b0000000000011101;
        weights1[17258] <= 16'b0000000000011110;
        weights1[17259] <= 16'b0000000000010111;
        weights1[17260] <= 16'b0000000000011100;
        weights1[17261] <= 16'b0000000000100111;
        weights1[17262] <= 16'b0000000000100001;
        weights1[17263] <= 16'b0000000000100000;
        weights1[17264] <= 16'b0000000000000111;
        weights1[17265] <= 16'b0000000000001110;
        weights1[17266] <= 16'b0000000000010010;
        weights1[17267] <= 16'b1111111111111111;
        weights1[17268] <= 16'b0000000000000101;
        weights1[17269] <= 16'b0000000000000110;
        weights1[17270] <= 16'b0000000000001001;
        weights1[17271] <= 16'b0000000000001000;
        weights1[17272] <= 16'b0000000000000100;
        weights1[17273] <= 16'b1111111111111011;
        weights1[17274] <= 16'b1111111111111011;
        weights1[17275] <= 16'b1111111111111011;
        weights1[17276] <= 16'b1111111111111111;
        weights1[17277] <= 16'b0000000000000001;
        weights1[17278] <= 16'b0000000000000011;
        weights1[17279] <= 16'b0000000000001110;
        weights1[17280] <= 16'b0000000000011111;
        weights1[17281] <= 16'b0000000000010100;
        weights1[17282] <= 16'b0000000000100011;
        weights1[17283] <= 16'b0000000000011111;
        weights1[17284] <= 16'b0000000000011101;
        weights1[17285] <= 16'b0000000000001001;
        weights1[17286] <= 16'b0000000000000000;
        weights1[17287] <= 16'b0000000000001000;
        weights1[17288] <= 16'b1111111111101100;
        weights1[17289] <= 16'b1111111111111000;
        weights1[17290] <= 16'b1111111111111101;
        weights1[17291] <= 16'b1111111111111100;
        weights1[17292] <= 16'b1111111111111010;
        weights1[17293] <= 16'b1111111111111001;
        weights1[17294] <= 16'b1111111111111111;
        weights1[17295] <= 16'b0000000000000100;
        weights1[17296] <= 16'b0000000000001001;
        weights1[17297] <= 16'b0000000000001000;
        weights1[17298] <= 16'b1111111111110010;
        weights1[17299] <= 16'b0000000000000000;
        weights1[17300] <= 16'b0000000000000100;
        weights1[17301] <= 16'b0000000000000101;
        weights1[17302] <= 16'b1111111111111110;
        weights1[17303] <= 16'b0000000000000011;
        weights1[17304] <= 16'b0000000000000001;
        weights1[17305] <= 16'b0000000000000111;
        weights1[17306] <= 16'b0000000000001011;
        weights1[17307] <= 16'b0000000000011011;
        weights1[17308] <= 16'b0000000000011101;
        weights1[17309] <= 16'b0000000000011001;
        weights1[17310] <= 16'b0000000000100010;
        weights1[17311] <= 16'b0000000000100111;
        weights1[17312] <= 16'b0000000000100101;
        weights1[17313] <= 16'b0000000000100110;
        weights1[17314] <= 16'b0000000000010011;
        weights1[17315] <= 16'b0000000000001001;
        weights1[17316] <= 16'b0000000000010001;
        weights1[17317] <= 16'b1111111111111110;
        weights1[17318] <= 16'b1111111111101110;
        weights1[17319] <= 16'b1111111111110110;
        weights1[17320] <= 16'b0000000000000111;
        weights1[17321] <= 16'b1111111111111110;
        weights1[17322] <= 16'b1111111111110011;
        weights1[17323] <= 16'b0000000000000110;
        weights1[17324] <= 16'b1111111111111110;
        weights1[17325] <= 16'b0000000000000011;
        weights1[17326] <= 16'b0000000000000100;
        weights1[17327] <= 16'b0000000000000111;
        weights1[17328] <= 16'b0000000000010010;
        weights1[17329] <= 16'b1111111111111100;
        weights1[17330] <= 16'b1111111111101110;
        weights1[17331] <= 16'b1111111111111000;
        weights1[17332] <= 16'b0000000000000010;
        weights1[17333] <= 16'b0000000000001100;
        weights1[17334] <= 16'b0000000000001000;
        weights1[17335] <= 16'b0000000000011100;
        weights1[17336] <= 16'b0000000000011100;
        weights1[17337] <= 16'b0000000000100011;
        weights1[17338] <= 16'b0000000000100101;
        weights1[17339] <= 16'b0000000000111101;
        weights1[17340] <= 16'b0000000001000101;
        weights1[17341] <= 16'b0000000000101011;
        weights1[17342] <= 16'b0000000000110000;
        weights1[17343] <= 16'b0000000000011010;
        weights1[17344] <= 16'b0000000000000110;
        weights1[17345] <= 16'b0000000000101100;
        weights1[17346] <= 16'b0000000000011001;
        weights1[17347] <= 16'b1111111111111111;
        weights1[17348] <= 16'b0000000000010011;
        weights1[17349] <= 16'b0000000000010000;
        weights1[17350] <= 16'b0000000000000100;
        weights1[17351] <= 16'b1111111111111100;
        weights1[17352] <= 16'b1111111111110111;
        weights1[17353] <= 16'b0000000000000000;
        weights1[17354] <= 16'b1111111111110001;
        weights1[17355] <= 16'b0000000000001001;
        weights1[17356] <= 16'b0000000000010000;
        weights1[17357] <= 16'b1111111111110101;
        weights1[17358] <= 16'b0000000000000000;
        weights1[17359] <= 16'b1111111111111000;
        weights1[17360] <= 16'b0000000000000110;
        weights1[17361] <= 16'b0000000000001100;
        weights1[17362] <= 16'b0000000000000110;
        weights1[17363] <= 16'b0000000000011000;
        weights1[17364] <= 16'b0000000000100110;
        weights1[17365] <= 16'b0000000000110001;
        weights1[17366] <= 16'b0000000001000101;
        weights1[17367] <= 16'b0000000000111100;
        weights1[17368] <= 16'b0000000000101101;
        weights1[17369] <= 16'b0000000000110010;
        weights1[17370] <= 16'b0000000001000001;
        weights1[17371] <= 16'b0000000000011110;
        weights1[17372] <= 16'b0000000000011010;
        weights1[17373] <= 16'b0000000000000110;
        weights1[17374] <= 16'b0000000000001010;
        weights1[17375] <= 16'b0000000000010001;
        weights1[17376] <= 16'b0000000000010001;
        weights1[17377] <= 16'b0000000000000101;
        weights1[17378] <= 16'b0000000000000101;
        weights1[17379] <= 16'b0000000000001111;
        weights1[17380] <= 16'b0000000000010011;
        weights1[17381] <= 16'b0000000000000001;
        weights1[17382] <= 16'b0000000000000000;
        weights1[17383] <= 16'b1111111111110101;
        weights1[17384] <= 16'b0000000000000100;
        weights1[17385] <= 16'b0000000000000001;
        weights1[17386] <= 16'b0000000000000000;
        weights1[17387] <= 16'b0000000000000001;
        weights1[17388] <= 16'b0000000000000010;
        weights1[17389] <= 16'b0000000000000001;
        weights1[17390] <= 16'b0000000000000010;
        weights1[17391] <= 16'b0000000000011110;
        weights1[17392] <= 16'b0000000000110010;
        weights1[17393] <= 16'b0000000000100111;
        weights1[17394] <= 16'b0000000000111101;
        weights1[17395] <= 16'b0000000001000111;
        weights1[17396] <= 16'b0000000000110100;
        weights1[17397] <= 16'b0000000000100110;
        weights1[17398] <= 16'b0000000000101110;
        weights1[17399] <= 16'b0000000001001101;
        weights1[17400] <= 16'b0000000000110011;
        weights1[17401] <= 16'b0000000000011001;
        weights1[17402] <= 16'b0000000000010101;
        weights1[17403] <= 16'b0000000000010001;
        weights1[17404] <= 16'b0000000000000111;
        weights1[17405] <= 16'b0000000000000101;
        weights1[17406] <= 16'b0000000000010100;
        weights1[17407] <= 16'b0000000000001010;
        weights1[17408] <= 16'b0000000000001000;
        weights1[17409] <= 16'b1111111111111111;
        weights1[17410] <= 16'b0000000000001010;
        weights1[17411] <= 16'b0000000000000101;
        weights1[17412] <= 16'b0000000000001010;
        weights1[17413] <= 16'b0000000000000111;
        weights1[17414] <= 16'b1111111111111001;
        weights1[17415] <= 16'b1111111111111110;
        weights1[17416] <= 16'b1111111111111100;
        weights1[17417] <= 16'b1111111111111101;
        weights1[17418] <= 16'b1111111111110111;
        weights1[17419] <= 16'b0000000000010000;
        weights1[17420] <= 16'b0000000000101100;
        weights1[17421] <= 16'b0000000000101000;
        weights1[17422] <= 16'b0000000000011100;
        weights1[17423] <= 16'b0000000001010101;
        weights1[17424] <= 16'b0000000001010011;
        weights1[17425] <= 16'b0000000001011101;
        weights1[17426] <= 16'b0000000000111011;
        weights1[17427] <= 16'b0000000001010001;
        weights1[17428] <= 16'b0000000001001001;
        weights1[17429] <= 16'b0000000000110110;
        weights1[17430] <= 16'b0000000000100101;
        weights1[17431] <= 16'b0000000000100011;
        weights1[17432] <= 16'b0000000000011101;
        weights1[17433] <= 16'b0000000000000100;
        weights1[17434] <= 16'b0000000000000101;
        weights1[17435] <= 16'b0000000000001100;
        weights1[17436] <= 16'b0000000000000111;
        weights1[17437] <= 16'b0000000000001001;
        weights1[17438] <= 16'b0000000000000110;
        weights1[17439] <= 16'b0000000000001100;
        weights1[17440] <= 16'b0000000000000011;
        weights1[17441] <= 16'b0000000000000101;
        weights1[17442] <= 16'b1111111111111101;
        weights1[17443] <= 16'b0000000000000010;
        weights1[17444] <= 16'b1111111111100111;
        weights1[17445] <= 16'b1111111111100001;
        weights1[17446] <= 16'b1111111111011100;
        weights1[17447] <= 16'b1111111111101000;
        weights1[17448] <= 16'b1111111111111111;
        weights1[17449] <= 16'b0000000000010001;
        weights1[17450] <= 16'b0000000000011110;
        weights1[17451] <= 16'b0000000000011011;
        weights1[17452] <= 16'b0000000000100101;
        weights1[17453] <= 16'b0000000000000110;
        weights1[17454] <= 16'b0000000000010101;
        weights1[17455] <= 16'b0000000000000011;
        weights1[17456] <= 16'b0000000000001011;
        weights1[17457] <= 16'b0000000000010111;
        weights1[17458] <= 16'b0000000000100010;
        weights1[17459] <= 16'b0000000000001010;
        weights1[17460] <= 16'b0000000000100011;
        weights1[17461] <= 16'b1111111111111111;
        weights1[17462] <= 16'b0000000000001111;
        weights1[17463] <= 16'b1111111111111100;
        weights1[17464] <= 16'b0000000000000100;
        weights1[17465] <= 16'b0000000000001001;
        weights1[17466] <= 16'b0000000000001101;
        weights1[17467] <= 16'b1111111111110101;
        weights1[17468] <= 16'b0000000000001110;
        weights1[17469] <= 16'b0000000000000111;
        weights1[17470] <= 16'b1111111111111111;
        weights1[17471] <= 16'b1111111111110110;
        weights1[17472] <= 16'b1111111111011111;
        weights1[17473] <= 16'b1111111111000111;
        weights1[17474] <= 16'b1111111110011110;
        weights1[17475] <= 16'b1111111110011000;
        weights1[17476] <= 16'b1111111110001011;
        weights1[17477] <= 16'b1111111110010111;
        weights1[17478] <= 16'b1111111110111111;
        weights1[17479] <= 16'b1111111110011110;
        weights1[17480] <= 16'b1111111110101001;
        weights1[17481] <= 16'b1111111110010001;
        weights1[17482] <= 16'b1111111110110000;
        weights1[17483] <= 16'b1111111110111110;
        weights1[17484] <= 16'b1111111110111111;
        weights1[17485] <= 16'b1111111111001000;
        weights1[17486] <= 16'b1111111111000111;
        weights1[17487] <= 16'b1111111111010110;
        weights1[17488] <= 16'b1111111111101001;
        weights1[17489] <= 16'b1111111111111010;
        weights1[17490] <= 16'b0000000000001001;
        weights1[17491] <= 16'b1111111111110011;
        weights1[17492] <= 16'b1111111111111111;
        weights1[17493] <= 16'b1111111111111110;
        weights1[17494] <= 16'b0000000000001010;
        weights1[17495] <= 16'b0000000000000011;
        weights1[17496] <= 16'b1111111111111011;
        weights1[17497] <= 16'b0000000000000001;
        weights1[17498] <= 16'b1111111111111011;
        weights1[17499] <= 16'b0000000000000100;
        weights1[17500] <= 16'b1111111111001100;
        weights1[17501] <= 16'b1111111110011001;
        weights1[17502] <= 16'b1111111101111011;
        weights1[17503] <= 16'b1111111101100001;
        weights1[17504] <= 16'b1111111101010101;
        weights1[17505] <= 16'b1111111100110101;
        weights1[17506] <= 16'b1111111100001100;
        weights1[17507] <= 16'b1111111011101100;
        weights1[17508] <= 16'b1111111011101111;
        weights1[17509] <= 16'b1111111100000000;
        weights1[17510] <= 16'b1111111100011101;
        weights1[17511] <= 16'b1111111100111100;
        weights1[17512] <= 16'b1111111101110100;
        weights1[17513] <= 16'b1111111110011001;
        weights1[17514] <= 16'b1111111111000011;
        weights1[17515] <= 16'b1111111111001111;
        weights1[17516] <= 16'b1111111111011000;
        weights1[17517] <= 16'b1111111111100111;
        weights1[17518] <= 16'b1111111111111000;
        weights1[17519] <= 16'b1111111111110001;
        weights1[17520] <= 16'b0000000000001100;
        weights1[17521] <= 16'b1111111111100100;
        weights1[17522] <= 16'b0000000000000101;
        weights1[17523] <= 16'b0000000000000110;
        weights1[17524] <= 16'b0000000000000011;
        weights1[17525] <= 16'b0000000000000001;
        weights1[17526] <= 16'b1111111111111100;
        weights1[17527] <= 16'b1111111111101001;
        weights1[17528] <= 16'b1111111110111011;
        weights1[17529] <= 16'b1111111101111011;
        weights1[17530] <= 16'b1111111101100000;
        weights1[17531] <= 16'b1111111101001011;
        weights1[17532] <= 16'b1111111100101110;
        weights1[17533] <= 16'b1111111011111010;
        weights1[17534] <= 16'b1111111011110111;
        weights1[17535] <= 16'b1111111011111010;
        weights1[17536] <= 16'b1111111100011011;
        weights1[17537] <= 16'b1111111110000001;
        weights1[17538] <= 16'b1111111110111000;
        weights1[17539] <= 16'b1111111111010110;
        weights1[17540] <= 16'b1111111111101000;
        weights1[17541] <= 16'b1111111111101110;
        weights1[17542] <= 16'b1111111111101011;
        weights1[17543] <= 16'b1111111111101101;
        weights1[17544] <= 16'b1111111111110111;
        weights1[17545] <= 16'b1111111111101001;
        weights1[17546] <= 16'b1111111111110101;
        weights1[17547] <= 16'b1111111111111001;
        weights1[17548] <= 16'b1111111111111001;
        weights1[17549] <= 16'b0000000000001100;
        weights1[17550] <= 16'b1111111111111001;
        weights1[17551] <= 16'b1111111111111100;
        weights1[17552] <= 16'b0000000000010100;
        weights1[17553] <= 16'b1111111111110111;
        weights1[17554] <= 16'b0000000000000110;
        weights1[17555] <= 16'b1111111111110000;
        weights1[17556] <= 16'b1111111111000000;
        weights1[17557] <= 16'b1111111110010100;
        weights1[17558] <= 16'b1111111101110011;
        weights1[17559] <= 16'b1111111101110000;
        weights1[17560] <= 16'b1111111101110010;
        weights1[17561] <= 16'b1111111110000111;
        weights1[17562] <= 16'b1111111110100110;
        weights1[17563] <= 16'b1111111111010111;
        weights1[17564] <= 16'b1111111111111101;
        weights1[17565] <= 16'b1111111111111110;
        weights1[17566] <= 16'b1111111111110111;
        weights1[17567] <= 16'b0000000000000000;
        weights1[17568] <= 16'b1111111111111000;
        weights1[17569] <= 16'b1111111111111001;
        weights1[17570] <= 16'b1111111111111011;
        weights1[17571] <= 16'b0000000000000010;
        weights1[17572] <= 16'b0000000000000010;
        weights1[17573] <= 16'b0000000000010101;
        weights1[17574] <= 16'b1111111111111011;
        weights1[17575] <= 16'b0000000000000010;
        weights1[17576] <= 16'b0000000000001100;
        weights1[17577] <= 16'b0000000000000000;
        weights1[17578] <= 16'b1111111111110010;
        weights1[17579] <= 16'b0000000000001000;
        weights1[17580] <= 16'b1111111111111101;
        weights1[17581] <= 16'b1111111111111100;
        weights1[17582] <= 16'b1111111111100111;
        weights1[17583] <= 16'b1111111111110001;
        weights1[17584] <= 16'b1111111111010100;
        weights1[17585] <= 16'b1111111110110010;
        weights1[17586] <= 16'b1111111111001000;
        weights1[17587] <= 16'b1111111111001010;
        weights1[17588] <= 16'b1111111111101011;
        weights1[17589] <= 16'b1111111111110110;
        weights1[17590] <= 16'b0000000000011101;
        weights1[17591] <= 16'b0000000000100111;
        weights1[17592] <= 16'b0000000000111001;
        weights1[17593] <= 16'b0000000000100001;
        weights1[17594] <= 16'b0000000000011110;
        weights1[17595] <= 16'b0000000000010111;
        weights1[17596] <= 16'b0000000000010001;
        weights1[17597] <= 16'b0000000000000110;
        weights1[17598] <= 16'b0000000000001010;
        weights1[17599] <= 16'b0000000000000100;
        weights1[17600] <= 16'b0000000000001000;
        weights1[17601] <= 16'b1111111111110010;
        weights1[17602] <= 16'b0000000000001100;
        weights1[17603] <= 16'b1111111111110100;
        weights1[17604] <= 16'b1111111111111111;
        weights1[17605] <= 16'b1111111111110111;
        weights1[17606] <= 16'b0000000000010011;
        weights1[17607] <= 16'b0000000000000001;
        weights1[17608] <= 16'b1111111111101110;
        weights1[17609] <= 16'b0000000000010010;
        weights1[17610] <= 16'b0000000000000010;
        weights1[17611] <= 16'b0000000000000011;
        weights1[17612] <= 16'b1111111111101110;
        weights1[17613] <= 16'b1111111111111011;
        weights1[17614] <= 16'b0000000000000101;
        weights1[17615] <= 16'b0000000000010011;
        weights1[17616] <= 16'b0000000000111010;
        weights1[17617] <= 16'b0000000000100101;
        weights1[17618] <= 16'b0000000000100000;
        weights1[17619] <= 16'b0000000000011100;
        weights1[17620] <= 16'b0000000000100000;
        weights1[17621] <= 16'b0000000000001100;
        weights1[17622] <= 16'b0000000000001111;
        weights1[17623] <= 16'b0000000000010001;
        weights1[17624] <= 16'b0000000000011000;
        weights1[17625] <= 16'b0000000000011110;
        weights1[17626] <= 16'b0000000000001000;
        weights1[17627] <= 16'b0000000000010001;
        weights1[17628] <= 16'b0000000000001001;
        weights1[17629] <= 16'b0000000000000010;
        weights1[17630] <= 16'b1111111111111011;
        weights1[17631] <= 16'b0000000000001100;
        weights1[17632] <= 16'b0000000000000001;
        weights1[17633] <= 16'b0000000000000000;
        weights1[17634] <= 16'b0000000000001001;
        weights1[17635] <= 16'b0000000000000000;
        weights1[17636] <= 16'b1111111111111110;
        weights1[17637] <= 16'b1111111111111010;
        weights1[17638] <= 16'b0000000000001001;
        weights1[17639] <= 16'b1111111111111000;
        weights1[17640] <= 16'b1111111111111011;
        weights1[17641] <= 16'b0000000000100101;
        weights1[17642] <= 16'b0000000000011010;
        weights1[17643] <= 16'b0000000000111001;
        weights1[17644] <= 16'b0000000000111001;
        weights1[17645] <= 16'b0000000000110000;
        weights1[17646] <= 16'b0000000000101001;
        weights1[17647] <= 16'b0000000000011100;
        weights1[17648] <= 16'b0000000000011111;
        weights1[17649] <= 16'b0000000000010110;
        weights1[17650] <= 16'b0000000000000000;
        weights1[17651] <= 16'b0000000000010100;
        weights1[17652] <= 16'b1111111111111010;
        weights1[17653] <= 16'b0000000000000001;
        weights1[17654] <= 16'b1111111111111100;
        weights1[17655] <= 16'b0000000000001001;
        weights1[17656] <= 16'b0000000000001011;
        weights1[17657] <= 16'b1111111111111001;
        weights1[17658] <= 16'b0000000000010010;
        weights1[17659] <= 16'b1111111111111101;
        weights1[17660] <= 16'b0000000000001111;
        weights1[17661] <= 16'b1111111111111110;
        weights1[17662] <= 16'b1111111111101110;
        weights1[17663] <= 16'b0000000000000011;
        weights1[17664] <= 16'b1111111111111010;
        weights1[17665] <= 16'b1111111111111100;
        weights1[17666] <= 16'b0000000000000001;
        weights1[17667] <= 16'b0000000000000011;
        weights1[17668] <= 16'b0000000000001101;
        weights1[17669] <= 16'b0000000000100010;
        weights1[17670] <= 16'b0000000000100001;
        weights1[17671] <= 16'b0000000000001100;
        weights1[17672] <= 16'b0000000000000000;
        weights1[17673] <= 16'b0000000000010011;
        weights1[17674] <= 16'b0000000000000111;
        weights1[17675] <= 16'b1111111111110101;
        weights1[17676] <= 16'b1111111111111011;
        weights1[17677] <= 16'b0000000000000111;
        weights1[17678] <= 16'b0000000000001010;
        weights1[17679] <= 16'b0000000000000011;
        weights1[17680] <= 16'b0000000000010010;
        weights1[17681] <= 16'b0000000000000100;
        weights1[17682] <= 16'b0000000000001000;
        weights1[17683] <= 16'b0000000000000010;
        weights1[17684] <= 16'b0000000000001111;
        weights1[17685] <= 16'b0000000000000011;
        weights1[17686] <= 16'b1111111111110111;
        weights1[17687] <= 16'b1111111111110101;
        weights1[17688] <= 16'b1111111111111110;
        weights1[17689] <= 16'b0000000000000110;
        weights1[17690] <= 16'b0000000000000100;
        weights1[17691] <= 16'b0000000000000001;
        weights1[17692] <= 16'b0000000000000011;
        weights1[17693] <= 16'b1111111111111100;
        weights1[17694] <= 16'b1111111111111011;
        weights1[17695] <= 16'b0000000000000101;
        weights1[17696] <= 16'b0000000000011000;
        weights1[17697] <= 16'b0000000000010010;
        weights1[17698] <= 16'b1111111111111111;
        weights1[17699] <= 16'b0000000000000010;
        weights1[17700] <= 16'b1111111111110100;
        weights1[17701] <= 16'b1111111111111000;
        weights1[17702] <= 16'b0000000000001010;
        weights1[17703] <= 16'b1111111111111000;
        weights1[17704] <= 16'b0000000000000011;
        weights1[17705] <= 16'b0000000000001000;
        weights1[17706] <= 16'b0000000000000111;
        weights1[17707] <= 16'b1111111111110111;
        weights1[17708] <= 16'b1111111111110011;
        weights1[17709] <= 16'b0000000000000111;
        weights1[17710] <= 16'b1111111111111010;
        weights1[17711] <= 16'b1111111111110110;
        weights1[17712] <= 16'b1111111111110011;
        weights1[17713] <= 16'b0000000000000010;
        weights1[17714] <= 16'b0000000000000000;
        weights1[17715] <= 16'b1111111111111000;
        weights1[17716] <= 16'b1111111111111101;
        weights1[17717] <= 16'b1111111111110110;
        weights1[17718] <= 16'b0000000000001011;
        weights1[17719] <= 16'b1111111111110001;
        weights1[17720] <= 16'b0000000000000101;
        weights1[17721] <= 16'b1111111111111110;
        weights1[17722] <= 16'b0000000000000101;
        weights1[17723] <= 16'b0000000000010101;
        weights1[17724] <= 16'b0000000000001111;
        weights1[17725] <= 16'b0000000000001110;
        weights1[17726] <= 16'b1111111111110001;
        weights1[17727] <= 16'b1111111111110110;
        weights1[17728] <= 16'b0000000000001000;
        weights1[17729] <= 16'b0000000000001110;
        weights1[17730] <= 16'b1111111111111011;
        weights1[17731] <= 16'b0000000000000000;
        weights1[17732] <= 16'b0000000000001010;
        weights1[17733] <= 16'b1111111111101000;
        weights1[17734] <= 16'b0000000000000010;
        weights1[17735] <= 16'b0000000000000001;
        weights1[17736] <= 16'b1111111111111101;
        weights1[17737] <= 16'b1111111111110101;
        weights1[17738] <= 16'b1111111111111010;
        weights1[17739] <= 16'b1111111111111110;
        weights1[17740] <= 16'b1111111111111111;
        weights1[17741] <= 16'b1111111111111011;
        weights1[17742] <= 16'b1111111111110100;
        weights1[17743] <= 16'b0000000000000001;
        weights1[17744] <= 16'b0000000000000010;
        weights1[17745] <= 16'b1111111111111010;
        weights1[17746] <= 16'b0000000000000101;
        weights1[17747] <= 16'b1111111111110111;
        weights1[17748] <= 16'b0000000000000100;
        weights1[17749] <= 16'b0000000000000101;
        weights1[17750] <= 16'b0000000000000111;
        weights1[17751] <= 16'b0000000000000011;
        weights1[17752] <= 16'b0000000000001101;
        weights1[17753] <= 16'b0000000000000011;
        weights1[17754] <= 16'b1111111111101010;
        weights1[17755] <= 16'b1111111111101101;
        weights1[17756] <= 16'b1111111111101110;
        weights1[17757] <= 16'b0000000000000000;
        weights1[17758] <= 16'b1111111111110100;
        weights1[17759] <= 16'b1111111111110111;
        weights1[17760] <= 16'b0000000000010011;
        weights1[17761] <= 16'b0000000000000110;
        weights1[17762] <= 16'b0000000000000010;
        weights1[17763] <= 16'b0000000000000111;
        weights1[17764] <= 16'b1111111111111100;
        weights1[17765] <= 16'b0000000000000000;
        weights1[17766] <= 16'b1111111111111110;
        weights1[17767] <= 16'b1111111111100110;
        weights1[17768] <= 16'b0000000000010010;
        weights1[17769] <= 16'b1111111111110101;
        weights1[17770] <= 16'b1111111111111000;
        weights1[17771] <= 16'b1111111111111011;
        weights1[17772] <= 16'b0000000000000110;
        weights1[17773] <= 16'b0000000000010100;
        weights1[17774] <= 16'b0000000000000110;
        weights1[17775] <= 16'b0000000000010100;
        weights1[17776] <= 16'b1111111111110000;
        weights1[17777] <= 16'b0000000000001010;
        weights1[17778] <= 16'b1111111111111101;
        weights1[17779] <= 16'b0000000000000111;
        weights1[17780] <= 16'b1111111111111001;
        weights1[17781] <= 16'b1111111111111000;
        weights1[17782] <= 16'b1111111111011010;
        weights1[17783] <= 16'b1111111111101101;
        weights1[17784] <= 16'b0000000000001110;
        weights1[17785] <= 16'b0000000000001111;
        weights1[17786] <= 16'b0000000000000010;
        weights1[17787] <= 16'b1111111111110100;
        weights1[17788] <= 16'b1111111111110110;
        weights1[17789] <= 16'b1111111111111011;
        weights1[17790] <= 16'b0000000000000010;
        weights1[17791] <= 16'b0000000000000001;
        weights1[17792] <= 16'b1111111111110100;
        weights1[17793] <= 16'b1111111111111010;
        weights1[17794] <= 16'b0000000000000100;
        weights1[17795] <= 16'b1111111111110100;
        weights1[17796] <= 16'b1111111111111010;
        weights1[17797] <= 16'b0000000000000010;
        weights1[17798] <= 16'b0000000000000110;
        weights1[17799] <= 16'b1111111111111101;
        weights1[17800] <= 16'b1111111111111001;
        weights1[17801] <= 16'b1111111111101101;
        weights1[17802] <= 16'b1111111111100101;
        weights1[17803] <= 16'b1111111111110100;
        weights1[17804] <= 16'b1111111111111101;
        weights1[17805] <= 16'b1111111111111001;
        weights1[17806] <= 16'b1111111111111110;
        weights1[17807] <= 16'b0000000000001000;
        weights1[17808] <= 16'b1111111111110101;
        weights1[17809] <= 16'b1111111111111111;
        weights1[17810] <= 16'b1111111111100110;
        weights1[17811] <= 16'b1111111111111110;
        weights1[17812] <= 16'b0000000000000101;
        weights1[17813] <= 16'b0000000000010100;
        weights1[17814] <= 16'b1111111111111001;
        weights1[17815] <= 16'b0000000000001000;
        weights1[17816] <= 16'b1111111111111111;
        weights1[17817] <= 16'b1111111111110101;
        weights1[17818] <= 16'b1111111111111111;
        weights1[17819] <= 16'b0000000000000000;
        weights1[17820] <= 16'b1111111111111000;
        weights1[17821] <= 16'b0000000000001010;
        weights1[17822] <= 16'b1111111111110111;
        weights1[17823] <= 16'b1111111111111111;
        weights1[17824] <= 16'b1111111111110001;
        weights1[17825] <= 16'b1111111111111110;
        weights1[17826] <= 16'b1111111111111001;
        weights1[17827] <= 16'b1111111111111101;
        weights1[17828] <= 16'b1111111111110111;
        weights1[17829] <= 16'b0000000000000101;
        weights1[17830] <= 16'b0000000000000111;
        weights1[17831] <= 16'b0000000000001000;
        weights1[17832] <= 16'b0000000000001000;
        weights1[17833] <= 16'b0000000000000011;
        weights1[17834] <= 16'b1111111111111100;
        weights1[17835] <= 16'b1111111111111011;
        weights1[17836] <= 16'b1111111111110100;
        weights1[17837] <= 16'b1111111111110100;
        weights1[17838] <= 16'b1111111111100101;
        weights1[17839] <= 16'b1111111111110111;
        weights1[17840] <= 16'b1111111111111010;
        weights1[17841] <= 16'b0000000000000001;
        weights1[17842] <= 16'b0000000000000000;
        weights1[17843] <= 16'b1111111111111000;
        weights1[17844] <= 16'b1111111111111110;
        weights1[17845] <= 16'b1111111111111100;
        weights1[17846] <= 16'b1111111111111001;
        weights1[17847] <= 16'b1111111111100010;
        weights1[17848] <= 16'b1111111111111111;
        weights1[17849] <= 16'b1111111111101011;
        weights1[17850] <= 16'b1111111111111110;
        weights1[17851] <= 16'b1111111111111101;
        weights1[17852] <= 16'b0000000000000111;
        weights1[17853] <= 16'b1111111111111000;
        weights1[17854] <= 16'b0000000000000100;
        weights1[17855] <= 16'b0000000000000100;
        weights1[17856] <= 16'b1111111111110111;
        weights1[17857] <= 16'b0000000000000010;
        weights1[17858] <= 16'b0000000000000100;
        weights1[17859] <= 16'b0000000000000101;
        weights1[17860] <= 16'b1111111111111010;
        weights1[17861] <= 16'b0000000000000000;
        weights1[17862] <= 16'b0000000000000000;
        weights1[17863] <= 16'b0000000000000100;
        weights1[17864] <= 16'b1111111111110110;
        weights1[17865] <= 16'b1111111111110101;
        weights1[17866] <= 16'b1111111111110100;
        weights1[17867] <= 16'b1111111111110001;
        weights1[17868] <= 16'b1111111111111101;
        weights1[17869] <= 16'b0000000000001000;
        weights1[17870] <= 16'b1111111111101100;
        weights1[17871] <= 16'b1111111111111111;
        weights1[17872] <= 16'b1111111111110000;
        weights1[17873] <= 16'b1111111111110100;
        weights1[17874] <= 16'b0000000000010100;
        weights1[17875] <= 16'b0000000000011000;
        weights1[17876] <= 16'b1111111111111000;
        weights1[17877] <= 16'b0000000000000001;
        weights1[17878] <= 16'b1111111111110111;
        weights1[17879] <= 16'b0000000000001011;
        weights1[17880] <= 16'b1111111111110111;
        weights1[17881] <= 16'b1111111111110011;
        weights1[17882] <= 16'b1111111111111101;
        weights1[17883] <= 16'b1111111111110000;
        weights1[17884] <= 16'b1111111111111010;
        weights1[17885] <= 16'b1111111111110110;
        weights1[17886] <= 16'b1111111111101111;
        weights1[17887] <= 16'b0000000000001001;
        weights1[17888] <= 16'b1111111111111010;
        weights1[17889] <= 16'b1111111111111111;
        weights1[17890] <= 16'b1111111111110100;
        weights1[17891] <= 16'b1111111111111111;
        weights1[17892] <= 16'b1111111111111010;
        weights1[17893] <= 16'b1111111111111000;
        weights1[17894] <= 16'b1111111111110101;
        weights1[17895] <= 16'b1111111111100101;
        weights1[17896] <= 16'b1111111111101100;
        weights1[17897] <= 16'b1111111111101110;
        weights1[17898] <= 16'b1111111111110110;
        weights1[17899] <= 16'b1111111111101110;
        weights1[17900] <= 16'b1111111111111000;
        weights1[17901] <= 16'b1111111111111111;
        weights1[17902] <= 16'b1111111111110101;
        weights1[17903] <= 16'b1111111111110110;
        weights1[17904] <= 16'b1111111111111011;
        weights1[17905] <= 16'b1111111111101111;
        weights1[17906] <= 16'b1111111111111111;
        weights1[17907] <= 16'b1111111111111111;
        weights1[17908] <= 16'b1111111111111010;
        weights1[17909] <= 16'b1111111111110000;
        weights1[17910] <= 16'b1111111111111000;
        weights1[17911] <= 16'b0000000000000100;
        weights1[17912] <= 16'b0000000000011110;
        weights1[17913] <= 16'b0000000000000111;
        weights1[17914] <= 16'b0000000000001000;
        weights1[17915] <= 16'b1111111111111011;
        weights1[17916] <= 16'b0000000000000010;
        weights1[17917] <= 16'b1111111111111000;
        weights1[17918] <= 16'b1111111111111010;
        weights1[17919] <= 16'b0000000000000001;
        weights1[17920] <= 16'b1111111111110111;
        weights1[17921] <= 16'b1111111111101110;
        weights1[17922] <= 16'b1111111111111010;
        weights1[17923] <= 16'b1111111111110100;
        weights1[17924] <= 16'b1111111111110010;
        weights1[17925] <= 16'b1111111111110011;
        weights1[17926] <= 16'b1111111111110010;
        weights1[17927] <= 16'b1111111111111001;
        weights1[17928] <= 16'b0000000000000000;
        weights1[17929] <= 16'b0000000000000001;
        weights1[17930] <= 16'b1111111111110111;
        weights1[17931] <= 16'b1111111111111101;
        weights1[17932] <= 16'b1111111111110101;
        weights1[17933] <= 16'b0000000000010010;
        weights1[17934] <= 16'b1111111111111000;
        weights1[17935] <= 16'b1111111111111011;
        weights1[17936] <= 16'b1111111111111001;
        weights1[17937] <= 16'b0000000000000011;
        weights1[17938] <= 16'b0000000000001010;
        weights1[17939] <= 16'b1111111111110110;
        weights1[17940] <= 16'b1111111111110100;
        weights1[17941] <= 16'b0000000000001011;
        weights1[17942] <= 16'b1111111111111011;
        weights1[17943] <= 16'b0000000000000010;
        weights1[17944] <= 16'b1111111111110101;
        weights1[17945] <= 16'b0000000000000000;
        weights1[17946] <= 16'b1111111111111101;
        weights1[17947] <= 16'b0000000000000101;
        weights1[17948] <= 16'b1111111111111000;
        weights1[17949] <= 16'b1111111111111000;
        weights1[17950] <= 16'b1111111111110011;
        weights1[17951] <= 16'b1111111111110110;
        weights1[17952] <= 16'b0000000000000001;
        weights1[17953] <= 16'b1111111111111011;
        weights1[17954] <= 16'b1111111111101000;
        weights1[17955] <= 16'b1111111111100010;
        weights1[17956] <= 16'b1111111111110100;
        weights1[17957] <= 16'b1111111111110000;
        weights1[17958] <= 16'b1111111111111110;
        weights1[17959] <= 16'b1111111111101011;
        weights1[17960] <= 16'b1111111111111001;
        weights1[17961] <= 16'b1111111111111111;
        weights1[17962] <= 16'b1111111111100110;
        weights1[17963] <= 16'b0000000000010001;
        weights1[17964] <= 16'b1111111111110110;
        weights1[17965] <= 16'b0000000000000110;
        weights1[17966] <= 16'b0000000000000101;
        weights1[17967] <= 16'b0000000000000100;
        weights1[17968] <= 16'b0000000000000101;
        weights1[17969] <= 16'b1111111111111111;
        weights1[17970] <= 16'b1111111111111100;
        weights1[17971] <= 16'b1111111111111011;
        weights1[17972] <= 16'b1111111111110110;
        weights1[17973] <= 16'b0000000000000011;
        weights1[17974] <= 16'b0000000000000000;
        weights1[17975] <= 16'b0000000000000001;
        weights1[17976] <= 16'b1111111111111100;
        weights1[17977] <= 16'b1111111111111110;
        weights1[17978] <= 16'b1111111111110111;
        weights1[17979] <= 16'b0000000000000100;
        weights1[17980] <= 16'b1111111111110111;
        weights1[17981] <= 16'b1111111111110011;
        weights1[17982] <= 16'b1111111111101111;
        weights1[17983] <= 16'b1111111111101010;
        weights1[17984] <= 16'b1111111111101011;
        weights1[17985] <= 16'b1111111111100111;
        weights1[17986] <= 16'b1111111111100111;
        weights1[17987] <= 16'b1111111111101100;
        weights1[17988] <= 16'b1111111111110011;
        weights1[17989] <= 16'b1111111111101011;
        weights1[17990] <= 16'b0000000000000110;
        weights1[17991] <= 16'b1111111111111110;
        weights1[17992] <= 16'b1111111111111010;
        weights1[17993] <= 16'b0000000000000000;
        weights1[17994] <= 16'b1111111111101011;
        weights1[17995] <= 16'b1111111111111101;
        weights1[17996] <= 16'b0000000000000110;
        weights1[17997] <= 16'b0000000000001000;
        weights1[17998] <= 16'b1111111111110111;
        weights1[17999] <= 16'b0000000000000000;
        weights1[18000] <= 16'b0000000000001010;
        weights1[18001] <= 16'b0000000000001001;
        weights1[18002] <= 16'b0000000000000000;
        weights1[18003] <= 16'b0000000000000100;
        weights1[18004] <= 16'b1111111111111111;
        weights1[18005] <= 16'b1111111111111100;
        weights1[18006] <= 16'b1111111111111101;
        weights1[18007] <= 16'b1111111111110011;
        weights1[18008] <= 16'b0000000000000011;
        weights1[18009] <= 16'b1111111111111001;
        weights1[18010] <= 16'b1111111111101101;
        weights1[18011] <= 16'b1111111111111001;
        weights1[18012] <= 16'b0000000000000010;
        weights1[18013] <= 16'b0000000000000111;
        weights1[18014] <= 16'b1111111111111011;
        weights1[18015] <= 16'b0000000000010011;
        weights1[18016] <= 16'b0000000000010110;
        weights1[18017] <= 16'b0000000000011011;
        weights1[18018] <= 16'b0000000000001110;
        weights1[18019] <= 16'b0000000000001010;
        weights1[18020] <= 16'b0000000000010101;
        weights1[18021] <= 16'b0000000000010100;
        weights1[18022] <= 16'b0000000000010001;
        weights1[18023] <= 16'b0000000000001011;
        weights1[18024] <= 16'b0000000000011000;
        weights1[18025] <= 16'b0000000000011000;
        weights1[18026] <= 16'b0000000000010010;
        weights1[18027] <= 16'b0000000000010101;
        weights1[18028] <= 16'b0000000000010010;
        weights1[18029] <= 16'b0000000000001000;
        weights1[18030] <= 16'b0000000000000110;
        weights1[18031] <= 16'b0000000000000011;
        weights1[18032] <= 16'b0000000000000000;
        weights1[18033] <= 16'b1111111111111111;
        weights1[18034] <= 16'b1111111111111111;
        weights1[18035] <= 16'b0000000000000000;
        weights1[18036] <= 16'b0000000000000000;
        weights1[18037] <= 16'b0000000000000000;
        weights1[18038] <= 16'b0000000000000001;
        weights1[18039] <= 16'b0000000000000010;
        weights1[18040] <= 16'b1111111111111001;
        weights1[18041] <= 16'b1111111111111110;
        weights1[18042] <= 16'b0000000000000000;
        weights1[18043] <= 16'b1111111111111100;
        weights1[18044] <= 16'b1111111111111011;
        weights1[18045] <= 16'b1111111111111110;
        weights1[18046] <= 16'b0000000000000001;
        weights1[18047] <= 16'b1111111111111101;
        weights1[18048] <= 16'b1111111111111111;
        weights1[18049] <= 16'b0000000000000011;
        weights1[18050] <= 16'b1111111111111110;
        weights1[18051] <= 16'b1111111111111111;
        weights1[18052] <= 16'b1111111111111110;
        weights1[18053] <= 16'b1111111111111100;
        weights1[18054] <= 16'b1111111111111111;
        weights1[18055] <= 16'b1111111111111111;
        weights1[18056] <= 16'b0000000000000000;
        weights1[18057] <= 16'b1111111111111111;
        weights1[18058] <= 16'b0000000000000000;
        weights1[18059] <= 16'b0000000000000000;
        weights1[18060] <= 16'b1111111111111111;
        weights1[18061] <= 16'b1111111111111110;
        weights1[18062] <= 16'b1111111111111110;
        weights1[18063] <= 16'b1111111111111110;
        weights1[18064] <= 16'b1111111111111111;
        weights1[18065] <= 16'b1111111111111011;
        weights1[18066] <= 16'b0000000000000000;
        weights1[18067] <= 16'b0000000000000000;
        weights1[18068] <= 16'b1111111111110111;
        weights1[18069] <= 16'b1111111111111010;
        weights1[18070] <= 16'b1111111111111000;
        weights1[18071] <= 16'b1111111111111101;
        weights1[18072] <= 16'b1111111111111101;
        weights1[18073] <= 16'b1111111111111010;
        weights1[18074] <= 16'b0000000000000001;
        weights1[18075] <= 16'b1111111111111110;
        weights1[18076] <= 16'b0000000000000100;
        weights1[18077] <= 16'b0000000000000011;
        weights1[18078] <= 16'b1111111111110111;
        weights1[18079] <= 16'b1111111111111000;
        weights1[18080] <= 16'b1111111111110111;
        weights1[18081] <= 16'b1111111111111010;
        weights1[18082] <= 16'b1111111111111110;
        weights1[18083] <= 16'b1111111111111111;
        weights1[18084] <= 16'b0000000000000000;
        weights1[18085] <= 16'b1111111111111101;
        weights1[18086] <= 16'b0000000000000000;
        weights1[18087] <= 16'b0000000000000000;
        weights1[18088] <= 16'b1111111111111111;
        weights1[18089] <= 16'b1111111111111111;
        weights1[18090] <= 16'b1111111111111111;
        weights1[18091] <= 16'b1111111111111100;
        weights1[18092] <= 16'b1111111111111101;
        weights1[18093] <= 16'b1111111111111100;
        weights1[18094] <= 16'b1111111111111011;
        weights1[18095] <= 16'b0000000000000000;
        weights1[18096] <= 16'b1111111111110000;
        weights1[18097] <= 16'b1111111111110010;
        weights1[18098] <= 16'b1111111111101111;
        weights1[18099] <= 16'b1111111111110101;
        weights1[18100] <= 16'b1111111111111001;
        weights1[18101] <= 16'b0000000000000011;
        weights1[18102] <= 16'b1111111111111000;
        weights1[18103] <= 16'b0000000000000100;
        weights1[18104] <= 16'b0000000000001000;
        weights1[18105] <= 16'b0000000000000010;
        weights1[18106] <= 16'b0000000000000111;
        weights1[18107] <= 16'b1111111111110011;
        weights1[18108] <= 16'b1111111111101010;
        weights1[18109] <= 16'b1111111111110111;
        weights1[18110] <= 16'b1111111111111110;
        weights1[18111] <= 16'b1111111111111100;
        weights1[18112] <= 16'b0000000000000000;
        weights1[18113] <= 16'b0000000000000100;
        weights1[18114] <= 16'b0000000000000000;
        weights1[18115] <= 16'b0000000000000000;
        weights1[18116] <= 16'b1111111111111111;
        weights1[18117] <= 16'b1111111111111111;
        weights1[18118] <= 16'b1111111111111110;
        weights1[18119] <= 16'b1111111111111100;
        weights1[18120] <= 16'b1111111111111001;
        weights1[18121] <= 16'b1111111111111000;
        weights1[18122] <= 16'b1111111111110011;
        weights1[18123] <= 16'b1111111111101000;
        weights1[18124] <= 16'b1111111111101100;
        weights1[18125] <= 16'b1111111111101010;
        weights1[18126] <= 16'b1111111111111010;
        weights1[18127] <= 16'b1111111111110101;
        weights1[18128] <= 16'b1111111111100010;
        weights1[18129] <= 16'b1111111111011110;
        weights1[18130] <= 16'b1111111111110111;
        weights1[18131] <= 16'b1111111111110100;
        weights1[18132] <= 16'b1111111111100101;
        weights1[18133] <= 16'b1111111111101010;
        weights1[18134] <= 16'b1111111111110001;
        weights1[18135] <= 16'b1111111111111000;
        weights1[18136] <= 16'b1111111111110100;
        weights1[18137] <= 16'b1111111111111011;
        weights1[18138] <= 16'b1111111111111100;
        weights1[18139] <= 16'b1111111111101111;
        weights1[18140] <= 16'b0000000000000111;
        weights1[18141] <= 16'b1111111111111010;
        weights1[18142] <= 16'b1111111111111100;
        weights1[18143] <= 16'b0000000000000010;
        weights1[18144] <= 16'b1111111111111110;
        weights1[18145] <= 16'b1111111111111101;
        weights1[18146] <= 16'b0000000000000000;
        weights1[18147] <= 16'b1111111111111011;
        weights1[18148] <= 16'b1111111111111010;
        weights1[18149] <= 16'b1111111111111011;
        weights1[18150] <= 16'b1111111111111100;
        weights1[18151] <= 16'b0000000000001001;
        weights1[18152] <= 16'b0000000000000000;
        weights1[18153] <= 16'b1111111111101000;
        weights1[18154] <= 16'b1111111111101001;
        weights1[18155] <= 16'b1111111111101011;
        weights1[18156] <= 16'b1111111111101101;
        weights1[18157] <= 16'b1111111111111010;
        weights1[18158] <= 16'b1111111111111011;
        weights1[18159] <= 16'b0000000000001110;
        weights1[18160] <= 16'b0000000000001100;
        weights1[18161] <= 16'b0000000000010101;
        weights1[18162] <= 16'b0000000000000111;
        weights1[18163] <= 16'b0000000000010011;
        weights1[18164] <= 16'b1111111111111000;
        weights1[18165] <= 16'b1111111111110101;
        weights1[18166] <= 16'b1111111111111110;
        weights1[18167] <= 16'b1111111111101010;
        weights1[18168] <= 16'b1111111111111001;
        weights1[18169] <= 16'b1111111111111110;
        weights1[18170] <= 16'b0000000000000010;
        weights1[18171] <= 16'b0000000000000001;
        weights1[18172] <= 16'b1111111111111110;
        weights1[18173] <= 16'b1111111111111001;
        weights1[18174] <= 16'b1111111111111011;
        weights1[18175] <= 16'b1111111111110011;
        weights1[18176] <= 16'b1111111111110010;
        weights1[18177] <= 16'b1111111111110011;
        weights1[18178] <= 16'b1111111111111000;
        weights1[18179] <= 16'b0000000000000010;
        weights1[18180] <= 16'b1111111111111000;
        weights1[18181] <= 16'b1111111111101010;
        weights1[18182] <= 16'b0000000000000110;
        weights1[18183] <= 16'b1111111111110101;
        weights1[18184] <= 16'b1111111111110010;
        weights1[18185] <= 16'b0000000000000000;
        weights1[18186] <= 16'b1111111111101111;
        weights1[18187] <= 16'b0000000000001111;
        weights1[18188] <= 16'b0000000000010000;
        weights1[18189] <= 16'b0000000000000101;
        weights1[18190] <= 16'b1111111111110101;
        weights1[18191] <= 16'b0000000000001010;
        weights1[18192] <= 16'b1111111111111111;
        weights1[18193] <= 16'b1111111111111100;
        weights1[18194] <= 16'b1111111111111011;
        weights1[18195] <= 16'b1111111111110110;
        weights1[18196] <= 16'b1111111111110101;
        weights1[18197] <= 16'b1111111111111011;
        weights1[18198] <= 16'b1111111111111111;
        weights1[18199] <= 16'b1111111111111101;
        weights1[18200] <= 16'b1111111111111100;
        weights1[18201] <= 16'b1111111111110111;
        weights1[18202] <= 16'b1111111111110010;
        weights1[18203] <= 16'b1111111111110110;
        weights1[18204] <= 16'b1111111111101011;
        weights1[18205] <= 16'b1111111111110100;
        weights1[18206] <= 16'b1111111111111011;
        weights1[18207] <= 16'b1111111111111111;
        weights1[18208] <= 16'b0000000000001011;
        weights1[18209] <= 16'b1111111111111100;
        weights1[18210] <= 16'b1111111111101101;
        weights1[18211] <= 16'b1111111111101011;
        weights1[18212] <= 16'b0000000000000011;
        weights1[18213] <= 16'b1111111111111011;
        weights1[18214] <= 16'b0000000000000001;
        weights1[18215] <= 16'b1111111111110001;
        weights1[18216] <= 16'b1111111111110001;
        weights1[18217] <= 16'b1111111111110000;
        weights1[18218] <= 16'b0000000000001010;
        weights1[18219] <= 16'b0000000000010111;
        weights1[18220] <= 16'b0000000000000110;
        weights1[18221] <= 16'b0000000000000110;
        weights1[18222] <= 16'b0000000000000001;
        weights1[18223] <= 16'b0000000000000101;
        weights1[18224] <= 16'b1111111111111010;
        weights1[18225] <= 16'b0000000000001100;
        weights1[18226] <= 16'b1111111111111100;
        weights1[18227] <= 16'b0000000000001011;
        weights1[18228] <= 16'b1111111111111000;
        weights1[18229] <= 16'b1111111111111000;
        weights1[18230] <= 16'b1111111111111010;
        weights1[18231] <= 16'b0000000000000111;
        weights1[18232] <= 16'b1111111111110111;
        weights1[18233] <= 16'b0000000000000111;
        weights1[18234] <= 16'b0000000000000111;
        weights1[18235] <= 16'b0000000000000110;
        weights1[18236] <= 16'b0000000000000110;
        weights1[18237] <= 16'b1111111111010100;
        weights1[18238] <= 16'b1111111111111011;
        weights1[18239] <= 16'b1111111111110011;
        weights1[18240] <= 16'b0000000000000000;
        weights1[18241] <= 16'b1111111111110110;
        weights1[18242] <= 16'b1111111111111110;
        weights1[18243] <= 16'b0000000000000100;
        weights1[18244] <= 16'b1111111111111101;
        weights1[18245] <= 16'b1111111111111011;
        weights1[18246] <= 16'b0000000000001000;
        weights1[18247] <= 16'b1111111111111010;
        weights1[18248] <= 16'b1111111111110111;
        weights1[18249] <= 16'b0000000000010000;
        weights1[18250] <= 16'b0000000000010000;
        weights1[18251] <= 16'b0000000000001110;
        weights1[18252] <= 16'b0000000000000110;
        weights1[18253] <= 16'b1111111111111101;
        weights1[18254] <= 16'b0000000000001100;
        weights1[18255] <= 16'b0000000000001000;
        weights1[18256] <= 16'b1111111111111100;
        weights1[18257] <= 16'b1111111111111011;
        weights1[18258] <= 16'b1111111111111001;
        weights1[18259] <= 16'b1111111111110100;
        weights1[18260] <= 16'b1111111111111100;
        weights1[18261] <= 16'b1111111111110000;
        weights1[18262] <= 16'b1111111111111001;
        weights1[18263] <= 16'b0000000000011011;
        weights1[18264] <= 16'b1111111111111100;
        weights1[18265] <= 16'b1111111111111100;
        weights1[18266] <= 16'b1111111111111000;
        weights1[18267] <= 16'b1111111111111000;
        weights1[18268] <= 16'b0000000000001001;
        weights1[18269] <= 16'b0000000000001100;
        weights1[18270] <= 16'b1111111111111100;
        weights1[18271] <= 16'b0000000000001000;
        weights1[18272] <= 16'b1111111111111111;
        weights1[18273] <= 16'b1111111111111001;
        weights1[18274] <= 16'b0000000000000000;
        weights1[18275] <= 16'b0000000000001101;
        weights1[18276] <= 16'b0000000000000000;
        weights1[18277] <= 16'b1111111111111110;
        weights1[18278] <= 16'b0000000000001100;
        weights1[18279] <= 16'b0000000000000110;
        weights1[18280] <= 16'b1111111111111111;
        weights1[18281] <= 16'b1111111111110011;
        weights1[18282] <= 16'b0000000000010100;
        weights1[18283] <= 16'b0000000000000101;
        weights1[18284] <= 16'b1111111111111101;
        weights1[18285] <= 16'b1111111111110111;
        weights1[18286] <= 16'b1111111111110111;
        weights1[18287] <= 16'b1111111111101101;
        weights1[18288] <= 16'b1111111111110111;
        weights1[18289] <= 16'b1111111111110110;
        weights1[18290] <= 16'b0000000000000110;
        weights1[18291] <= 16'b0000000000010001;
        weights1[18292] <= 16'b0000000000010011;
        weights1[18293] <= 16'b0000000000010000;
        weights1[18294] <= 16'b1111111111100111;
        weights1[18295] <= 16'b1111111111101000;
        weights1[18296] <= 16'b1111111111101000;
        weights1[18297] <= 16'b1111111111111101;
        weights1[18298] <= 16'b1111111111111010;
        weights1[18299] <= 16'b0000000000000111;
        weights1[18300] <= 16'b0000000000000010;
        weights1[18301] <= 16'b0000000000000110;
        weights1[18302] <= 16'b1111111111110100;
        weights1[18303] <= 16'b1111111111110110;
        weights1[18304] <= 16'b0000000000000110;
        weights1[18305] <= 16'b0000000000001011;
        weights1[18306] <= 16'b1111111111111101;
        weights1[18307] <= 16'b0000000000011011;
        weights1[18308] <= 16'b0000000000000011;
        weights1[18309] <= 16'b0000000000010011;
        weights1[18310] <= 16'b0000000000001010;
        weights1[18311] <= 16'b0000000000000011;
        weights1[18312] <= 16'b1111111111111000;
        weights1[18313] <= 16'b0000000000000100;
        weights1[18314] <= 16'b0000000000000111;
        weights1[18315] <= 16'b1111111111110010;
        weights1[18316] <= 16'b1111111111110011;
        weights1[18317] <= 16'b0000000000000011;
        weights1[18318] <= 16'b1111111111111101;
        weights1[18319] <= 16'b1111111111111111;
        weights1[18320] <= 16'b0000000000010110;
        weights1[18321] <= 16'b0000000000000011;
        weights1[18322] <= 16'b0000000000010111;
        weights1[18323] <= 16'b0000000000000100;
        weights1[18324] <= 16'b1111111111110000;
        weights1[18325] <= 16'b1111111111111100;
        weights1[18326] <= 16'b1111111111110101;
        weights1[18327] <= 16'b1111111111111001;
        weights1[18328] <= 16'b1111111111110111;
        weights1[18329] <= 16'b0000000000000111;
        weights1[18330] <= 16'b1111111111110100;
        weights1[18331] <= 16'b1111111111111101;
        weights1[18332] <= 16'b0000000000010100;
        weights1[18333] <= 16'b1111111111111101;
        weights1[18334] <= 16'b1111111111101011;
        weights1[18335] <= 16'b0000000000001010;
        weights1[18336] <= 16'b0000000000010011;
        weights1[18337] <= 16'b1111111111100101;
        weights1[18338] <= 16'b0000000000000111;
        weights1[18339] <= 16'b1111111111111111;
        weights1[18340] <= 16'b1111111111111111;
        weights1[18341] <= 16'b0000000000000111;
        weights1[18342] <= 16'b0000000000000101;
        weights1[18343] <= 16'b0000000000000000;
        weights1[18344] <= 16'b1111111111111110;
        weights1[18345] <= 16'b1111111111111000;
        weights1[18346] <= 16'b0000000000001011;
        weights1[18347] <= 16'b0000000000000100;
        weights1[18348] <= 16'b1111111111111001;
        weights1[18349] <= 16'b1111111111111100;
        weights1[18350] <= 16'b1111111111110111;
        weights1[18351] <= 16'b0000000000001010;
        weights1[18352] <= 16'b0000000000000101;
        weights1[18353] <= 16'b1111111111101100;
        weights1[18354] <= 16'b1111111111111110;
        weights1[18355] <= 16'b1111111111101100;
        weights1[18356] <= 16'b1111111111110100;
        weights1[18357] <= 16'b1111111111111001;
        weights1[18358] <= 16'b0000000000001000;
        weights1[18359] <= 16'b0000000000000100;
        weights1[18360] <= 16'b1111111111111101;
        weights1[18361] <= 16'b1111111111101110;
        weights1[18362] <= 16'b0000000000010011;
        weights1[18363] <= 16'b0000000000010001;
        weights1[18364] <= 16'b1111111111111100;
        weights1[18365] <= 16'b1111111111111101;
        weights1[18366] <= 16'b0000000000001110;
        weights1[18367] <= 16'b0000000000001011;
        weights1[18368] <= 16'b0000000000000110;
        weights1[18369] <= 16'b0000000000000111;
        weights1[18370] <= 16'b0000000000000110;
        weights1[18371] <= 16'b0000000000001110;
        weights1[18372] <= 16'b0000000000010110;
        weights1[18373] <= 16'b0000000000010101;
        weights1[18374] <= 16'b1111111111111111;
        weights1[18375] <= 16'b0000000000011110;
        weights1[18376] <= 16'b0000000000001001;
        weights1[18377] <= 16'b1111111111110000;
        weights1[18378] <= 16'b1111111111110000;
        weights1[18379] <= 16'b0000000000000101;
        weights1[18380] <= 16'b1111111111100010;
        weights1[18381] <= 16'b1111111111100101;
        weights1[18382] <= 16'b1111111111011011;
        weights1[18383] <= 16'b1111111111101101;
        weights1[18384] <= 16'b1111111111100001;
        weights1[18385] <= 16'b1111111111110101;
        weights1[18386] <= 16'b1111111111110011;
        weights1[18387] <= 16'b1111111111101000;
        weights1[18388] <= 16'b0000000000001000;
        weights1[18389] <= 16'b1111111111110101;
        weights1[18390] <= 16'b1111111111111001;
        weights1[18391] <= 16'b1111111111110011;
        weights1[18392] <= 16'b0000000000000000;
        weights1[18393] <= 16'b0000000000001000;
        weights1[18394] <= 16'b0000000000001100;
        weights1[18395] <= 16'b1111111111111100;
        weights1[18396] <= 16'b1111111111111010;
        weights1[18397] <= 16'b1111111111111011;
        weights1[18398] <= 16'b1111111111111110;
        weights1[18399] <= 16'b0000000000000110;
        weights1[18400] <= 16'b0000000000010101;
        weights1[18401] <= 16'b1111111111111011;
        weights1[18402] <= 16'b1111111111101010;
        weights1[18403] <= 16'b1111111111101111;
        weights1[18404] <= 16'b0000000000000001;
        weights1[18405] <= 16'b0000000000001001;
        weights1[18406] <= 16'b1111111111110111;
        weights1[18407] <= 16'b1111111111101000;
        weights1[18408] <= 16'b1111111111100011;
        weights1[18409] <= 16'b1111111111100011;
        weights1[18410] <= 16'b1111111111101001;
        weights1[18411] <= 16'b1111111111100110;
        weights1[18412] <= 16'b1111111111011110;
        weights1[18413] <= 16'b1111111111110010;
        weights1[18414] <= 16'b0000000000000110;
        weights1[18415] <= 16'b0000000000001001;
        weights1[18416] <= 16'b0000000000001101;
        weights1[18417] <= 16'b0000000000001010;
        weights1[18418] <= 16'b0000000000010100;
        weights1[18419] <= 16'b1111111111110110;
        weights1[18420] <= 16'b0000000000010100;
        weights1[18421] <= 16'b0000000000010110;
        weights1[18422] <= 16'b1111111111111000;
        weights1[18423] <= 16'b1111111111011110;
        weights1[18424] <= 16'b1111111111110100;
        weights1[18425] <= 16'b1111111111101110;
        weights1[18426] <= 16'b1111111111110101;
        weights1[18427] <= 16'b1111111111111010;
        weights1[18428] <= 16'b0000000000000001;
        weights1[18429] <= 16'b1111111111110001;
        weights1[18430] <= 16'b0000000000001001;
        weights1[18431] <= 16'b1111111111100111;
        weights1[18432] <= 16'b1111111111110010;
        weights1[18433] <= 16'b1111111111101000;
        weights1[18434] <= 16'b1111111111011011;
        weights1[18435] <= 16'b1111111111010001;
        weights1[18436] <= 16'b1111111111001001;
        weights1[18437] <= 16'b0000000000000000;
        weights1[18438] <= 16'b1111111111110100;
        weights1[18439] <= 16'b1111111111110100;
        weights1[18440] <= 16'b1111111111110100;
        weights1[18441] <= 16'b1111111111110100;
        weights1[18442] <= 16'b1111111111010101;
        weights1[18443] <= 16'b1111111111101111;
        weights1[18444] <= 16'b0000000000000001;
        weights1[18445] <= 16'b0000000000100101;
        weights1[18446] <= 16'b0000000000010001;
        weights1[18447] <= 16'b0000000000011110;
        weights1[18448] <= 16'b0000000000101000;
        weights1[18449] <= 16'b0000000000010001;
        weights1[18450] <= 16'b1111111111101100;
        weights1[18451] <= 16'b1111111111010101;
        weights1[18452] <= 16'b1111111111110111;
        weights1[18453] <= 16'b1111111111101110;
        weights1[18454] <= 16'b1111111111100100;
        weights1[18455] <= 16'b1111111111011111;
        weights1[18456] <= 16'b1111111111100000;
        weights1[18457] <= 16'b1111111111100010;
        weights1[18458] <= 16'b1111111111101110;
        weights1[18459] <= 16'b1111111111101101;
        weights1[18460] <= 16'b1111111111010011;
        weights1[18461] <= 16'b1111111110110001;
        weights1[18462] <= 16'b1111111111001100;
        weights1[18463] <= 16'b1111111111010101;
        weights1[18464] <= 16'b1111111111111101;
        weights1[18465] <= 16'b1111111111111111;
        weights1[18466] <= 16'b0000000000000110;
        weights1[18467] <= 16'b1111111111111110;
        weights1[18468] <= 16'b1111111111100001;
        weights1[18469] <= 16'b1111111111101101;
        weights1[18470] <= 16'b0000000000000110;
        weights1[18471] <= 16'b1111111111101001;
        weights1[18472] <= 16'b1111111111111011;
        weights1[18473] <= 16'b0000000000010000;
        weights1[18474] <= 16'b0000000000101011;
        weights1[18475] <= 16'b0000000000101010;
        weights1[18476] <= 16'b0000000000001101;
        weights1[18477] <= 16'b1111111111000101;
        weights1[18478] <= 16'b1111111110110010;
        weights1[18479] <= 16'b1111111110110101;
        weights1[18480] <= 16'b1111111111101111;
        weights1[18481] <= 16'b1111111111101100;
        weights1[18482] <= 16'b1111111111010001;
        weights1[18483] <= 16'b1111111110111101;
        weights1[18484] <= 16'b1111111111010011;
        weights1[18485] <= 16'b1111111111010000;
        weights1[18486] <= 16'b1111111110111011;
        weights1[18487] <= 16'b1111111110111010;
        weights1[18488] <= 16'b1111111110011101;
        weights1[18489] <= 16'b1111111111001101;
        weights1[18490] <= 16'b1111111111010001;
        weights1[18491] <= 16'b1111111111111111;
        weights1[18492] <= 16'b0000000000010000;
        weights1[18493] <= 16'b0000000000010010;
        weights1[18494] <= 16'b0000000000010001;
        weights1[18495] <= 16'b0000000000010010;
        weights1[18496] <= 16'b1111111111110110;
        weights1[18497] <= 16'b1111111111101111;
        weights1[18498] <= 16'b1111111111110001;
        weights1[18499] <= 16'b1111111111110000;
        weights1[18500] <= 16'b1111111111111011;
        weights1[18501] <= 16'b0000000000001000;
        weights1[18502] <= 16'b1111111111111000;
        weights1[18503] <= 16'b1111111111001101;
        weights1[18504] <= 16'b1111111110110100;
        weights1[18505] <= 16'b1111111110010110;
        weights1[18506] <= 16'b1111111110101011;
        weights1[18507] <= 16'b1111111110110011;
        weights1[18508] <= 16'b1111111111101100;
        weights1[18509] <= 16'b1111111111011110;
        weights1[18510] <= 16'b1111111111001000;
        weights1[18511] <= 16'b1111111110110000;
        weights1[18512] <= 16'b1111111110111000;
        weights1[18513] <= 16'b1111111110100011;
        weights1[18514] <= 16'b1111111110010110;
        weights1[18515] <= 16'b1111111110011011;
        weights1[18516] <= 16'b1111111111010011;
        weights1[18517] <= 16'b1111111111110111;
        weights1[18518] <= 16'b0000000000000100;
        weights1[18519] <= 16'b0000000000011001;
        weights1[18520] <= 16'b0000000000011000;
        weights1[18521] <= 16'b0000000000010111;
        weights1[18522] <= 16'b0000000000000010;
        weights1[18523] <= 16'b0000000000011000;
        weights1[18524] <= 16'b0000000000000110;
        weights1[18525] <= 16'b1111111111110101;
        weights1[18526] <= 16'b1111111111011111;
        weights1[18527] <= 16'b1111111111010101;
        weights1[18528] <= 16'b1111111110110000;
        weights1[18529] <= 16'b1111111110101010;
        weights1[18530] <= 16'b1111111101111100;
        weights1[18531] <= 16'b1111111101101101;
        weights1[18532] <= 16'b1111111101111011;
        weights1[18533] <= 16'b1111111110100100;
        weights1[18534] <= 16'b1111111110100011;
        weights1[18535] <= 16'b1111111110110110;
        weights1[18536] <= 16'b1111111111101011;
        weights1[18537] <= 16'b1111111111011001;
        weights1[18538] <= 16'b1111111111001011;
        weights1[18539] <= 16'b1111111110111000;
        weights1[18540] <= 16'b1111111110110010;
        weights1[18541] <= 16'b1111111110100101;
        weights1[18542] <= 16'b1111111111010000;
        weights1[18543] <= 16'b1111111111100100;
        weights1[18544] <= 16'b1111111111111110;
        weights1[18545] <= 16'b0000000000011001;
        weights1[18546] <= 16'b0000000000011110;
        weights1[18547] <= 16'b0000000000100010;
        weights1[18548] <= 16'b0000000000000101;
        weights1[18549] <= 16'b0000000000010100;
        weights1[18550] <= 16'b0000000000000000;
        weights1[18551] <= 16'b0000000000001001;
        weights1[18552] <= 16'b1111111111111101;
        weights1[18553] <= 16'b1111111111100001;
        weights1[18554] <= 16'b1111111111010111;
        weights1[18555] <= 16'b1111111110110111;
        weights1[18556] <= 16'b1111111101111011;
        weights1[18557] <= 16'b1111111100111010;
        weights1[18558] <= 16'b1111111100101101;
        weights1[18559] <= 16'b1111111101011110;
        weights1[18560] <= 16'b1111111101110110;
        weights1[18561] <= 16'b1111111110100010;
        weights1[18562] <= 16'b1111111110100110;
        weights1[18563] <= 16'b1111111110110001;
        weights1[18564] <= 16'b1111111111101011;
        weights1[18565] <= 16'b1111111111100000;
        weights1[18566] <= 16'b1111111111010001;
        weights1[18567] <= 16'b1111111111010010;
        weights1[18568] <= 16'b1111111111001011;
        weights1[18569] <= 16'b1111111111011111;
        weights1[18570] <= 16'b1111111111100101;
        weights1[18571] <= 16'b0000000000010000;
        weights1[18572] <= 16'b0000000000011011;
        weights1[18573] <= 16'b0000000000011111;
        weights1[18574] <= 16'b1111111111111101;
        weights1[18575] <= 16'b0000000000010111;
        weights1[18576] <= 16'b0000000000010110;
        weights1[18577] <= 16'b0000000000010011;
        weights1[18578] <= 16'b0000000000010111;
        weights1[18579] <= 16'b1111111111111110;
        weights1[18580] <= 16'b0000000000000110;
        weights1[18581] <= 16'b1111111111111110;
        weights1[18582] <= 16'b1111111111011010;
        weights1[18583] <= 16'b1111111111000100;
        weights1[18584] <= 16'b1111111110000111;
        weights1[18585] <= 16'b1111111101101010;
        weights1[18586] <= 16'b1111111101101001;
        weights1[18587] <= 16'b1111111101111110;
        weights1[18588] <= 16'b1111111110000100;
        weights1[18589] <= 16'b1111111110011111;
        weights1[18590] <= 16'b1111111110100101;
        weights1[18591] <= 16'b1111111111000000;
        weights1[18592] <= 16'b1111111111101101;
        weights1[18593] <= 16'b1111111111100100;
        weights1[18594] <= 16'b1111111111011100;
        weights1[18595] <= 16'b1111111111100010;
        weights1[18596] <= 16'b1111111111111011;
        weights1[18597] <= 16'b0000000000000010;
        weights1[18598] <= 16'b0000000000100100;
        weights1[18599] <= 16'b0000000000100101;
        weights1[18600] <= 16'b0000000000001111;
        weights1[18601] <= 16'b0000000000011110;
        weights1[18602] <= 16'b0000000000100001;
        weights1[18603] <= 16'b0000000000001001;
        weights1[18604] <= 16'b0000000000000111;
        weights1[18605] <= 16'b0000000000010100;
        weights1[18606] <= 16'b0000000000010111;
        weights1[18607] <= 16'b0000000000010000;
        weights1[18608] <= 16'b0000000000000001;
        weights1[18609] <= 16'b0000000000010000;
        weights1[18610] <= 16'b1111111111110010;
        weights1[18611] <= 16'b1111111111011001;
        weights1[18612] <= 16'b0000000000000010;
        weights1[18613] <= 16'b1111111111011111;
        weights1[18614] <= 16'b1111111111001111;
        weights1[18615] <= 16'b1111111110101100;
        weights1[18616] <= 16'b1111111110110000;
        weights1[18617] <= 16'b1111111110110110;
        weights1[18618] <= 16'b1111111110111010;
        weights1[18619] <= 16'b1111111111001100;
        weights1[18620] <= 16'b1111111111110100;
        weights1[18621] <= 16'b1111111111110011;
        weights1[18622] <= 16'b1111111111111110;
        weights1[18623] <= 16'b0000000000000111;
        weights1[18624] <= 16'b0000000000001010;
        weights1[18625] <= 16'b0000000000011111;
        weights1[18626] <= 16'b0000000000101100;
        weights1[18627] <= 16'b0000000000000111;
        weights1[18628] <= 16'b0000000000010000;
        weights1[18629] <= 16'b0000000000001001;
        weights1[18630] <= 16'b0000000000011111;
        weights1[18631] <= 16'b0000000000100001;
        weights1[18632] <= 16'b0000000000101101;
        weights1[18633] <= 16'b0000000000100110;
        weights1[18634] <= 16'b0000000000001010;
        weights1[18635] <= 16'b0000000000111000;
        weights1[18636] <= 16'b0000000000100000;
        weights1[18637] <= 16'b0000000000100011;
        weights1[18638] <= 16'b0000000000111110;
        weights1[18639] <= 16'b0000000000101001;
        weights1[18640] <= 16'b0000000000101100;
        weights1[18641] <= 16'b0000000000101101;
        weights1[18642] <= 16'b0000000000100011;
        weights1[18643] <= 16'b0000000000001000;
        weights1[18644] <= 16'b1111111111011100;
        weights1[18645] <= 16'b1111111111010111;
        weights1[18646] <= 16'b1111111111011000;
        weights1[18647] <= 16'b1111111111100001;
        weights1[18648] <= 16'b0000000000000111;
        weights1[18649] <= 16'b0000000000001110;
        weights1[18650] <= 16'b0000000000001111;
        weights1[18651] <= 16'b0000000000010100;
        weights1[18652] <= 16'b0000000000010000;
        weights1[18653] <= 16'b0000000000100010;
        weights1[18654] <= 16'b0000000000001001;
        weights1[18655] <= 16'b0000000000000001;
        weights1[18656] <= 16'b0000000000011001;
        weights1[18657] <= 16'b0000000000010101;
        weights1[18658] <= 16'b0000000000011110;
        weights1[18659] <= 16'b0000000000011000;
        weights1[18660] <= 16'b0000000000101010;
        weights1[18661] <= 16'b0000000000110001;
        weights1[18662] <= 16'b0000000000100000;
        weights1[18663] <= 16'b0000000000101110;
        weights1[18664] <= 16'b0000000000100111;
        weights1[18665] <= 16'b0000000000101110;
        weights1[18666] <= 16'b0000000001001101;
        weights1[18667] <= 16'b0000000000110111;
        weights1[18668] <= 16'b0000000000111011;
        weights1[18669] <= 16'b0000000001010111;
        weights1[18670] <= 16'b0000000001000101;
        weights1[18671] <= 16'b0000000000100001;
        weights1[18672] <= 16'b0000000000010011;
        weights1[18673] <= 16'b1111111111110011;
        weights1[18674] <= 16'b1111111111111001;
        weights1[18675] <= 16'b1111111111110011;
        weights1[18676] <= 16'b0000000000001011;
        weights1[18677] <= 16'b0000000000011011;
        weights1[18678] <= 16'b0000000000011001;
        weights1[18679] <= 16'b0000000000010011;
        weights1[18680] <= 16'b0000000000100101;
        weights1[18681] <= 16'b0000000000010010;
        weights1[18682] <= 16'b0000000000000100;
        weights1[18683] <= 16'b0000000000001010;
        weights1[18684] <= 16'b0000000000011111;
        weights1[18685] <= 16'b0000000000001100;
        weights1[18686] <= 16'b0000000000011110;
        weights1[18687] <= 16'b0000000000010001;
        weights1[18688] <= 16'b0000000000011110;
        weights1[18689] <= 16'b0000000000100011;
        weights1[18690] <= 16'b0000000000011011;
        weights1[18691] <= 16'b0000000000100110;
        weights1[18692] <= 16'b0000000001000110;
        weights1[18693] <= 16'b0000000000010100;
        weights1[18694] <= 16'b0000000000100001;
        weights1[18695] <= 16'b0000000001001000;
        weights1[18696] <= 16'b0000000000111110;
        weights1[18697] <= 16'b0000000000101111;
        weights1[18698] <= 16'b0000000001010100;
        weights1[18699] <= 16'b0000000001000000;
        weights1[18700] <= 16'b0000000000101111;
        weights1[18701] <= 16'b0000000000011001;
        weights1[18702] <= 16'b0000000000001111;
        weights1[18703] <= 16'b0000000000001011;
        weights1[18704] <= 16'b0000000000000001;
        weights1[18705] <= 16'b0000000000000111;
        weights1[18706] <= 16'b0000000000000001;
        weights1[18707] <= 16'b0000000000000100;
        weights1[18708] <= 16'b0000000000001010;
        weights1[18709] <= 16'b0000000000010011;
        weights1[18710] <= 16'b1111111111111110;
        weights1[18711] <= 16'b1111111111111000;
        weights1[18712] <= 16'b0000000000001000;
        weights1[18713] <= 16'b0000000000010111;
        weights1[18714] <= 16'b0000000000000101;
        weights1[18715] <= 16'b0000000000011110;
        weights1[18716] <= 16'b0000000000100000;
        weights1[18717] <= 16'b0000000000010100;
        weights1[18718] <= 16'b0000000000010101;
        weights1[18719] <= 16'b0000000000011110;
        weights1[18720] <= 16'b0000000000000111;
        weights1[18721] <= 16'b0000000000110011;
        weights1[18722] <= 16'b0000000000101101;
        weights1[18723] <= 16'b0000000000100011;
        weights1[18724] <= 16'b0000000000100110;
        weights1[18725] <= 16'b0000000000101011;
        weights1[18726] <= 16'b0000000001011111;
        weights1[18727] <= 16'b0000000000110111;
        weights1[18728] <= 16'b0000000000101011;
        weights1[18729] <= 16'b0000000000101000;
        weights1[18730] <= 16'b0000000000011110;
        weights1[18731] <= 16'b0000000000001100;
        weights1[18732] <= 16'b0000000000000001;
        weights1[18733] <= 16'b0000000000000100;
        weights1[18734] <= 16'b0000000000000000;
        weights1[18735] <= 16'b0000000000001001;
        weights1[18736] <= 16'b0000000000010100;
        weights1[18737] <= 16'b0000000000011111;
        weights1[18738] <= 16'b0000000000010100;
        weights1[18739] <= 16'b0000000000010011;
        weights1[18740] <= 16'b0000000000001010;
        weights1[18741] <= 16'b0000000000001101;
        weights1[18742] <= 16'b0000000000001011;
        weights1[18743] <= 16'b1111111111110100;
        weights1[18744] <= 16'b0000000000001011;
        weights1[18745] <= 16'b0000000000010111;
        weights1[18746] <= 16'b0000000000001010;
        weights1[18747] <= 16'b0000000000011000;
        weights1[18748] <= 16'b0000000000001000;
        weights1[18749] <= 16'b0000000000011000;
        weights1[18750] <= 16'b0000000000010110;
        weights1[18751] <= 16'b0000000000100011;
        weights1[18752] <= 16'b0000000000110010;
        weights1[18753] <= 16'b0000000000001101;
        weights1[18754] <= 16'b0000000000101111;
        weights1[18755] <= 16'b0000000000110111;
        weights1[18756] <= 16'b0000000000110010;
        weights1[18757] <= 16'b0000000000100100;
        weights1[18758] <= 16'b0000000000011001;
        weights1[18759] <= 16'b0000000000000111;
        weights1[18760] <= 16'b0000000000000000;
        weights1[18761] <= 16'b1111111111111111;
        weights1[18762] <= 16'b0000000000000110;
        weights1[18763] <= 16'b0000000000001110;
        weights1[18764] <= 16'b0000000000000000;
        weights1[18765] <= 16'b0000000000000100;
        weights1[18766] <= 16'b0000000000011011;
        weights1[18767] <= 16'b0000000000011001;
        weights1[18768] <= 16'b0000000000010100;
        weights1[18769] <= 16'b0000000000010100;
        weights1[18770] <= 16'b0000000000000010;
        weights1[18771] <= 16'b0000000000010000;
        weights1[18772] <= 16'b0000000000001011;
        weights1[18773] <= 16'b0000000000000101;
        weights1[18774] <= 16'b0000000000001111;
        weights1[18775] <= 16'b0000000000000111;
        weights1[18776] <= 16'b0000000000010110;
        weights1[18777] <= 16'b0000000000000010;
        weights1[18778] <= 16'b0000000000001111;
        weights1[18779] <= 16'b0000000000001111;
        weights1[18780] <= 16'b0000000000001110;
        weights1[18781] <= 16'b0000000000011010;
        weights1[18782] <= 16'b0000000000111110;
        weights1[18783] <= 16'b0000000000110001;
        weights1[18784] <= 16'b0000000000101010;
        weights1[18785] <= 16'b0000000000010010;
        weights1[18786] <= 16'b0000000000001011;
        weights1[18787] <= 16'b0000000000000100;
        weights1[18788] <= 16'b0000000000000010;
        weights1[18789] <= 16'b1111111111111111;
        weights1[18790] <= 16'b1111111111111111;
        weights1[18791] <= 16'b0000000000000001;
        weights1[18792] <= 16'b1111111111111001;
        weights1[18793] <= 16'b0000000000001010;
        weights1[18794] <= 16'b0000000000010000;
        weights1[18795] <= 16'b1111111111111101;
        weights1[18796] <= 16'b0000000000001111;
        weights1[18797] <= 16'b0000000000001011;
        weights1[18798] <= 16'b1111111111111011;
        weights1[18799] <= 16'b0000000000000110;
        weights1[18800] <= 16'b1111111111111110;
        weights1[18801] <= 16'b1111111111111111;
        weights1[18802] <= 16'b1111111111111011;
        weights1[18803] <= 16'b0000000000010011;
        weights1[18804] <= 16'b0000000000010000;
        weights1[18805] <= 16'b0000000000010110;
        weights1[18806] <= 16'b0000000000000110;
        weights1[18807] <= 16'b1111111111111100;
        weights1[18808] <= 16'b0000000000010001;
        weights1[18809] <= 16'b0000000000101001;
        weights1[18810] <= 16'b0000000000100110;
        weights1[18811] <= 16'b0000000000011101;
        weights1[18812] <= 16'b0000000000010111;
        weights1[18813] <= 16'b0000000000001000;
        weights1[18814] <= 16'b0000000000000100;
        weights1[18815] <= 16'b0000000000000100;
        weights1[18816] <= 16'b0000000000000000;
        weights1[18817] <= 16'b0000000000000000;
        weights1[18818] <= 16'b0000000000000001;
        weights1[18819] <= 16'b0000000000000010;
        weights1[18820] <= 16'b0000000000000111;
        weights1[18821] <= 16'b0000000000000101;
        weights1[18822] <= 16'b0000000000000101;
        weights1[18823] <= 16'b1111111111110000;
        weights1[18824] <= 16'b1111111111011100;
        weights1[18825] <= 16'b1111111111001001;
        weights1[18826] <= 16'b1111111110110111;
        weights1[18827] <= 16'b1111111110111010;
        weights1[18828] <= 16'b1111111111001111;
        weights1[18829] <= 16'b1111111111110011;
        weights1[18830] <= 16'b0000000000011001;
        weights1[18831] <= 16'b0000000000100011;
        weights1[18832] <= 16'b0000000000100101;
        weights1[18833] <= 16'b0000000000011110;
        weights1[18834] <= 16'b1111111111111110;
        weights1[18835] <= 16'b1111111111011011;
        weights1[18836] <= 16'b1111111111001000;
        weights1[18837] <= 16'b1111111111000011;
        weights1[18838] <= 16'b1111111111001100;
        weights1[18839] <= 16'b1111111111011011;
        weights1[18840] <= 16'b1111111111110111;
        weights1[18841] <= 16'b0000000000000011;
        weights1[18842] <= 16'b0000000000000010;
        weights1[18843] <= 16'b1111111111111111;
        weights1[18844] <= 16'b0000000000000000;
        weights1[18845] <= 16'b0000000000000000;
        weights1[18846] <= 16'b0000000000000011;
        weights1[18847] <= 16'b0000000000000111;
        weights1[18848] <= 16'b0000000000001000;
        weights1[18849] <= 16'b0000000000000101;
        weights1[18850] <= 16'b1111111111111101;
        weights1[18851] <= 16'b1111111111101101;
        weights1[18852] <= 16'b1111111111010010;
        weights1[18853] <= 16'b1111111110110011;
        weights1[18854] <= 16'b1111111110100000;
        weights1[18855] <= 16'b1111111110101011;
        weights1[18856] <= 16'b1111111111011000;
        weights1[18857] <= 16'b0000000000000100;
        weights1[18858] <= 16'b0000000000100100;
        weights1[18859] <= 16'b0000000000101110;
        weights1[18860] <= 16'b0000000000011100;
        weights1[18861] <= 16'b0000000000000111;
        weights1[18862] <= 16'b1111111111011111;
        weights1[18863] <= 16'b1111111110101110;
        weights1[18864] <= 16'b1111111110010111;
        weights1[18865] <= 16'b1111111110101100;
        weights1[18866] <= 16'b1111111111000011;
        weights1[18867] <= 16'b1111111111010110;
        weights1[18868] <= 16'b1111111111110101;
        weights1[18869] <= 16'b0000000000000010;
        weights1[18870] <= 16'b0000000000000111;
        weights1[18871] <= 16'b0000000000000011;
        weights1[18872] <= 16'b0000000000000000;
        weights1[18873] <= 16'b0000000000000001;
        weights1[18874] <= 16'b0000000000000000;
        weights1[18875] <= 16'b0000000000001010;
        weights1[18876] <= 16'b0000000000001001;
        weights1[18877] <= 16'b0000000000001110;
        weights1[18878] <= 16'b0000000000000001;
        weights1[18879] <= 16'b1111111111110010;
        weights1[18880] <= 16'b1111111110111011;
        weights1[18881] <= 16'b1111111110011110;
        weights1[18882] <= 16'b1111111110000101;
        weights1[18883] <= 16'b1111111110010101;
        weights1[18884] <= 16'b1111111111100111;
        weights1[18885] <= 16'b0000000000101110;
        weights1[18886] <= 16'b0000000000101111;
        weights1[18887] <= 16'b0000000000101100;
        weights1[18888] <= 16'b0000000000101010;
        weights1[18889] <= 16'b0000000000010100;
        weights1[18890] <= 16'b1111111111010000;
        weights1[18891] <= 16'b1111111110001011;
        weights1[18892] <= 16'b1111111101110111;
        weights1[18893] <= 16'b1111111110011000;
        weights1[18894] <= 16'b1111111111001011;
        weights1[18895] <= 16'b1111111111100110;
        weights1[18896] <= 16'b1111111111110101;
        weights1[18897] <= 16'b0000000000000010;
        weights1[18898] <= 16'b0000000000000011;
        weights1[18899] <= 16'b0000000000000100;
        weights1[18900] <= 16'b0000000000000000;
        weights1[18901] <= 16'b0000000000000001;
        weights1[18902] <= 16'b0000000000010000;
        weights1[18903] <= 16'b0000000000010110;
        weights1[18904] <= 16'b0000000000011110;
        weights1[18905] <= 16'b0000000000011111;
        weights1[18906] <= 16'b0000000000010100;
        weights1[18907] <= 16'b1111111111111011;
        weights1[18908] <= 16'b1111111110111001;
        weights1[18909] <= 16'b1111111110011000;
        weights1[18910] <= 16'b1111111110000011;
        weights1[18911] <= 16'b1111111110010110;
        weights1[18912] <= 16'b1111111111011111;
        weights1[18913] <= 16'b0000000000101000;
        weights1[18914] <= 16'b0000000000111111;
        weights1[18915] <= 16'b0000000000101111;
        weights1[18916] <= 16'b0000000000001110;
        weights1[18917] <= 16'b0000000000100000;
        weights1[18918] <= 16'b1111111110111010;
        weights1[18919] <= 16'b1111111101100001;
        weights1[18920] <= 16'b1111111101100111;
        weights1[18921] <= 16'b1111111110011111;
        weights1[18922] <= 16'b1111111111001000;
        weights1[18923] <= 16'b1111111111101001;
        weights1[18924] <= 16'b0000000000000111;
        weights1[18925] <= 16'b0000000000010111;
        weights1[18926] <= 16'b0000000000010101;
        weights1[18927] <= 16'b0000000000001000;
        weights1[18928] <= 16'b0000000000000000;
        weights1[18929] <= 16'b0000000000001000;
        weights1[18930] <= 16'b0000000000010101;
        weights1[18931] <= 16'b0000000000011110;
        weights1[18932] <= 16'b0000000000100110;
        weights1[18933] <= 16'b0000000000100001;
        weights1[18934] <= 16'b0000000000010100;
        weights1[18935] <= 16'b1111111111111111;
        weights1[18936] <= 16'b1111111110111010;
        weights1[18937] <= 16'b1111111101111111;
        weights1[18938] <= 16'b1111111101010101;
        weights1[18939] <= 16'b1111111110100110;
        weights1[18940] <= 16'b1111111111011110;
        weights1[18941] <= 16'b0000000001001011;
        weights1[18942] <= 16'b0000000000101110;
        weights1[18943] <= 16'b0000000000100001;
        weights1[18944] <= 16'b0000000000110101;
        weights1[18945] <= 16'b1111111111011110;
        weights1[18946] <= 16'b1111111110011001;
        weights1[18947] <= 16'b1111111101000111;
        weights1[18948] <= 16'b1111111101010111;
        weights1[18949] <= 16'b1111111110110100;
        weights1[18950] <= 16'b1111111111111100;
        weights1[18951] <= 16'b0000000000001011;
        weights1[18952] <= 16'b0000000000100001;
        weights1[18953] <= 16'b0000000000101100;
        weights1[18954] <= 16'b0000000000100000;
        weights1[18955] <= 16'b0000000000010010;
        weights1[18956] <= 16'b0000000000000010;
        weights1[18957] <= 16'b0000000000000110;
        weights1[18958] <= 16'b0000000000001010;
        weights1[18959] <= 16'b0000000000011010;
        weights1[18960] <= 16'b0000000000100011;
        weights1[18961] <= 16'b0000000000100101;
        weights1[18962] <= 16'b0000000000011101;
        weights1[18963] <= 16'b0000000000001110;
        weights1[18964] <= 16'b1111111111010001;
        weights1[18965] <= 16'b1111111110011011;
        weights1[18966] <= 16'b1111111101100001;
        weights1[18967] <= 16'b1111111111000101;
        weights1[18968] <= 16'b0000000000010010;
        weights1[18969] <= 16'b0000000000101000;
        weights1[18970] <= 16'b0000000000111000;
        weights1[18971] <= 16'b0000000000111001;
        weights1[18972] <= 16'b0000000000000010;
        weights1[18973] <= 16'b1111111111000100;
        weights1[18974] <= 16'b1111111101100100;
        weights1[18975] <= 16'b1111111101001100;
        weights1[18976] <= 16'b1111111101111101;
        weights1[18977] <= 16'b1111111111111011;
        weights1[18978] <= 16'b0000000000011011;
        weights1[18979] <= 16'b0000000000010011;
        weights1[18980] <= 16'b0000000000011000;
        weights1[18981] <= 16'b0000000000101100;
        weights1[18982] <= 16'b0000000000010101;
        weights1[18983] <= 16'b0000000000010110;
        weights1[18984] <= 16'b1111111111111100;
        weights1[18985] <= 16'b0000000000000011;
        weights1[18986] <= 16'b0000000000000011;
        weights1[18987] <= 16'b0000000000000010;
        weights1[18988] <= 16'b0000000000010101;
        weights1[18989] <= 16'b0000000000101100;
        weights1[18990] <= 16'b0000000000101101;
        weights1[18991] <= 16'b0000000000100101;
        weights1[18992] <= 16'b1111111111011001;
        weights1[18993] <= 16'b1111111101111010;
        weights1[18994] <= 16'b1111111101110100;
        weights1[18995] <= 16'b1111111111110110;
        weights1[18996] <= 16'b0000000000001001;
        weights1[18997] <= 16'b0000000000100010;
        weights1[18998] <= 16'b0000000000100001;
        weights1[18999] <= 16'b0000000000100100;
        weights1[19000] <= 16'b0000000000001001;
        weights1[19001] <= 16'b1111111110111111;
        weights1[19002] <= 16'b1111111101010001;
        weights1[19003] <= 16'b1111111101010010;
        weights1[19004] <= 16'b1111111111011001;
        weights1[19005] <= 16'b0000000000110101;
        weights1[19006] <= 16'b0000000000101100;
        weights1[19007] <= 16'b0000000000110111;
        weights1[19008] <= 16'b0000000000011011;
        weights1[19009] <= 16'b0000000000011010;
        weights1[19010] <= 16'b0000000000011011;
        weights1[19011] <= 16'b0000000000011101;
        weights1[19012] <= 16'b0000000000000011;
        weights1[19013] <= 16'b1111111111111111;
        weights1[19014] <= 16'b0000000000000100;
        weights1[19015] <= 16'b0000000000001001;
        weights1[19016] <= 16'b1111111111111101;
        weights1[19017] <= 16'b0000000000011100;
        weights1[19018] <= 16'b0000000000100110;
        weights1[19019] <= 16'b0000000000110110;
        weights1[19020] <= 16'b1111111111001001;
        weights1[19021] <= 16'b1111111110011101;
        weights1[19022] <= 16'b1111111110110011;
        weights1[19023] <= 16'b1111111111101101;
        weights1[19024] <= 16'b0000000000000110;
        weights1[19025] <= 16'b0000000000100010;
        weights1[19026] <= 16'b0000000000110000;
        weights1[19027] <= 16'b0000000000011001;
        weights1[19028] <= 16'b1111111111110001;
        weights1[19029] <= 16'b1111111110100000;
        weights1[19030] <= 16'b1111111101010011;
        weights1[19031] <= 16'b1111111110100011;
        weights1[19032] <= 16'b0000000000000001;
        weights1[19033] <= 16'b0000000000101101;
        weights1[19034] <= 16'b0000000000100000;
        weights1[19035] <= 16'b0000000000101000;
        weights1[19036] <= 16'b0000000000011000;
        weights1[19037] <= 16'b0000000000000000;
        weights1[19038] <= 16'b0000000000001110;
        weights1[19039] <= 16'b0000000000001000;
        weights1[19040] <= 16'b0000000000000001;
        weights1[19041] <= 16'b1111111111111000;
        weights1[19042] <= 16'b1111111111111001;
        weights1[19043] <= 16'b1111111111111100;
        weights1[19044] <= 16'b0000000000001111;
        weights1[19045] <= 16'b0000000000011001;
        weights1[19046] <= 16'b0000000000011011;
        weights1[19047] <= 16'b0000000000100100;
        weights1[19048] <= 16'b1111111111011010;
        weights1[19049] <= 16'b1111111111000001;
        weights1[19050] <= 16'b1111111111001101;
        weights1[19051] <= 16'b1111111111001111;
        weights1[19052] <= 16'b0000000000010101;
        weights1[19053] <= 16'b0000000000100001;
        weights1[19054] <= 16'b0000000000101010;
        weights1[19055] <= 16'b0000000000010010;
        weights1[19056] <= 16'b1111111111111101;
        weights1[19057] <= 16'b1111111110001101;
        weights1[19058] <= 16'b1111111100111100;
        weights1[19059] <= 16'b1111111111110011;
        weights1[19060] <= 16'b0000000000111111;
        weights1[19061] <= 16'b0000000000010001;
        weights1[19062] <= 16'b0000000000011111;
        weights1[19063] <= 16'b0000000000000101;
        weights1[19064] <= 16'b0000000000001100;
        weights1[19065] <= 16'b0000000000011001;
        weights1[19066] <= 16'b0000000000001101;
        weights1[19067] <= 16'b0000000000001000;
        weights1[19068] <= 16'b1111111111111011;
        weights1[19069] <= 16'b1111111111111010;
        weights1[19070] <= 16'b0000000000000110;
        weights1[19071] <= 16'b1111111111111000;
        weights1[19072] <= 16'b1111111111101111;
        weights1[19073] <= 16'b0000000000011111;
        weights1[19074] <= 16'b0000000000110100;
        weights1[19075] <= 16'b0000000000100100;
        weights1[19076] <= 16'b1111111111101000;
        weights1[19077] <= 16'b1111111111001011;
        weights1[19078] <= 16'b1111111111000101;
        weights1[19079] <= 16'b0000000000000000;
        weights1[19080] <= 16'b0000000000000011;
        weights1[19081] <= 16'b0000000000011000;
        weights1[19082] <= 16'b0000000000100000;
        weights1[19083] <= 16'b0000000000010000;
        weights1[19084] <= 16'b1111111111110011;
        weights1[19085] <= 16'b1111111110000010;
        weights1[19086] <= 16'b1111111110110110;
        weights1[19087] <= 16'b0000000000011000;
        weights1[19088] <= 16'b0000000000011110;
        weights1[19089] <= 16'b0000000000100111;
        weights1[19090] <= 16'b0000000000000001;
        weights1[19091] <= 16'b0000000000010101;
        weights1[19092] <= 16'b0000000000001100;
        weights1[19093] <= 16'b0000000000100100;
        weights1[19094] <= 16'b0000000000001111;
        weights1[19095] <= 16'b0000000000010000;
        weights1[19096] <= 16'b1111111111111100;
        weights1[19097] <= 16'b0000000000000001;
        weights1[19098] <= 16'b1111111111110101;
        weights1[19099] <= 16'b0000000000000011;
        weights1[19100] <= 16'b1111111111101000;
        weights1[19101] <= 16'b0000000000000010;
        weights1[19102] <= 16'b0000000000001110;
        weights1[19103] <= 16'b0000000000011101;
        weights1[19104] <= 16'b0000000000001001;
        weights1[19105] <= 16'b1111111111011100;
        weights1[19106] <= 16'b1111111111011111;
        weights1[19107] <= 16'b1111111111101000;
        weights1[19108] <= 16'b1111111111111110;
        weights1[19109] <= 16'b0000000000010011;
        weights1[19110] <= 16'b0000000000001101;
        weights1[19111] <= 16'b0000000000010011;
        weights1[19112] <= 16'b1111111111100010;
        weights1[19113] <= 16'b1111111110100010;
        weights1[19114] <= 16'b1111111111010101;
        weights1[19115] <= 16'b0000000000001110;
        weights1[19116] <= 16'b0000000000100110;
        weights1[19117] <= 16'b0000000000001001;
        weights1[19118] <= 16'b0000000000011100;
        weights1[19119] <= 16'b0000000000000010;
        weights1[19120] <= 16'b0000000000000111;
        weights1[19121] <= 16'b0000000000011100;
        weights1[19122] <= 16'b0000000000010100;
        weights1[19123] <= 16'b1111111111110110;
        weights1[19124] <= 16'b1111111111111111;
        weights1[19125] <= 16'b0000000000000100;
        weights1[19126] <= 16'b1111111111111100;
        weights1[19127] <= 16'b0000000000000100;
        weights1[19128] <= 16'b1111111111111110;
        weights1[19129] <= 16'b1111111111111110;
        weights1[19130] <= 16'b0000000000001100;
        weights1[19131] <= 16'b0000000000001101;
        weights1[19132] <= 16'b1111111111111000;
        weights1[19133] <= 16'b1111111111101010;
        weights1[19134] <= 16'b1111111111100100;
        weights1[19135] <= 16'b1111111111110110;
        weights1[19136] <= 16'b1111111111111110;
        weights1[19137] <= 16'b1111111111111010;
        weights1[19138] <= 16'b0000000000001011;
        weights1[19139] <= 16'b0000000000000011;
        weights1[19140] <= 16'b1111111111011000;
        weights1[19141] <= 16'b1111111111011100;
        weights1[19142] <= 16'b1111111111100101;
        weights1[19143] <= 16'b0000000000100101;
        weights1[19144] <= 16'b0000000000001011;
        weights1[19145] <= 16'b0000000000010110;
        weights1[19146] <= 16'b0000000000001000;
        weights1[19147] <= 16'b0000000000001001;
        weights1[19148] <= 16'b0000000000000010;
        weights1[19149] <= 16'b0000000000011010;
        weights1[19150] <= 16'b0000000000000000;
        weights1[19151] <= 16'b1111111111110110;
        weights1[19152] <= 16'b1111111111111011;
        weights1[19153] <= 16'b1111111111111101;
        weights1[19154] <= 16'b0000000000001111;
        weights1[19155] <= 16'b0000000000001000;
        weights1[19156] <= 16'b0000000000000111;
        weights1[19157] <= 16'b1111111111101111;
        weights1[19158] <= 16'b1111111111110100;
        weights1[19159] <= 16'b0000000000000010;
        weights1[19160] <= 16'b0000000000010110;
        weights1[19161] <= 16'b1111111111110000;
        weights1[19162] <= 16'b0000000000001100;
        weights1[19163] <= 16'b1111111111110010;
        weights1[19164] <= 16'b1111111111111101;
        weights1[19165] <= 16'b1111111111111111;
        weights1[19166] <= 16'b0000000000001001;
        weights1[19167] <= 16'b1111111111111111;
        weights1[19168] <= 16'b1111111111001111;
        weights1[19169] <= 16'b1111111111101001;
        weights1[19170] <= 16'b1111111111111010;
        weights1[19171] <= 16'b0000000000001000;
        weights1[19172] <= 16'b0000000000000100;
        weights1[19173] <= 16'b0000000000010000;
        weights1[19174] <= 16'b1111111111110011;
        weights1[19175] <= 16'b0000000000001001;
        weights1[19176] <= 16'b1111111111110000;
        weights1[19177] <= 16'b0000000000000100;
        weights1[19178] <= 16'b1111111111101001;
        weights1[19179] <= 16'b1111111111100110;
        weights1[19180] <= 16'b1111111111111100;
        weights1[19181] <= 16'b1111111111111111;
        weights1[19182] <= 16'b1111111111111110;
        weights1[19183] <= 16'b1111111111111111;
        weights1[19184] <= 16'b0000000000001001;
        weights1[19185] <= 16'b0000000000000011;
        weights1[19186] <= 16'b1111111111111101;
        weights1[19187] <= 16'b0000000000000011;
        weights1[19188] <= 16'b0000000000001000;
        weights1[19189] <= 16'b1111111111101010;
        weights1[19190] <= 16'b0000000000000010;
        weights1[19191] <= 16'b1111111111101110;
        weights1[19192] <= 16'b1111111111111111;
        weights1[19193] <= 16'b0000000000001000;
        weights1[19194] <= 16'b1111111111111001;
        weights1[19195] <= 16'b1111111111110010;
        weights1[19196] <= 16'b1111111111101011;
        weights1[19197] <= 16'b0000000000001001;
        weights1[19198] <= 16'b0000000000001001;
        weights1[19199] <= 16'b0000000000001101;
        weights1[19200] <= 16'b0000000000011011;
        weights1[19201] <= 16'b0000000000000100;
        weights1[19202] <= 16'b0000000000001101;
        weights1[19203] <= 16'b0000000000001010;
        weights1[19204] <= 16'b1111111111111001;
        weights1[19205] <= 16'b1111111111010000;
        weights1[19206] <= 16'b1111111111011100;
        weights1[19207] <= 16'b1111111111100100;
        weights1[19208] <= 16'b1111111111111010;
        weights1[19209] <= 16'b0000000000000011;
        weights1[19210] <= 16'b1111111111111110;
        weights1[19211] <= 16'b0000000000000100;
        weights1[19212] <= 16'b0000000000000011;
        weights1[19213] <= 16'b0000000000011011;
        weights1[19214] <= 16'b0000000000001101;
        weights1[19215] <= 16'b1111111111111010;
        weights1[19216] <= 16'b0000000000000111;
        weights1[19217] <= 16'b0000000000000110;
        weights1[19218] <= 16'b0000000000001101;
        weights1[19219] <= 16'b1111111111111000;
        weights1[19220] <= 16'b1111111111111101;
        weights1[19221] <= 16'b0000000000000010;
        weights1[19222] <= 16'b0000000000001000;
        weights1[19223] <= 16'b1111111111101100;
        weights1[19224] <= 16'b0000000000000011;
        weights1[19225] <= 16'b1111111111111110;
        weights1[19226] <= 16'b0000000000010000;
        weights1[19227] <= 16'b1111111111101110;
        weights1[19228] <= 16'b0000000000001010;
        weights1[19229] <= 16'b1111111111111101;
        weights1[19230] <= 16'b0000000000001110;
        weights1[19231] <= 16'b1111111111110010;
        weights1[19232] <= 16'b1111111111100110;
        weights1[19233] <= 16'b0000000000000010;
        weights1[19234] <= 16'b0000000000000000;
        weights1[19235] <= 16'b1111111111111010;
        weights1[19236] <= 16'b0000000000000010;
        weights1[19237] <= 16'b0000000000000011;
        weights1[19238] <= 16'b1111111111110111;
        weights1[19239] <= 16'b1111111111111101;
        weights1[19240] <= 16'b1111111111110011;
        weights1[19241] <= 16'b1111111111111010;
        weights1[19242] <= 16'b1111111111110110;
        weights1[19243] <= 16'b0000000000000111;
        weights1[19244] <= 16'b0000000000000110;
        weights1[19245] <= 16'b0000000000000001;
        weights1[19246] <= 16'b1111111111111110;
        weights1[19247] <= 16'b1111111111111101;
        weights1[19248] <= 16'b1111111111111110;
        weights1[19249] <= 16'b1111111111110111;
        weights1[19250] <= 16'b0000000000001110;
        weights1[19251] <= 16'b0000000000000111;
        weights1[19252] <= 16'b0000000000000101;
        weights1[19253] <= 16'b1111111111110111;
        weights1[19254] <= 16'b0000000000011000;
        weights1[19255] <= 16'b1111111111111100;
        weights1[19256] <= 16'b0000000000000101;
        weights1[19257] <= 16'b1111111111111000;
        weights1[19258] <= 16'b1111111111110000;
        weights1[19259] <= 16'b0000000000001101;
        weights1[19260] <= 16'b0000000000000000;
        weights1[19261] <= 16'b1111111111111110;
        weights1[19262] <= 16'b1111111111111101;
        weights1[19263] <= 16'b1111111111111010;
        weights1[19264] <= 16'b1111111111111010;
        weights1[19265] <= 16'b1111111111110110;
        weights1[19266] <= 16'b0000000000000001;
        weights1[19267] <= 16'b0000000000000100;
        weights1[19268] <= 16'b0000000000000000;
        weights1[19269] <= 16'b0000000000010001;
        weights1[19270] <= 16'b0000000000000111;
        weights1[19271] <= 16'b1111111111111001;
        weights1[19272] <= 16'b0000000000001101;
        weights1[19273] <= 16'b1111111111101111;
        weights1[19274] <= 16'b0000000000000100;
        weights1[19275] <= 16'b0000000000000010;
        weights1[19276] <= 16'b1111111111110110;
        weights1[19277] <= 16'b1111111111111100;
        weights1[19278] <= 16'b0000000000000010;
        weights1[19279] <= 16'b0000000000001011;
        weights1[19280] <= 16'b1111111111110010;
        weights1[19281] <= 16'b1111111111110111;
        weights1[19282] <= 16'b0000000000001010;
        weights1[19283] <= 16'b1111111111100110;
        weights1[19284] <= 16'b0000000000000000;
        weights1[19285] <= 16'b1111111111111010;
        weights1[19286] <= 16'b1111111111100110;
        weights1[19287] <= 16'b1111111111111001;
        weights1[19288] <= 16'b1111111111111010;
        weights1[19289] <= 16'b1111111111111011;
        weights1[19290] <= 16'b0000000000000011;
        weights1[19291] <= 16'b1111111111110111;
        weights1[19292] <= 16'b1111111111110110;
        weights1[19293] <= 16'b1111111111111100;
        weights1[19294] <= 16'b0000000000001111;
        weights1[19295] <= 16'b1111111111111100;
        weights1[19296] <= 16'b0000000000001110;
        weights1[19297] <= 16'b0000000000000011;
        weights1[19298] <= 16'b0000000000000110;
        weights1[19299] <= 16'b0000000000000100;
        weights1[19300] <= 16'b1111111111111110;
        weights1[19301] <= 16'b0000000000001010;
        weights1[19302] <= 16'b0000000000000111;
        weights1[19303] <= 16'b1111111111110101;
        weights1[19304] <= 16'b1111111111111000;
        weights1[19305] <= 16'b0000000000001110;
        weights1[19306] <= 16'b0000000000000101;
        weights1[19307] <= 16'b0000000000001111;
        weights1[19308] <= 16'b0000000000001111;
        weights1[19309] <= 16'b1111111111111010;
        weights1[19310] <= 16'b0000000000000101;
        weights1[19311] <= 16'b0000000000011100;
        weights1[19312] <= 16'b1111111111101111;
        weights1[19313] <= 16'b0000000000000001;
        weights1[19314] <= 16'b0000000000000110;
        weights1[19315] <= 16'b0000000000001011;
        weights1[19316] <= 16'b0000000000000001;
        weights1[19317] <= 16'b1111111111101110;
        weights1[19318] <= 16'b0000000000000111;
        weights1[19319] <= 16'b0000000000001101;
        weights1[19320] <= 16'b1111111111111001;
        weights1[19321] <= 16'b1111111111110001;
        weights1[19322] <= 16'b0000000000001100;
        weights1[19323] <= 16'b0000000000000101;
        weights1[19324] <= 16'b0000000000000111;
        weights1[19325] <= 16'b0000000000000111;
        weights1[19326] <= 16'b1111111111101110;
        weights1[19327] <= 16'b1111111111111010;
        weights1[19328] <= 16'b0000000000001011;
        weights1[19329] <= 16'b1111111111101111;
        weights1[19330] <= 16'b0000000000000000;
        weights1[19331] <= 16'b1111111111111100;
        weights1[19332] <= 16'b0000000000000111;
        weights1[19333] <= 16'b0000000000001000;
        weights1[19334] <= 16'b0000000000001011;
        weights1[19335] <= 16'b0000000000000001;
        weights1[19336] <= 16'b1111111111111110;
        weights1[19337] <= 16'b0000000000000000;
        weights1[19338] <= 16'b1111111111110111;
        weights1[19339] <= 16'b0000000000000111;
        weights1[19340] <= 16'b0000000000000100;
        weights1[19341] <= 16'b0000000000000110;
        weights1[19342] <= 16'b1111111111111010;
        weights1[19343] <= 16'b0000000000010011;
        weights1[19344] <= 16'b1111111111111010;
        weights1[19345] <= 16'b1111111111111100;
        weights1[19346] <= 16'b1111111111111110;
        weights1[19347] <= 16'b0000000000000001;
        weights1[19348] <= 16'b1111111111111110;
        weights1[19349] <= 16'b1111111111110111;
        weights1[19350] <= 16'b1111111111111111;
        weights1[19351] <= 16'b0000000000010011;
        weights1[19352] <= 16'b0000000000000101;
        weights1[19353] <= 16'b1111111111110110;
        weights1[19354] <= 16'b0000000000001011;
        weights1[19355] <= 16'b0000000000000111;
        weights1[19356] <= 16'b1111111111110110;
        weights1[19357] <= 16'b1111111111101111;
        weights1[19358] <= 16'b1111111111111101;
        weights1[19359] <= 16'b1111111111111100;
        weights1[19360] <= 16'b0000000000001011;
        weights1[19361] <= 16'b0000000000000000;
        weights1[19362] <= 16'b0000000000010100;
        weights1[19363] <= 16'b1111111111110100;
        weights1[19364] <= 16'b0000000000010011;
        weights1[19365] <= 16'b0000000000000011;
        weights1[19366] <= 16'b0000000000001100;
        weights1[19367] <= 16'b0000000000000110;
        weights1[19368] <= 16'b1111111111111010;
        weights1[19369] <= 16'b1111111111110101;
        weights1[19370] <= 16'b0000000000000001;
        weights1[19371] <= 16'b0000000000001010;
        weights1[19372] <= 16'b0000000000011001;
        weights1[19373] <= 16'b0000000000001000;
        weights1[19374] <= 16'b1111111111111111;
        weights1[19375] <= 16'b1111111111111001;
        weights1[19376] <= 16'b0000000000000000;
        weights1[19377] <= 16'b0000000000000010;
        weights1[19378] <= 16'b1111111111111000;
        weights1[19379] <= 16'b0000000000000110;
        weights1[19380] <= 16'b0000000000000011;
        weights1[19381] <= 16'b1111111111111100;
        weights1[19382] <= 16'b0000000000001111;
        weights1[19383] <= 16'b1111111111111010;
        weights1[19384] <= 16'b0000000000001101;
        weights1[19385] <= 16'b1111111111111001;
        weights1[19386] <= 16'b1111111111111101;
        weights1[19387] <= 16'b0000000000001010;
        weights1[19388] <= 16'b0000000000000011;
        weights1[19389] <= 16'b0000000000001001;
        weights1[19390] <= 16'b0000000000001011;
        weights1[19391] <= 16'b0000000000001001;
        weights1[19392] <= 16'b0000000000000011;
        weights1[19393] <= 16'b1111111111111011;
        weights1[19394] <= 16'b1111111111111111;
        weights1[19395] <= 16'b1111111111110100;
        weights1[19396] <= 16'b0000000000010110;
        weights1[19397] <= 16'b0000000000000100;
        weights1[19398] <= 16'b1111111111101010;
        weights1[19399] <= 16'b1111111111111100;
        weights1[19400] <= 16'b1111111111110110;
        weights1[19401] <= 16'b1111111111110011;
        weights1[19402] <= 16'b1111111111111011;
        weights1[19403] <= 16'b0000000000000001;
        weights1[19404] <= 16'b0000000000000000;
        weights1[19405] <= 16'b0000000000001011;
        weights1[19406] <= 16'b0000000000000110;
        weights1[19407] <= 16'b1111111111111100;
        weights1[19408] <= 16'b1111111111111111;
        weights1[19409] <= 16'b1111111111110010;
        weights1[19410] <= 16'b0000000000000000;
        weights1[19411] <= 16'b1111111111110000;
        weights1[19412] <= 16'b1111111111100011;
        weights1[19413] <= 16'b0000000000001111;
        weights1[19414] <= 16'b1111111111110100;
        weights1[19415] <= 16'b1111111111110011;
        weights1[19416] <= 16'b1111111111111110;
        weights1[19417] <= 16'b1111111111111000;
        weights1[19418] <= 16'b0000000000000011;
        weights1[19419] <= 16'b0000000000000000;
        weights1[19420] <= 16'b1111111111110110;
        weights1[19421] <= 16'b0000000000001001;
        weights1[19422] <= 16'b1111111111111111;
        weights1[19423] <= 16'b1111111111110010;
        weights1[19424] <= 16'b1111111111101111;
        weights1[19425] <= 16'b0000000000010001;
        weights1[19426] <= 16'b0000000000001000;
        weights1[19427] <= 16'b0000000000001010;
        weights1[19428] <= 16'b1111111111111011;
        weights1[19429] <= 16'b0000000000011100;
        weights1[19430] <= 16'b1111111111111000;
        weights1[19431] <= 16'b1111111111110111;
        weights1[19432] <= 16'b0000000000000100;
        weights1[19433] <= 16'b1111111111111101;
        weights1[19434] <= 16'b0000000000001110;
        weights1[19435] <= 16'b0000000000000000;
        weights1[19436] <= 16'b0000000000000110;
        weights1[19437] <= 16'b1111111111110111;
        weights1[19438] <= 16'b0000000000010000;
        weights1[19439] <= 16'b0000000000000000;
        weights1[19440] <= 16'b1111111111111111;
        weights1[19441] <= 16'b1111111111100101;
        weights1[19442] <= 16'b1111111111101001;
        weights1[19443] <= 16'b1111111111111001;
        weights1[19444] <= 16'b0000000000010010;
        weights1[19445] <= 16'b1111111111110011;
        weights1[19446] <= 16'b1111111111101111;
        weights1[19447] <= 16'b0000000000000101;
        weights1[19448] <= 16'b0000000000001100;
        weights1[19449] <= 16'b0000000000000001;
        weights1[19450] <= 16'b0000000000000100;
        weights1[19451] <= 16'b0000000000000101;
        weights1[19452] <= 16'b1111111111110011;
        weights1[19453] <= 16'b1111111111111011;
        weights1[19454] <= 16'b0000000000000101;
        weights1[19455] <= 16'b0000000000000000;
        weights1[19456] <= 16'b1111111111111000;
        weights1[19457] <= 16'b1111111111110100;
        weights1[19458] <= 16'b1111111111111010;
        weights1[19459] <= 16'b1111111111111010;
        weights1[19460] <= 16'b0000000000000101;
        weights1[19461] <= 16'b0000000000000010;
        weights1[19462] <= 16'b0000000000000110;
        weights1[19463] <= 16'b1111111111111101;
        weights1[19464] <= 16'b1111111111111110;
        weights1[19465] <= 16'b0000000000000011;
        weights1[19466] <= 16'b0000000000001010;
        weights1[19467] <= 16'b0000000000000101;
        weights1[19468] <= 16'b0000000000000011;
        weights1[19469] <= 16'b0000000000010111;
        weights1[19470] <= 16'b0000000000001000;
        weights1[19471] <= 16'b1111111111111001;
        weights1[19472] <= 16'b1111111111101000;
        weights1[19473] <= 16'b0000000000000101;
        weights1[19474] <= 16'b1111111111110001;
        weights1[19475] <= 16'b0000000000000011;
        weights1[19476] <= 16'b1111111111110001;
        weights1[19477] <= 16'b0000000000001001;
        weights1[19478] <= 16'b1111111111111000;
        weights1[19479] <= 16'b0000000000010101;
        weights1[19480] <= 16'b1111111111111111;
        weights1[19481] <= 16'b1111111111111000;
        weights1[19482] <= 16'b1111111111101011;
        weights1[19483] <= 16'b1111111111111100;
        weights1[19484] <= 16'b1111111111101111;
        weights1[19485] <= 16'b1111111111111001;
        weights1[19486] <= 16'b0000000000000001;
        weights1[19487] <= 16'b1111111111110101;
        weights1[19488] <= 16'b0000000000001000;
        weights1[19489] <= 16'b0000000000001001;
        weights1[19490] <= 16'b0000000000000100;
        weights1[19491] <= 16'b1111111111111001;
        weights1[19492] <= 16'b1111111111111000;
        weights1[19493] <= 16'b0000000000000000;
        weights1[19494] <= 16'b0000000000000001;
        weights1[19495] <= 16'b0000000000000000;
        weights1[19496] <= 16'b1111111111111001;
        weights1[19497] <= 16'b0000000000000100;
        weights1[19498] <= 16'b0000000000000010;
        weights1[19499] <= 16'b0000000000000000;
        weights1[19500] <= 16'b1111111111111000;
        weights1[19501] <= 16'b1111111111111111;
        weights1[19502] <= 16'b1111111111101011;
        weights1[19503] <= 16'b1111111111101001;
        weights1[19504] <= 16'b1111111111111000;
        weights1[19505] <= 16'b1111111111101101;
        weights1[19506] <= 16'b0000000000001101;
        weights1[19507] <= 16'b0000000000000110;
        weights1[19508] <= 16'b1111111111111000;
        weights1[19509] <= 16'b0000000000000100;
        weights1[19510] <= 16'b0000000000000100;
        weights1[19511] <= 16'b0000000000001011;
        weights1[19512] <= 16'b1111111111110100;
        weights1[19513] <= 16'b1111111111111110;
        weights1[19514] <= 16'b0000000000000000;
        weights1[19515] <= 16'b1111111111111100;
        weights1[19516] <= 16'b0000000000001001;
        weights1[19517] <= 16'b0000000000000010;
        weights1[19518] <= 16'b0000000000000100;
        weights1[19519] <= 16'b1111111111111111;
        weights1[19520] <= 16'b1111111111110101;
        weights1[19521] <= 16'b1111111111111101;
        weights1[19522] <= 16'b1111111111110110;
        weights1[19523] <= 16'b1111111111111001;
        weights1[19524] <= 16'b1111111111110010;
        weights1[19525] <= 16'b0000000000000000;
        weights1[19526] <= 16'b0000000000000011;
        weights1[19527] <= 16'b0000000000001000;
        weights1[19528] <= 16'b1111111111110110;
        weights1[19529] <= 16'b1111111111101110;
        weights1[19530] <= 16'b1111111111110000;
        weights1[19531] <= 16'b0000000000000000;
        weights1[19532] <= 16'b1111111111110101;
        weights1[19533] <= 16'b1111111111110001;
        weights1[19534] <= 16'b1111111111111101;
        weights1[19535] <= 16'b1111111111111001;
        weights1[19536] <= 16'b0000000000000010;
        weights1[19537] <= 16'b1111111111101000;
        weights1[19538] <= 16'b0000000000000001;
        weights1[19539] <= 16'b0000000000000110;
        weights1[19540] <= 16'b1111111111111110;
        weights1[19541] <= 16'b1111111111110101;
        weights1[19542] <= 16'b1111111111111000;
        weights1[19543] <= 16'b1111111111111100;
        weights1[19544] <= 16'b0000000000000000;
        weights1[19545] <= 16'b0000000000000010;
        weights1[19546] <= 16'b0000000000000001;
        weights1[19547] <= 16'b1111111111110011;
        weights1[19548] <= 16'b1111111111111101;
        weights1[19549] <= 16'b1111111111110101;
        weights1[19550] <= 16'b1111111111110111;
        weights1[19551] <= 16'b1111111111111110;
        weights1[19552] <= 16'b1111111111111000;
        weights1[19553] <= 16'b0000000000000001;
        weights1[19554] <= 16'b1111111111110011;
        weights1[19555] <= 16'b1111111111111010;
        weights1[19556] <= 16'b1111111111111110;
        weights1[19557] <= 16'b1111111111111000;
        weights1[19558] <= 16'b0000000000000110;
        weights1[19559] <= 16'b1111111111110111;
        weights1[19560] <= 16'b0000000000000000;
        weights1[19561] <= 16'b1111111111110111;
        weights1[19562] <= 16'b1111111111111010;
        weights1[19563] <= 16'b1111111111110111;
        weights1[19564] <= 16'b0000000000000001;
        weights1[19565] <= 16'b0000000000001110;
        weights1[19566] <= 16'b0000000000001001;
        weights1[19567] <= 16'b0000000000001100;
        weights1[19568] <= 16'b1111111111110011;
        weights1[19569] <= 16'b1111111111110110;
        weights1[19570] <= 16'b1111111111110110;
        weights1[19571] <= 16'b0000000000000011;
        weights1[19572] <= 16'b1111111111111101;
        weights1[19573] <= 16'b1111111111111111;
        weights1[19574] <= 16'b1111111111111110;
        weights1[19575] <= 16'b1111111111111010;
        weights1[19576] <= 16'b1111111111101110;
        weights1[19577] <= 16'b1111111111111110;
        weights1[19578] <= 16'b1111111111111101;
        weights1[19579] <= 16'b1111111111101110;
        weights1[19580] <= 16'b1111111111111011;
        weights1[19581] <= 16'b1111111111111000;
        weights1[19582] <= 16'b1111111111110011;
        weights1[19583] <= 16'b1111111111110011;
        weights1[19584] <= 16'b0000000000000100;
        weights1[19585] <= 16'b1111111111111010;
        weights1[19586] <= 16'b1111111111111100;
        weights1[19587] <= 16'b1111111111111111;
        weights1[19588] <= 16'b1111111111111111;
        weights1[19589] <= 16'b1111111111111110;
        weights1[19590] <= 16'b1111111111111000;
        weights1[19591] <= 16'b1111111111101101;
        weights1[19592] <= 16'b1111111111101011;
        weights1[19593] <= 16'b1111111111110101;
        weights1[19594] <= 16'b1111111111110011;
        weights1[19595] <= 16'b1111111111111010;
        weights1[19596] <= 16'b1111111111110111;
        weights1[19597] <= 16'b1111111111111000;
        weights1[19598] <= 16'b1111111111111001;
        weights1[19599] <= 16'b0000000000000100;
        weights1[19600] <= 16'b0000000000000000;
        weights1[19601] <= 16'b0000000000000000;
        weights1[19602] <= 16'b1111111111111110;
        weights1[19603] <= 16'b1111111111111110;
        weights1[19604] <= 16'b1111111111111110;
        weights1[19605] <= 16'b1111111111110111;
        weights1[19606] <= 16'b1111111111110000;
        weights1[19607] <= 16'b1111111111100110;
        weights1[19608] <= 16'b1111111111100100;
        weights1[19609] <= 16'b1111111111011011;
        weights1[19610] <= 16'b1111111111001110;
        weights1[19611] <= 16'b1111111111010100;
        weights1[19612] <= 16'b1111111111011000;
        weights1[19613] <= 16'b1111111111100111;
        weights1[19614] <= 16'b1111111111100100;
        weights1[19615] <= 16'b1111111111111100;
        weights1[19616] <= 16'b0000000000001110;
        weights1[19617] <= 16'b0000000000000111;
        weights1[19618] <= 16'b0000000000011011;
        weights1[19619] <= 16'b0000000000010000;
        weights1[19620] <= 16'b0000000000011001;
        weights1[19621] <= 16'b0000000000010010;
        weights1[19622] <= 16'b0000000000011111;
        weights1[19623] <= 16'b0000000000011111;
        weights1[19624] <= 16'b0000000000011001;
        weights1[19625] <= 16'b0000000000010010;
        weights1[19626] <= 16'b0000000000001010;
        weights1[19627] <= 16'b0000000000000101;
        weights1[19628] <= 16'b0000000000000000;
        weights1[19629] <= 16'b1111111111111110;
        weights1[19630] <= 16'b1111111111111100;
        weights1[19631] <= 16'b1111111111111100;
        weights1[19632] <= 16'b1111111111110101;
        weights1[19633] <= 16'b1111111111110110;
        weights1[19634] <= 16'b1111111111101001;
        weights1[19635] <= 16'b1111111111011111;
        weights1[19636] <= 16'b1111111111010110;
        weights1[19637] <= 16'b1111111111001110;
        weights1[19638] <= 16'b1111111111010001;
        weights1[19639] <= 16'b1111111111101010;
        weights1[19640] <= 16'b1111111111100110;
        weights1[19641] <= 16'b1111111111110111;
        weights1[19642] <= 16'b1111111111111110;
        weights1[19643] <= 16'b0000000000000100;
        weights1[19644] <= 16'b0000000000010110;
        weights1[19645] <= 16'b0000000000010011;
        weights1[19646] <= 16'b0000000000010101;
        weights1[19647] <= 16'b0000000000010110;
        weights1[19648] <= 16'b0000000000010101;
        weights1[19649] <= 16'b0000000000100000;
        weights1[19650] <= 16'b0000000000011110;
        weights1[19651] <= 16'b0000000000011100;
        weights1[19652] <= 16'b0000000000011101;
        weights1[19653] <= 16'b0000000000010101;
        weights1[19654] <= 16'b0000000000001001;
        weights1[19655] <= 16'b0000000000000011;
        weights1[19656] <= 16'b0000000000000000;
        weights1[19657] <= 16'b1111111111111100;
        weights1[19658] <= 16'b1111111111111001;
        weights1[19659] <= 16'b1111111111110111;
        weights1[19660] <= 16'b1111111111101111;
        weights1[19661] <= 16'b1111111111110000;
        weights1[19662] <= 16'b1111111111100010;
        weights1[19663] <= 16'b1111111111011101;
        weights1[19664] <= 16'b1111111111011001;
        weights1[19665] <= 16'b1111111111001110;
        weights1[19666] <= 16'b1111111111100111;
        weights1[19667] <= 16'b1111111111101111;
        weights1[19668] <= 16'b0000000000000010;
        weights1[19669] <= 16'b1111111111110101;
        weights1[19670] <= 16'b0000000000000110;
        weights1[19671] <= 16'b0000000000010111;
        weights1[19672] <= 16'b1111111111111101;
        weights1[19673] <= 16'b0000000000011011;
        weights1[19674] <= 16'b0000000000001110;
        weights1[19675] <= 16'b0000000000011001;
        weights1[19676] <= 16'b0000000000101010;
        weights1[19677] <= 16'b0000000000100001;
        weights1[19678] <= 16'b0000000000100100;
        weights1[19679] <= 16'b0000000000100111;
        weights1[19680] <= 16'b0000000000011011;
        weights1[19681] <= 16'b0000000000010010;
        weights1[19682] <= 16'b0000000000010001;
        weights1[19683] <= 16'b0000000000000110;
        weights1[19684] <= 16'b1111111111111110;
        weights1[19685] <= 16'b1111111111111010;
        weights1[19686] <= 16'b1111111111110100;
        weights1[19687] <= 16'b1111111111101110;
        weights1[19688] <= 16'b1111111111101000;
        weights1[19689] <= 16'b1111111111110000;
        weights1[19690] <= 16'b1111111111100100;
        weights1[19691] <= 16'b1111111111010101;
        weights1[19692] <= 16'b1111111111110010;
        weights1[19693] <= 16'b1111111111101000;
        weights1[19694] <= 16'b0000000000000111;
        weights1[19695] <= 16'b0000000000010000;
        weights1[19696] <= 16'b1111111111111110;
        weights1[19697] <= 16'b0000000000001000;
        weights1[19698] <= 16'b1111111111111100;
        weights1[19699] <= 16'b0000000000001011;
        weights1[19700] <= 16'b0000000000001010;
        weights1[19701] <= 16'b0000000000010011;
        weights1[19702] <= 16'b0000000000011010;
        weights1[19703] <= 16'b0000000000001001;
        weights1[19704] <= 16'b0000000000010011;
        weights1[19705] <= 16'b0000000000011010;
        weights1[19706] <= 16'b0000000000011011;
        weights1[19707] <= 16'b0000000000010001;
        weights1[19708] <= 16'b0000000000001111;
        weights1[19709] <= 16'b0000000000001011;
        weights1[19710] <= 16'b0000000000010100;
        weights1[19711] <= 16'b0000000000001001;
        weights1[19712] <= 16'b1111111111111011;
        weights1[19713] <= 16'b1111111111110100;
        weights1[19714] <= 16'b1111111111101101;
        weights1[19715] <= 16'b1111111111100100;
        weights1[19716] <= 16'b1111111111100101;
        weights1[19717] <= 16'b1111111111110001;
        weights1[19718] <= 16'b1111111111100100;
        weights1[19719] <= 16'b1111111111110011;
        weights1[19720] <= 16'b1111111111110101;
        weights1[19721] <= 16'b0000000000010011;
        weights1[19722] <= 16'b0000000000011111;
        weights1[19723] <= 16'b0000000000101001;
        weights1[19724] <= 16'b1111111111111111;
        weights1[19725] <= 16'b0000000000011111;
        weights1[19726] <= 16'b0000000000100100;
        weights1[19727] <= 16'b0000000000011000;
        weights1[19728] <= 16'b0000000000011001;
        weights1[19729] <= 16'b0000000000010101;
        weights1[19730] <= 16'b0000000000100000;
        weights1[19731] <= 16'b0000000000001100;
        weights1[19732] <= 16'b0000000000001000;
        weights1[19733] <= 16'b0000000000011010;
        weights1[19734] <= 16'b0000000000001011;
        weights1[19735] <= 16'b0000000000011011;
        weights1[19736] <= 16'b0000000000011100;
        weights1[19737] <= 16'b0000000000011000;
        weights1[19738] <= 16'b0000000000100111;
        weights1[19739] <= 16'b0000000000010101;
        weights1[19740] <= 16'b1111111111111010;
        weights1[19741] <= 16'b1111111111101111;
        weights1[19742] <= 16'b1111111111100111;
        weights1[19743] <= 16'b1111111111011110;
        weights1[19744] <= 16'b1111111111100110;
        weights1[19745] <= 16'b1111111111101001;
        weights1[19746] <= 16'b1111111111111111;
        weights1[19747] <= 16'b1111111111111100;
        weights1[19748] <= 16'b0000000000100101;
        weights1[19749] <= 16'b0000000000101000;
        weights1[19750] <= 16'b0000000000110100;
        weights1[19751] <= 16'b0000000000011101;
        weights1[19752] <= 16'b0000000000111101;
        weights1[19753] <= 16'b0000000000100001;
        weights1[19754] <= 16'b0000000000010001;
        weights1[19755] <= 16'b0000000000101000;
        weights1[19756] <= 16'b0000000000010001;
        weights1[19757] <= 16'b0000000000010111;
        weights1[19758] <= 16'b0000000000011010;
        weights1[19759] <= 16'b0000000000011101;
        weights1[19760] <= 16'b0000000000100110;
        weights1[19761] <= 16'b0000000000100010;
        weights1[19762] <= 16'b0000000000011110;
        weights1[19763] <= 16'b0000000000101011;
        weights1[19764] <= 16'b0000000000111100;
        weights1[19765] <= 16'b0000000000110000;
        weights1[19766] <= 16'b0000000000100100;
        weights1[19767] <= 16'b0000000000100010;
        weights1[19768] <= 16'b1111111111110111;
        weights1[19769] <= 16'b1111111111101110;
        weights1[19770] <= 16'b1111111111100010;
        weights1[19771] <= 16'b1111111111101001;
        weights1[19772] <= 16'b1111111111101101;
        weights1[19773] <= 16'b1111111111111110;
        weights1[19774] <= 16'b1111111111110101;
        weights1[19775] <= 16'b0000000000001101;
        weights1[19776] <= 16'b0000000000011110;
        weights1[19777] <= 16'b0000000001000010;
        weights1[19778] <= 16'b0000000001000101;
        weights1[19779] <= 16'b0000000001000001;
        weights1[19780] <= 16'b0000000000111100;
        weights1[19781] <= 16'b0000000000011111;
        weights1[19782] <= 16'b0000000000010101;
        weights1[19783] <= 16'b0000000000100001;
        weights1[19784] <= 16'b0000000001000000;
        weights1[19785] <= 16'b0000000000010000;
        weights1[19786] <= 16'b0000000000011110;
        weights1[19787] <= 16'b0000000000100100;
        weights1[19788] <= 16'b0000000000010011;
        weights1[19789] <= 16'b0000000000100100;
        weights1[19790] <= 16'b0000000000101111;
        weights1[19791] <= 16'b0000000000100110;
        weights1[19792] <= 16'b0000000000100101;
        weights1[19793] <= 16'b0000000000101000;
        weights1[19794] <= 16'b0000000000101100;
        weights1[19795] <= 16'b0000000000100101;
        weights1[19796] <= 16'b1111111111110100;
        weights1[19797] <= 16'b1111111111101100;
        weights1[19798] <= 16'b1111111111101010;
        weights1[19799] <= 16'b1111111111110110;
        weights1[19800] <= 16'b1111111111110101;
        weights1[19801] <= 16'b0000000000000101;
        weights1[19802] <= 16'b0000000000001000;
        weights1[19803] <= 16'b0000000000011110;
        weights1[19804] <= 16'b0000000000100101;
        weights1[19805] <= 16'b0000000000100010;
        weights1[19806] <= 16'b0000000000111010;
        weights1[19807] <= 16'b0000000001000011;
        weights1[19808] <= 16'b0000000001000110;
        weights1[19809] <= 16'b0000000000100010;
        weights1[19810] <= 16'b0000000000101011;
        weights1[19811] <= 16'b0000000000011111;
        weights1[19812] <= 16'b0000000000010101;
        weights1[19813] <= 16'b0000000000011110;
        weights1[19814] <= 16'b0000000000011111;
        weights1[19815] <= 16'b0000000000011110;
        weights1[19816] <= 16'b0000000000101000;
        weights1[19817] <= 16'b0000000000000001;
        weights1[19818] <= 16'b0000000000000111;
        weights1[19819] <= 16'b1111111111111101;
        weights1[19820] <= 16'b0000000000100010;
        weights1[19821] <= 16'b0000000000011100;
        weights1[19822] <= 16'b0000000000100110;
        weights1[19823] <= 16'b0000000000101011;
        weights1[19824] <= 16'b1111111111101100;
        weights1[19825] <= 16'b1111111111101010;
        weights1[19826] <= 16'b1111111111110100;
        weights1[19827] <= 16'b1111111111101000;
        weights1[19828] <= 16'b1111111111011011;
        weights1[19829] <= 16'b0000000000011010;
        weights1[19830] <= 16'b0000000000001001;
        weights1[19831] <= 16'b0000000000100011;
        weights1[19832] <= 16'b0000000000100011;
        weights1[19833] <= 16'b0000000000101101;
        weights1[19834] <= 16'b0000000001000001;
        weights1[19835] <= 16'b0000000001001000;
        weights1[19836] <= 16'b0000000000111100;
        weights1[19837] <= 16'b0000000000011100;
        weights1[19838] <= 16'b0000000001000010;
        weights1[19839] <= 16'b0000000001001000;
        weights1[19840] <= 16'b0000000000100000;
        weights1[19841] <= 16'b0000000000011011;
        weights1[19842] <= 16'b0000000000010011;
        weights1[19843] <= 16'b1111111111111001;
        weights1[19844] <= 16'b0000000000001001;
        weights1[19845] <= 16'b1111111111010101;
        weights1[19846] <= 16'b0000000000000111;
        weights1[19847] <= 16'b0000000000000000;
        weights1[19848] <= 16'b0000000000010001;
        weights1[19849] <= 16'b0000000000001011;
        weights1[19850] <= 16'b0000000000010101;
        weights1[19851] <= 16'b0000000000100010;
        weights1[19852] <= 16'b1111111111101101;
        weights1[19853] <= 16'b1111111111110001;
        weights1[19854] <= 16'b1111111111111101;
        weights1[19855] <= 16'b0000000000000101;
        weights1[19856] <= 16'b1111111111110110;
        weights1[19857] <= 16'b0000000000001010;
        weights1[19858] <= 16'b0000000000001101;
        weights1[19859] <= 16'b0000000000010001;
        weights1[19860] <= 16'b0000000000110010;
        weights1[19861] <= 16'b0000000000110001;
        weights1[19862] <= 16'b0000000001010011;
        weights1[19863] <= 16'b0000000000101110;
        weights1[19864] <= 16'b0000000000000101;
        weights1[19865] <= 16'b1111111111100010;
        weights1[19866] <= 16'b1111111111100100;
        weights1[19867] <= 16'b0000000000011110;
        weights1[19868] <= 16'b0000000000011010;
        weights1[19869] <= 16'b1111111111101110;
        weights1[19870] <= 16'b1111111111101101;
        weights1[19871] <= 16'b1111111111110100;
        weights1[19872] <= 16'b1111111111111011;
        weights1[19873] <= 16'b1111111111111010;
        weights1[19874] <= 16'b1111111111110011;
        weights1[19875] <= 16'b1111111111110011;
        weights1[19876] <= 16'b0000000000001010;
        weights1[19877] <= 16'b0000000000010010;
        weights1[19878] <= 16'b0000000000001111;
        weights1[19879] <= 16'b0000000000010100;
        weights1[19880] <= 16'b1111111111110000;
        weights1[19881] <= 16'b1111111111110101;
        weights1[19882] <= 16'b0000000000000101;
        weights1[19883] <= 16'b0000000000001011;
        weights1[19884] <= 16'b0000000000001010;
        weights1[19885] <= 16'b0000000000001010;
        weights1[19886] <= 16'b0000000000001100;
        weights1[19887] <= 16'b0000000000000010;
        weights1[19888] <= 16'b0000000000010011;
        weights1[19889] <= 16'b0000000000100010;
        weights1[19890] <= 16'b0000000001000101;
        weights1[19891] <= 16'b0000000000110011;
        weights1[19892] <= 16'b1111111111100000;
        weights1[19893] <= 16'b1111111110000010;
        weights1[19894] <= 16'b1111111110000010;
        weights1[19895] <= 16'b1111111111011000;
        weights1[19896] <= 16'b1111111111101000;
        weights1[19897] <= 16'b1111111111110101;
        weights1[19898] <= 16'b1111111111100100;
        weights1[19899] <= 16'b1111111111100110;
        weights1[19900] <= 16'b1111111111110000;
        weights1[19901] <= 16'b1111111111111011;
        weights1[19902] <= 16'b1111111111011111;
        weights1[19903] <= 16'b0000000000000000;
        weights1[19904] <= 16'b1111111111111111;
        weights1[19905] <= 16'b0000000000001100;
        weights1[19906] <= 16'b0000000000001101;
        weights1[19907] <= 16'b0000000000010100;
        weights1[19908] <= 16'b1111111111111001;
        weights1[19909] <= 16'b0000000000000110;
        weights1[19910] <= 16'b0000000000010110;
        weights1[19911] <= 16'b0000000000010111;
        weights1[19912] <= 16'b0000000000011010;
        weights1[19913] <= 16'b0000000000010001;
        weights1[19914] <= 16'b0000000000011000;
        weights1[19915] <= 16'b0000000000010111;
        weights1[19916] <= 16'b0000000000010101;
        weights1[19917] <= 16'b0000000000001101;
        weights1[19918] <= 16'b0000000000101100;
        weights1[19919] <= 16'b0000000000000100;
        weights1[19920] <= 16'b1111111110111000;
        weights1[19921] <= 16'b1111111101110101;
        weights1[19922] <= 16'b1111111101110110;
        weights1[19923] <= 16'b1111111111000001;
        weights1[19924] <= 16'b0000000000000000;
        weights1[19925] <= 16'b1111111111011001;
        weights1[19926] <= 16'b1111111111100100;
        weights1[19927] <= 16'b1111111111010010;
        weights1[19928] <= 16'b1111111111100110;
        weights1[19929] <= 16'b1111111111100011;
        weights1[19930] <= 16'b1111111111100011;
        weights1[19931] <= 16'b1111111111101111;
        weights1[19932] <= 16'b1111111111111010;
        weights1[19933] <= 16'b1111111111111110;
        weights1[19934] <= 16'b0000000000011000;
        weights1[19935] <= 16'b0000000000010100;
        weights1[19936] <= 16'b1111111111111011;
        weights1[19937] <= 16'b0000000000010101;
        weights1[19938] <= 16'b0000000000011011;
        weights1[19939] <= 16'b0000000000100001;
        weights1[19940] <= 16'b0000000000100101;
        weights1[19941] <= 16'b0000000000010011;
        weights1[19942] <= 16'b0000000000000110;
        weights1[19943] <= 16'b0000000000011100;
        weights1[19944] <= 16'b0000000000010001;
        weights1[19945] <= 16'b0000000000001100;
        weights1[19946] <= 16'b0000000000011001;
        weights1[19947] <= 16'b0000000000011100;
        weights1[19948] <= 16'b1111111111010100;
        weights1[19949] <= 16'b1111111110101000;
        weights1[19950] <= 16'b1111111110011111;
        weights1[19951] <= 16'b1111111111100010;
        weights1[19952] <= 16'b1111111111110010;
        weights1[19953] <= 16'b1111111111110001;
        weights1[19954] <= 16'b1111111111110101;
        weights1[19955] <= 16'b1111111111010111;
        weights1[19956] <= 16'b1111111111110111;
        weights1[19957] <= 16'b1111111111011101;
        weights1[19958] <= 16'b1111111111101100;
        weights1[19959] <= 16'b1111111111110011;
        weights1[19960] <= 16'b1111111111110010;
        weights1[19961] <= 16'b0000000000000001;
        weights1[19962] <= 16'b0000000000001001;
        weights1[19963] <= 16'b0000000000010101;
        weights1[19964] <= 16'b1111111111111000;
        weights1[19965] <= 16'b0000000000001001;
        weights1[19966] <= 16'b0000000000010110;
        weights1[19967] <= 16'b0000000000100010;
        weights1[19968] <= 16'b0000000000110000;
        weights1[19969] <= 16'b0000000000001101;
        weights1[19970] <= 16'b0000000000001110;
        weights1[19971] <= 16'b0000000000101111;
        weights1[19972] <= 16'b1111111111110001;
        weights1[19973] <= 16'b0000000000011100;
        weights1[19974] <= 16'b0000000000010010;
        weights1[19975] <= 16'b0000000000000110;
        weights1[19976] <= 16'b1111111111000110;
        weights1[19977] <= 16'b1111111110110011;
        weights1[19978] <= 16'b1111111110011010;
        weights1[19979] <= 16'b1111111110111101;
        weights1[19980] <= 16'b1111111111100011;
        weights1[19981] <= 16'b1111111111111010;
        weights1[19982] <= 16'b1111111111111111;
        weights1[19983] <= 16'b1111111111011011;
        weights1[19984] <= 16'b1111111111111110;
        weights1[19985] <= 16'b1111111111101110;
        weights1[19986] <= 16'b1111111111110100;
        weights1[19987] <= 16'b1111111111111111;
        weights1[19988] <= 16'b1111111111110100;
        weights1[19989] <= 16'b1111111111110111;
        weights1[19990] <= 16'b0000000000010010;
        weights1[19991] <= 16'b0000000000011000;
        weights1[19992] <= 16'b0000000000000100;
        weights1[19993] <= 16'b0000000000001110;
        weights1[19994] <= 16'b0000000000011010;
        weights1[19995] <= 16'b0000000000010011;
        weights1[19996] <= 16'b0000000000100010;
        weights1[19997] <= 16'b0000000000001000;
        weights1[19998] <= 16'b1111111111111101;
        weights1[19999] <= 16'b0000000000000110;
        weights1[20000] <= 16'b0000000000001010;
        weights1[20001] <= 16'b0000000000011010;
        weights1[20002] <= 16'b0000000000000011;
        weights1[20003] <= 16'b1111111111011111;
        weights1[20004] <= 16'b1111111111011101;
        weights1[20005] <= 16'b1111111110110000;
        weights1[20006] <= 16'b1111111110111111;
        weights1[20007] <= 16'b1111111111001011;
        weights1[20008] <= 16'b1111111111110100;
        weights1[20009] <= 16'b1111111111011010;
        weights1[20010] <= 16'b1111111111101011;
        weights1[20011] <= 16'b1111111111110100;
        weights1[20012] <= 16'b1111111111111001;
        weights1[20013] <= 16'b0000000000000111;
        weights1[20014] <= 16'b1111111111111011;
        weights1[20015] <= 16'b1111111111110010;
        weights1[20016] <= 16'b1111111111110101;
        weights1[20017] <= 16'b1111111111111101;
        weights1[20018] <= 16'b0000000000011100;
        weights1[20019] <= 16'b0000000000011011;
        weights1[20020] <= 16'b1111111111111101;
        weights1[20021] <= 16'b0000000000000010;
        weights1[20022] <= 16'b0000000000001111;
        weights1[20023] <= 16'b0000000000011101;
        weights1[20024] <= 16'b1111111111111001;
        weights1[20025] <= 16'b0000000000000111;
        weights1[20026] <= 16'b1111111111111001;
        weights1[20027] <= 16'b0000000000000010;
        weights1[20028] <= 16'b0000000000010100;
        weights1[20029] <= 16'b1111111111110001;
        weights1[20030] <= 16'b0000000000001000;
        weights1[20031] <= 16'b1111111111101011;
        weights1[20032] <= 16'b1111111111001111;
        weights1[20033] <= 16'b1111111111000000;
        weights1[20034] <= 16'b1111111110110100;
        weights1[20035] <= 16'b1111111111010001;
        weights1[20036] <= 16'b1111111111011101;
        weights1[20037] <= 16'b1111111111101000;
        weights1[20038] <= 16'b1111111111111000;
        weights1[20039] <= 16'b0000000000000000;
        weights1[20040] <= 16'b0000000000000001;
        weights1[20041] <= 16'b0000000000000110;
        weights1[20042] <= 16'b1111111111110001;
        weights1[20043] <= 16'b1111111111110001;
        weights1[20044] <= 16'b1111111111100011;
        weights1[20045] <= 16'b1111111111110111;
        weights1[20046] <= 16'b0000000000001110;
        weights1[20047] <= 16'b0000000000001101;
        weights1[20048] <= 16'b1111111111111111;
        weights1[20049] <= 16'b0000000000001001;
        weights1[20050] <= 16'b0000000000000101;
        weights1[20051] <= 16'b0000000000001011;
        weights1[20052] <= 16'b1111111111011110;
        weights1[20053] <= 16'b0000000000000100;
        weights1[20054] <= 16'b1111111111110100;
        weights1[20055] <= 16'b1111111111110011;
        weights1[20056] <= 16'b1111111111111010;
        weights1[20057] <= 16'b1111111111101001;
        weights1[20058] <= 16'b1111111111110101;
        weights1[20059] <= 16'b1111111111100001;
        weights1[20060] <= 16'b1111111111100000;
        weights1[20061] <= 16'b1111111110110000;
        weights1[20062] <= 16'b1111111111000010;
        weights1[20063] <= 16'b1111111111101101;
        weights1[20064] <= 16'b1111111111011010;
        weights1[20065] <= 16'b1111111111100100;
        weights1[20066] <= 16'b1111111111101001;
        weights1[20067] <= 16'b1111111111101110;
        weights1[20068] <= 16'b1111111111111101;
        weights1[20069] <= 16'b0000000000001000;
        weights1[20070] <= 16'b0000000000000000;
        weights1[20071] <= 16'b1111111111100111;
        weights1[20072] <= 16'b1111111111101010;
        weights1[20073] <= 16'b1111111111110010;
        weights1[20074] <= 16'b1111111111111111;
        weights1[20075] <= 16'b0000000000000000;
        weights1[20076] <= 16'b0000000000000111;
        weights1[20077] <= 16'b0000000000000101;
        weights1[20078] <= 16'b0000000000000000;
        weights1[20079] <= 16'b0000000000001001;
        weights1[20080] <= 16'b1111111111110110;
        weights1[20081] <= 16'b0000000000001010;
        weights1[20082] <= 16'b1111111111101101;
        weights1[20083] <= 16'b1111111111101011;
        weights1[20084] <= 16'b1111111111110011;
        weights1[20085] <= 16'b1111111111100101;
        weights1[20086] <= 16'b1111111111101111;
        weights1[20087] <= 16'b1111111111101011;
        weights1[20088] <= 16'b1111111111010111;
        weights1[20089] <= 16'b1111111111000110;
        weights1[20090] <= 16'b1111111110111110;
        weights1[20091] <= 16'b1111111111010000;
        weights1[20092] <= 16'b0000000000000100;
        weights1[20093] <= 16'b1111111111101011;
        weights1[20094] <= 16'b0000000000001010;
        weights1[20095] <= 16'b1111111111110011;
        weights1[20096] <= 16'b0000000000001000;
        weights1[20097] <= 16'b1111111111110110;
        weights1[20098] <= 16'b1111111111011001;
        weights1[20099] <= 16'b1111111111100110;
        weights1[20100] <= 16'b1111111111100101;
        weights1[20101] <= 16'b1111111111101100;
        weights1[20102] <= 16'b1111111111111010;
        weights1[20103] <= 16'b1111111111111010;
        weights1[20104] <= 16'b0000000000000111;
        weights1[20105] <= 16'b0000000000000011;
        weights1[20106] <= 16'b1111111111111111;
        weights1[20107] <= 16'b0000000000000110;
        weights1[20108] <= 16'b1111111111110001;
        weights1[20109] <= 16'b0000000000000010;
        weights1[20110] <= 16'b1111111111111001;
        weights1[20111] <= 16'b1111111111111001;
        weights1[20112] <= 16'b1111111111111000;
        weights1[20113] <= 16'b1111111111111001;
        weights1[20114] <= 16'b1111111111111110;
        weights1[20115] <= 16'b1111111111101101;
        weights1[20116] <= 16'b1111111111100010;
        weights1[20117] <= 16'b1111111111011001;
        weights1[20118] <= 16'b1111111111011100;
        weights1[20119] <= 16'b1111111111101111;
        weights1[20120] <= 16'b1111111111001000;
        weights1[20121] <= 16'b1111111111111000;
        weights1[20122] <= 16'b0000000000000001;
        weights1[20123] <= 16'b0000000000000001;
        weights1[20124] <= 16'b1111111111111010;
        weights1[20125] <= 16'b1111111111111101;
        weights1[20126] <= 16'b0000000000000001;
        weights1[20127] <= 16'b1111111111101001;
        weights1[20128] <= 16'b1111111111101101;
        weights1[20129] <= 16'b1111111111110011;
        weights1[20130] <= 16'b1111111111110000;
        weights1[20131] <= 16'b1111111111110100;
        weights1[20132] <= 16'b0000000000000101;
        weights1[20133] <= 16'b0000000000000000;
        weights1[20134] <= 16'b1111111111110110;
        weights1[20135] <= 16'b0000000000000100;
        weights1[20136] <= 16'b1111111111101110;
        weights1[20137] <= 16'b1111111111110010;
        weights1[20138] <= 16'b1111111111101001;
        weights1[20139] <= 16'b1111111111100111;
        weights1[20140] <= 16'b1111111111111000;
        weights1[20141] <= 16'b1111111111111110;
        weights1[20142] <= 16'b1111111111101100;
        weights1[20143] <= 16'b1111111111110000;
        weights1[20144] <= 16'b1111111111100011;
        weights1[20145] <= 16'b1111111111001000;
        weights1[20146] <= 16'b1111111111111010;
        weights1[20147] <= 16'b1111111111111110;
        weights1[20148] <= 16'b1111111111100010;
        weights1[20149] <= 16'b0000000000001101;
        weights1[20150] <= 16'b0000000000000101;
        weights1[20151] <= 16'b1111111111101111;
        weights1[20152] <= 16'b0000000000001111;
        weights1[20153] <= 16'b1111111111111100;
        weights1[20154] <= 16'b1111111111111110;
        weights1[20155] <= 16'b1111111111101110;
        weights1[20156] <= 16'b1111111111111111;
        weights1[20157] <= 16'b1111111111110000;
        weights1[20158] <= 16'b1111111111101001;
        weights1[20159] <= 16'b1111111111110000;
        weights1[20160] <= 16'b0000000000000001;
        weights1[20161] <= 16'b1111111111111011;
        weights1[20162] <= 16'b1111111111111001;
        weights1[20163] <= 16'b0000000000000000;
        weights1[20164] <= 16'b0000000000000010;
        weights1[20165] <= 16'b0000000000000100;
        weights1[20166] <= 16'b1111111111111110;
        weights1[20167] <= 16'b1111111111100111;
        weights1[20168] <= 16'b0000000000000100;
        weights1[20169] <= 16'b1111111111110101;
        weights1[20170] <= 16'b1111111111110101;
        weights1[20171] <= 16'b1111111111111100;
        weights1[20172] <= 16'b1111111111100010;
        weights1[20173] <= 16'b1111111111101010;
        weights1[20174] <= 16'b1111111111110011;
        weights1[20175] <= 16'b1111111111101010;
        weights1[20176] <= 16'b0000000000000001;
        weights1[20177] <= 16'b0000000000001010;
        weights1[20178] <= 16'b0000000000000000;
        weights1[20179] <= 16'b0000000000001000;
        weights1[20180] <= 16'b1111111111101001;
        weights1[20181] <= 16'b0000000000010000;
        weights1[20182] <= 16'b1111111111111001;
        weights1[20183] <= 16'b1111111111101111;
        weights1[20184] <= 16'b1111111111011100;
        weights1[20185] <= 16'b1111111111101110;
        weights1[20186] <= 16'b1111111111101100;
        weights1[20187] <= 16'b1111111111110100;
        weights1[20188] <= 16'b0000000000001000;
        weights1[20189] <= 16'b0000000000001111;
        weights1[20190] <= 16'b0000000000001110;
        weights1[20191] <= 16'b1111111111110101;
        weights1[20192] <= 16'b1111111111111001;
        weights1[20193] <= 16'b1111111111111101;
        weights1[20194] <= 16'b1111111111111101;
        weights1[20195] <= 16'b1111111111110011;
        weights1[20196] <= 16'b1111111111110100;
        weights1[20197] <= 16'b0000000000001111;
        weights1[20198] <= 16'b0000000000001100;
        weights1[20199] <= 16'b0000000000001100;
        weights1[20200] <= 16'b0000000000001100;
        weights1[20201] <= 16'b1111111111101110;
        weights1[20202] <= 16'b0000000000000001;
        weights1[20203] <= 16'b0000000000001001;
        weights1[20204] <= 16'b0000000000000110;
        weights1[20205] <= 16'b1111111111010001;
        weights1[20206] <= 16'b1111111111101000;
        weights1[20207] <= 16'b1111111111100110;
        weights1[20208] <= 16'b1111111111110111;
        weights1[20209] <= 16'b1111111111111001;
        weights1[20210] <= 16'b1111111111100101;
        weights1[20211] <= 16'b1111111111101010;
        weights1[20212] <= 16'b1111111111100110;
        weights1[20213] <= 16'b1111111111110010;
        weights1[20214] <= 16'b1111111111110101;
        weights1[20215] <= 16'b1111111111110110;
        weights1[20216] <= 16'b0000000000000111;
        weights1[20217] <= 16'b0000000000001110;
        weights1[20218] <= 16'b0000000000001001;
        weights1[20219] <= 16'b1111111111110111;
        weights1[20220] <= 16'b1111111111110111;
        weights1[20221] <= 16'b1111111111110001;
        weights1[20222] <= 16'b1111111111100001;
        weights1[20223] <= 16'b1111111111110110;
        weights1[20224] <= 16'b0000000000000111;
        weights1[20225] <= 16'b1111111111110010;
        weights1[20226] <= 16'b0000000000000001;
        weights1[20227] <= 16'b1111111111101101;
        weights1[20228] <= 16'b1111111111111110;
        weights1[20229] <= 16'b0000000000011000;
        weights1[20230] <= 16'b0000000000010101;
        weights1[20231] <= 16'b0000000000000110;
        weights1[20232] <= 16'b0000000000010110;
        weights1[20233] <= 16'b1111111111101111;
        weights1[20234] <= 16'b0000000000001110;
        weights1[20235] <= 16'b1111111111100010;
        weights1[20236] <= 16'b0000000000000101;
        weights1[20237] <= 16'b1111111111110111;
        weights1[20238] <= 16'b1111111111101011;
        weights1[20239] <= 16'b1111111111011011;
        weights1[20240] <= 16'b1111111111011011;
        weights1[20241] <= 16'b1111111111100110;
        weights1[20242] <= 16'b1111111111110011;
        weights1[20243] <= 16'b1111111111111000;
        weights1[20244] <= 16'b0000000000001000;
        weights1[20245] <= 16'b0000000000001001;
        weights1[20246] <= 16'b1111111111111111;
        weights1[20247] <= 16'b0000000000000100;
        weights1[20248] <= 16'b1111111111111111;
        weights1[20249] <= 16'b1111111111111110;
        weights1[20250] <= 16'b1111111111101010;
        weights1[20251] <= 16'b1111111111110111;
        weights1[20252] <= 16'b1111111111110011;
        weights1[20253] <= 16'b1111111111101011;
        weights1[20254] <= 16'b1111111111111101;
        weights1[20255] <= 16'b1111111111111010;
        weights1[20256] <= 16'b1111111111111011;
        weights1[20257] <= 16'b1111111111111010;
        weights1[20258] <= 16'b0000000000011111;
        weights1[20259] <= 16'b1111111111101100;
        weights1[20260] <= 16'b0000000000000111;
        weights1[20261] <= 16'b1111111111111110;
        weights1[20262] <= 16'b1111111111101110;
        weights1[20263] <= 16'b1111111111110011;
        weights1[20264] <= 16'b1111111111100111;
        weights1[20265] <= 16'b1111111111101101;
        weights1[20266] <= 16'b1111111111110110;
        weights1[20267] <= 16'b1111111111100110;
        weights1[20268] <= 16'b1111111111100011;
        weights1[20269] <= 16'b1111111111101110;
        weights1[20270] <= 16'b1111111111110110;
        weights1[20271] <= 16'b1111111111111010;
        weights1[20272] <= 16'b0000000000000111;
        weights1[20273] <= 16'b0000000000001011;
        weights1[20274] <= 16'b0000000000001011;
        weights1[20275] <= 16'b0000000000001001;
        weights1[20276] <= 16'b0000000000001101;
        weights1[20277] <= 16'b1111111111111111;
        weights1[20278] <= 16'b1111111111110110;
        weights1[20279] <= 16'b1111111111101001;
        weights1[20280] <= 16'b1111111111101110;
        weights1[20281] <= 16'b0000000000000000;
        weights1[20282] <= 16'b1111111111101101;
        weights1[20283] <= 16'b0000000000000000;
        weights1[20284] <= 16'b1111111111111011;
        weights1[20285] <= 16'b0000000000001011;
        weights1[20286] <= 16'b1111111111110011;
        weights1[20287] <= 16'b0000000000000010;
        weights1[20288] <= 16'b1111111111110010;
        weights1[20289] <= 16'b0000000000001101;
        weights1[20290] <= 16'b1111111111110110;
        weights1[20291] <= 16'b1111111111100011;
        weights1[20292] <= 16'b1111111111011111;
        weights1[20293] <= 16'b1111111111101011;
        weights1[20294] <= 16'b1111111111100100;
        weights1[20295] <= 16'b1111111111011110;
        weights1[20296] <= 16'b1111111111101101;
        weights1[20297] <= 16'b1111111111110001;
        weights1[20298] <= 16'b1111111111111100;
        weights1[20299] <= 16'b1111111111111110;
        weights1[20300] <= 16'b0000000000000011;
        weights1[20301] <= 16'b0000000000000001;
        weights1[20302] <= 16'b0000000000001101;
        weights1[20303] <= 16'b0000000000010000;
        weights1[20304] <= 16'b0000000000010100;
        weights1[20305] <= 16'b1111111111110110;
        weights1[20306] <= 16'b0000000000000111;
        weights1[20307] <= 16'b0000000000000001;
        weights1[20308] <= 16'b1111111111110011;
        weights1[20309] <= 16'b1111111111101111;
        weights1[20310] <= 16'b1111111111100111;
        weights1[20311] <= 16'b1111111111111010;
        weights1[20312] <= 16'b0000000000000011;
        weights1[20313] <= 16'b0000000000000100;
        weights1[20314] <= 16'b0000000000000000;
        weights1[20315] <= 16'b0000000000010100;
        weights1[20316] <= 16'b1111111111110001;
        weights1[20317] <= 16'b1111111111110110;
        weights1[20318] <= 16'b1111111111110111;
        weights1[20319] <= 16'b1111111111100110;
        weights1[20320] <= 16'b1111111111100000;
        weights1[20321] <= 16'b1111111111101001;
        weights1[20322] <= 16'b1111111111101010;
        weights1[20323] <= 16'b1111111111101100;
        weights1[20324] <= 16'b1111111111110100;
        weights1[20325] <= 16'b1111111111111010;
        weights1[20326] <= 16'b1111111111111100;
        weights1[20327] <= 16'b1111111111111101;
        weights1[20328] <= 16'b0000000000000010;
        weights1[20329] <= 16'b0000000000000000;
        weights1[20330] <= 16'b0000000000000000;
        weights1[20331] <= 16'b0000000000000110;
        weights1[20332] <= 16'b0000000000001101;
        weights1[20333] <= 16'b0000000000000010;
        weights1[20334] <= 16'b0000000000001110;
        weights1[20335] <= 16'b0000000000010001;
        weights1[20336] <= 16'b0000000000010011;
        weights1[20337] <= 16'b0000000000010011;
        weights1[20338] <= 16'b0000000000001110;
        weights1[20339] <= 16'b0000000000100011;
        weights1[20340] <= 16'b0000000000001111;
        weights1[20341] <= 16'b0000000000011100;
        weights1[20342] <= 16'b0000000000010010;
        weights1[20343] <= 16'b0000000000001011;
        weights1[20344] <= 16'b0000000000000110;
        weights1[20345] <= 16'b0000000000001000;
        weights1[20346] <= 16'b1111111111111011;
        weights1[20347] <= 16'b0000000000000011;
        weights1[20348] <= 16'b1111111111111010;
        weights1[20349] <= 16'b1111111111110010;
        weights1[20350] <= 16'b1111111111110000;
        weights1[20351] <= 16'b1111111111110010;
        weights1[20352] <= 16'b1111111111110110;
        weights1[20353] <= 16'b1111111111111101;
        weights1[20354] <= 16'b0000000000000000;
        weights1[20355] <= 16'b0000000000000000;
        weights1[20356] <= 16'b0000000000000001;
        weights1[20357] <= 16'b0000000000000000;
        weights1[20358] <= 16'b1111111111111100;
        weights1[20359] <= 16'b1111111111111010;
        weights1[20360] <= 16'b0000000000000000;
        weights1[20361] <= 16'b1111111111111101;
        weights1[20362] <= 16'b0000000000000010;
        weights1[20363] <= 16'b0000000000001101;
        weights1[20364] <= 16'b0000000000001100;
        weights1[20365] <= 16'b0000000000010010;
        weights1[20366] <= 16'b0000000000000011;
        weights1[20367] <= 16'b0000000000000101;
        weights1[20368] <= 16'b0000000000000000;
        weights1[20369] <= 16'b0000000000000010;
        weights1[20370] <= 16'b0000000000001000;
        weights1[20371] <= 16'b0000000000001000;
        weights1[20372] <= 16'b1111111111111100;
        weights1[20373] <= 16'b1111111111111100;
        weights1[20374] <= 16'b1111111111110011;
        weights1[20375] <= 16'b1111111111111011;
        weights1[20376] <= 16'b1111111111111000;
        weights1[20377] <= 16'b1111111111110100;
        weights1[20378] <= 16'b1111111111110011;
        weights1[20379] <= 16'b1111111111111010;
        weights1[20380] <= 16'b1111111111111111;
        weights1[20381] <= 16'b0000000000000000;
        weights1[20382] <= 16'b0000000000000000;
        weights1[20383] <= 16'b0000000000000000;
        weights1[20384] <= 16'b1111111111111111;
        weights1[20385] <= 16'b1111111111111111;
        weights1[20386] <= 16'b1111111111111110;
        weights1[20387] <= 16'b1111111111111111;
        weights1[20388] <= 16'b0000000000000001;
        weights1[20389] <= 16'b1111111111111110;
        weights1[20390] <= 16'b0000000000000001;
        weights1[20391] <= 16'b1111111111111101;
        weights1[20392] <= 16'b1111111111101110;
        weights1[20393] <= 16'b1111111111101111;
        weights1[20394] <= 16'b1111111111110011;
        weights1[20395] <= 16'b1111111111110011;
        weights1[20396] <= 16'b1111111111101010;
        weights1[20397] <= 16'b1111111111111001;
        weights1[20398] <= 16'b1111111111101011;
        weights1[20399] <= 16'b1111111111110011;
        weights1[20400] <= 16'b1111111111101011;
        weights1[20401] <= 16'b1111111111101010;
        weights1[20402] <= 16'b1111111111101011;
        weights1[20403] <= 16'b1111111111101101;
        weights1[20404] <= 16'b1111111111101100;
        weights1[20405] <= 16'b1111111111101110;
        weights1[20406] <= 16'b1111111111110011;
        weights1[20407] <= 16'b1111111111110010;
        weights1[20408] <= 16'b1111111111110001;
        weights1[20409] <= 16'b1111111111111010;
        weights1[20410] <= 16'b1111111111111100;
        weights1[20411] <= 16'b1111111111111110;
        weights1[20412] <= 16'b1111111111111110;
        weights1[20413] <= 16'b1111111111111110;
        weights1[20414] <= 16'b1111111111111110;
        weights1[20415] <= 16'b1111111111111010;
        weights1[20416] <= 16'b0000000000000001;
        weights1[20417] <= 16'b0000000000000010;
        weights1[20418] <= 16'b0000000000000111;
        weights1[20419] <= 16'b0000000000000000;
        weights1[20420] <= 16'b1111111111111101;
        weights1[20421] <= 16'b1111111111110000;
        weights1[20422] <= 16'b1111111111101111;
        weights1[20423] <= 16'b1111111111101110;
        weights1[20424] <= 16'b1111111111111111;
        weights1[20425] <= 16'b1111111111111011;
        weights1[20426] <= 16'b1111111111111111;
        weights1[20427] <= 16'b1111111111101011;
        weights1[20428] <= 16'b0000000000000010;
        weights1[20429] <= 16'b1111111111100011;
        weights1[20430] <= 16'b1111111111011101;
        weights1[20431] <= 16'b1111111111110001;
        weights1[20432] <= 16'b1111111111101011;
        weights1[20433] <= 16'b1111111111100000;
        weights1[20434] <= 16'b1111111111101010;
        weights1[20435] <= 16'b1111111111110101;
        weights1[20436] <= 16'b1111111111110010;
        weights1[20437] <= 16'b1111111111110100;
        weights1[20438] <= 16'b1111111111110011;
        weights1[20439] <= 16'b1111111111111100;
        weights1[20440] <= 16'b1111111111111101;
        weights1[20441] <= 16'b0000000000000000;
        weights1[20442] <= 16'b0000000000000001;
        weights1[20443] <= 16'b1111111111111111;
        weights1[20444] <= 16'b0000000000000010;
        weights1[20445] <= 16'b0000000000000100;
        weights1[20446] <= 16'b0000000000010001;
        weights1[20447] <= 16'b1111111111111100;
        weights1[20448] <= 16'b0000000000000011;
        weights1[20449] <= 16'b0000000000001100;
        weights1[20450] <= 16'b0000000000001110;
        weights1[20451] <= 16'b0000000000000000;
        weights1[20452] <= 16'b1111111111111010;
        weights1[20453] <= 16'b0000000000001011;
        weights1[20454] <= 16'b0000000000000101;
        weights1[20455] <= 16'b1111111111111011;
        weights1[20456] <= 16'b0000000000000011;
        weights1[20457] <= 16'b1111111111111001;
        weights1[20458] <= 16'b1111111111100000;
        weights1[20459] <= 16'b1111111111110100;
        weights1[20460] <= 16'b1111111111101110;
        weights1[20461] <= 16'b1111111111100011;
        weights1[20462] <= 16'b1111111111110101;
        weights1[20463] <= 16'b1111111111101101;
        weights1[20464] <= 16'b1111111111110100;
        weights1[20465] <= 16'b1111111111111001;
        weights1[20466] <= 16'b1111111111110001;
        weights1[20467] <= 16'b1111111111110101;
        weights1[20468] <= 16'b1111111111111110;
        weights1[20469] <= 16'b0000000000000010;
        weights1[20470] <= 16'b1111111111111111;
        weights1[20471] <= 16'b0000000000000101;
        weights1[20472] <= 16'b0000000000001011;
        weights1[20473] <= 16'b1111111111111001;
        weights1[20474] <= 16'b1111111111111100;
        weights1[20475] <= 16'b1111111111111111;
        weights1[20476] <= 16'b1111111111111001;
        weights1[20477] <= 16'b1111111111110011;
        weights1[20478] <= 16'b1111111111110100;
        weights1[20479] <= 16'b0000000000001010;
        weights1[20480] <= 16'b1111111111110000;
        weights1[20481] <= 16'b1111111111110011;
        weights1[20482] <= 16'b1111111111011111;
        weights1[20483] <= 16'b1111111111111111;
        weights1[20484] <= 16'b1111111111111100;
        weights1[20485] <= 16'b1111111111110110;
        weights1[20486] <= 16'b1111111111111111;
        weights1[20487] <= 16'b0000000000000100;
        weights1[20488] <= 16'b1111111111101010;
        weights1[20489] <= 16'b1111111111110011;
        weights1[20490] <= 16'b1111111111101001;
        weights1[20491] <= 16'b1111111111100110;
        weights1[20492] <= 16'b1111111111101011;
        weights1[20493] <= 16'b1111111111101110;
        weights1[20494] <= 16'b1111111111100111;
        weights1[20495] <= 16'b1111111111110110;
        weights1[20496] <= 16'b0000000000000000;
        weights1[20497] <= 16'b0000000000000110;
        weights1[20498] <= 16'b1111111111111100;
        weights1[20499] <= 16'b1111111111111101;
        weights1[20500] <= 16'b1111111111101110;
        weights1[20501] <= 16'b1111111111110110;
        weights1[20502] <= 16'b1111111111101101;
        weights1[20503] <= 16'b1111111111111100;
        weights1[20504] <= 16'b1111111111111100;
        weights1[20505] <= 16'b0000000000001011;
        weights1[20506] <= 16'b0000000000000110;
        weights1[20507] <= 16'b1111111111111010;
        weights1[20508] <= 16'b0000000000101100;
        weights1[20509] <= 16'b1111111111111100;
        weights1[20510] <= 16'b0000000000000010;
        weights1[20511] <= 16'b0000000000000101;
        weights1[20512] <= 16'b1111111111101110;
        weights1[20513] <= 16'b1111111111100111;
        weights1[20514] <= 16'b1111111111101111;
        weights1[20515] <= 16'b1111111111101111;
        weights1[20516] <= 16'b0000000000000001;
        weights1[20517] <= 16'b1111111111110101;
        weights1[20518] <= 16'b1111111111110100;
        weights1[20519] <= 16'b1111111111101011;
        weights1[20520] <= 16'b0000000000001001;
        weights1[20521] <= 16'b1111111111110010;
        weights1[20522] <= 16'b1111111111110001;
        weights1[20523] <= 16'b1111111111111011;
        weights1[20524] <= 16'b0000000000000010;
        weights1[20525] <= 16'b1111111111111110;
        weights1[20526] <= 16'b1111111111111101;
        weights1[20527] <= 16'b1111111111111100;
        weights1[20528] <= 16'b1111111111110111;
        weights1[20529] <= 16'b1111111111101110;
        weights1[20530] <= 16'b0000000000000010;
        weights1[20531] <= 16'b1111111111110000;
        weights1[20532] <= 16'b1111111111111011;
        weights1[20533] <= 16'b0000000000000101;
        weights1[20534] <= 16'b1111111111111010;
        weights1[20535] <= 16'b1111111111110111;
        weights1[20536] <= 16'b1111111111111001;
        weights1[20537] <= 16'b1111111111111001;
        weights1[20538] <= 16'b0000000000000011;
        weights1[20539] <= 16'b0000000000010111;
        weights1[20540] <= 16'b1111111111110110;
        weights1[20541] <= 16'b1111111111110010;
        weights1[20542] <= 16'b0000000000010000;
        weights1[20543] <= 16'b0000000000000001;
        weights1[20544] <= 16'b0000000000000011;
        weights1[20545] <= 16'b0000000000000100;
        weights1[20546] <= 16'b0000000000100101;
        weights1[20547] <= 16'b0000000000000011;
        weights1[20548] <= 16'b0000000000000010;
        weights1[20549] <= 16'b1111111111111110;
        weights1[20550] <= 16'b1111111111111101;
        weights1[20551] <= 16'b0000000000000010;
        weights1[20552] <= 16'b1111111111111111;
        weights1[20553] <= 16'b1111111111110100;
        weights1[20554] <= 16'b1111111111110111;
        weights1[20555] <= 16'b1111111111101111;
        weights1[20556] <= 16'b1111111111110111;
        weights1[20557] <= 16'b1111111111111101;
        weights1[20558] <= 16'b1111111111110110;
        weights1[20559] <= 16'b1111111111111000;
        weights1[20560] <= 16'b0000000000000001;
        weights1[20561] <= 16'b1111111111011001;
        weights1[20562] <= 16'b1111111111101001;
        weights1[20563] <= 16'b1111111111110000;
        weights1[20564] <= 16'b0000000000001011;
        weights1[20565] <= 16'b1111111111101011;
        weights1[20566] <= 16'b1111111111111001;
        weights1[20567] <= 16'b1111111111101100;
        weights1[20568] <= 16'b0000000000000001;
        weights1[20569] <= 16'b1111111111111000;
        weights1[20570] <= 16'b1111111111110110;
        weights1[20571] <= 16'b1111111111110000;
        weights1[20572] <= 16'b1111111111101110;
        weights1[20573] <= 16'b0000000000000100;
        weights1[20574] <= 16'b1111111111101100;
        weights1[20575] <= 16'b1111111111110001;
        weights1[20576] <= 16'b1111111111111101;
        weights1[20577] <= 16'b1111111111101001;
        weights1[20578] <= 16'b1111111111111001;
        weights1[20579] <= 16'b1111111111111101;
        weights1[20580] <= 16'b1111111111111010;
        weights1[20581] <= 16'b1111111111110001;
        weights1[20582] <= 16'b1111111111111001;
        weights1[20583] <= 16'b1111111111011110;
        weights1[20584] <= 16'b1111111111100110;
        weights1[20585] <= 16'b1111111111101001;
        weights1[20586] <= 16'b1111111111101011;
        weights1[20587] <= 16'b1111111111100111;
        weights1[20588] <= 16'b1111111111111000;
        weights1[20589] <= 16'b1111111111100101;
        weights1[20590] <= 16'b1111111111100010;
        weights1[20591] <= 16'b1111111111101100;
        weights1[20592] <= 16'b1111111111010101;
        weights1[20593] <= 16'b1111111111101001;
        weights1[20594] <= 16'b1111111111110101;
        weights1[20595] <= 16'b1111111111101010;
        weights1[20596] <= 16'b1111111111101001;
        weights1[20597] <= 16'b0000000000001110;
        weights1[20598] <= 16'b1111111111111000;
        weights1[20599] <= 16'b1111111111101011;
        weights1[20600] <= 16'b1111111111110111;
        weights1[20601] <= 16'b1111111111101000;
        weights1[20602] <= 16'b0000000000011001;
        weights1[20603] <= 16'b1111111111100010;
        weights1[20604] <= 16'b0000000000000000;
        weights1[20605] <= 16'b1111111111110110;
        weights1[20606] <= 16'b0000000000000010;
        weights1[20607] <= 16'b1111111111100111;
        weights1[20608] <= 16'b1111111111110101;
        weights1[20609] <= 16'b1111111111101101;
        weights1[20610] <= 16'b1111111111110000;
        weights1[20611] <= 16'b1111111111101001;
        weights1[20612] <= 16'b1111111111101000;
        weights1[20613] <= 16'b1111111111011111;
        weights1[20614] <= 16'b1111111111101100;
        weights1[20615] <= 16'b1111111111110101;
        weights1[20616] <= 16'b1111111111011000;
        weights1[20617] <= 16'b1111111111010010;
        weights1[20618] <= 16'b1111111111111100;
        weights1[20619] <= 16'b1111111111100000;
        weights1[20620] <= 16'b1111111111110100;
        weights1[20621] <= 16'b1111111111110100;
        weights1[20622] <= 16'b1111111111011100;
        weights1[20623] <= 16'b0000000000000101;
        weights1[20624] <= 16'b1111111111111101;
        weights1[20625] <= 16'b1111111111100000;
        weights1[20626] <= 16'b1111111111111001;
        weights1[20627] <= 16'b0000000000001001;
        weights1[20628] <= 16'b0000000000001110;
        weights1[20629] <= 16'b1111111111110001;
        weights1[20630] <= 16'b1111111111111100;
        weights1[20631] <= 16'b1111111111111011;
        weights1[20632] <= 16'b0000000000000010;
        weights1[20633] <= 16'b0000000000001111;
        weights1[20634] <= 16'b1111111111110100;
        weights1[20635] <= 16'b1111111111100110;
        weights1[20636] <= 16'b1111111111101110;
        weights1[20637] <= 16'b1111111111101010;
        weights1[20638] <= 16'b1111111111101000;
        weights1[20639] <= 16'b1111111111101001;
        weights1[20640] <= 16'b1111111111100000;
        weights1[20641] <= 16'b1111111111100111;
        weights1[20642] <= 16'b1111111111001101;
        weights1[20643] <= 16'b1111111111001000;
        weights1[20644] <= 16'b1111111111000100;
        weights1[20645] <= 16'b1111111111110001;
        weights1[20646] <= 16'b1111111111101101;
        weights1[20647] <= 16'b1111111111010010;
        weights1[20648] <= 16'b1111111111100000;
        weights1[20649] <= 16'b1111111111111110;
        weights1[20650] <= 16'b1111111111101100;
        weights1[20651] <= 16'b1111111111011010;
        weights1[20652] <= 16'b1111111111111010;
        weights1[20653] <= 16'b1111111111100100;
        weights1[20654] <= 16'b1111111111100111;
        weights1[20655] <= 16'b1111111111101010;
        weights1[20656] <= 16'b1111111111111011;
        weights1[20657] <= 16'b1111111111110010;
        weights1[20658] <= 16'b1111111111110101;
        weights1[20659] <= 16'b1111111111110000;
        weights1[20660] <= 16'b0000000000000010;
        weights1[20661] <= 16'b0000000000001110;
        weights1[20662] <= 16'b1111111111110001;
        weights1[20663] <= 16'b1111111111010110;
        weights1[20664] <= 16'b1111111111101100;
        weights1[20665] <= 16'b1111111111100000;
        weights1[20666] <= 16'b1111111111100111;
        weights1[20667] <= 16'b1111111111010101;
        weights1[20668] <= 16'b1111111111001111;
        weights1[20669] <= 16'b1111111111001111;
        weights1[20670] <= 16'b1111111111010101;
        weights1[20671] <= 16'b1111111111001111;
        weights1[20672] <= 16'b1111111110110100;
        weights1[20673] <= 16'b1111111111001110;
        weights1[20674] <= 16'b1111111111000110;
        weights1[20675] <= 16'b1111111111010111;
        weights1[20676] <= 16'b1111111111010011;
        weights1[20677] <= 16'b1111111111001111;
        weights1[20678] <= 16'b1111111111010111;
        weights1[20679] <= 16'b1111111111010100;
        weights1[20680] <= 16'b1111111111101011;
        weights1[20681] <= 16'b1111111111110000;
        weights1[20682] <= 16'b1111111111101111;
        weights1[20683] <= 16'b1111111111100110;
        weights1[20684] <= 16'b1111111111010000;
        weights1[20685] <= 16'b1111111111111101;
        weights1[20686] <= 16'b1111111111110000;
        weights1[20687] <= 16'b1111111111011101;
        weights1[20688] <= 16'b1111111111100000;
        weights1[20689] <= 16'b1111111111111010;
        weights1[20690] <= 16'b1111111111100010;
        weights1[20691] <= 16'b1111111111001111;
        weights1[20692] <= 16'b1111111111101100;
        weights1[20693] <= 16'b1111111111011111;
        weights1[20694] <= 16'b1111111111001010;
        weights1[20695] <= 16'b1111111110111011;
        weights1[20696] <= 16'b1111111111100000;
        weights1[20697] <= 16'b1111111111101100;
        weights1[20698] <= 16'b1111111111001110;
        weights1[20699] <= 16'b1111111111100111;
        weights1[20700] <= 16'b1111111111010010;
        weights1[20701] <= 16'b1111111111000000;
        weights1[20702] <= 16'b1111111111001011;
        weights1[20703] <= 16'b1111111111011011;
        weights1[20704] <= 16'b1111111111010100;
        weights1[20705] <= 16'b1111111111001011;
        weights1[20706] <= 16'b1111111111000011;
        weights1[20707] <= 16'b1111111111000010;
        weights1[20708] <= 16'b1111111111001100;
        weights1[20709] <= 16'b1111111111010011;
        weights1[20710] <= 16'b1111111111000001;
        weights1[20711] <= 16'b1111111111100000;
        weights1[20712] <= 16'b1111111111001110;
        weights1[20713] <= 16'b1111111111010100;
        weights1[20714] <= 16'b1111111111010010;
        weights1[20715] <= 16'b1111111111100010;
        weights1[20716] <= 16'b1111111111001111;
        weights1[20717] <= 16'b1111111111100001;
        weights1[20718] <= 16'b1111111111001100;
        weights1[20719] <= 16'b1111111111010010;
        weights1[20720] <= 16'b1111111111101011;
        weights1[20721] <= 16'b1111111111100100;
        weights1[20722] <= 16'b1111111111001111;
        weights1[20723] <= 16'b1111111111011001;
        weights1[20724] <= 16'b1111111111010100;
        weights1[20725] <= 16'b1111111111110111;
        weights1[20726] <= 16'b1111111111010100;
        weights1[20727] <= 16'b1111111111011011;
        weights1[20728] <= 16'b1111111111111010;
        weights1[20729] <= 16'b1111111111000111;
        weights1[20730] <= 16'b1111111111101001;
        weights1[20731] <= 16'b1111111111001100;
        weights1[20732] <= 16'b1111111111010111;
        weights1[20733] <= 16'b1111111110110101;
        weights1[20734] <= 16'b1111111110101110;
        weights1[20735] <= 16'b1111111110101100;
        weights1[20736] <= 16'b1111111111010101;
        weights1[20737] <= 16'b1111111111001010;
        weights1[20738] <= 16'b1111111111001010;
        weights1[20739] <= 16'b1111111111011010;
        weights1[20740] <= 16'b1111111111100110;
        weights1[20741] <= 16'b1111111110111111;
        weights1[20742] <= 16'b1111111111000010;
        weights1[20743] <= 16'b1111111110111011;
        weights1[20744] <= 16'b1111111111001101;
        weights1[20745] <= 16'b1111111111000001;
        weights1[20746] <= 16'b1111111111000001;
        weights1[20747] <= 16'b1111111111000100;
        weights1[20748] <= 16'b1111111111101110;
        weights1[20749] <= 16'b1111111111101110;
        weights1[20750] <= 16'b1111111111101011;
        weights1[20751] <= 16'b1111111111101101;
        weights1[20752] <= 16'b1111111111110001;
        weights1[20753] <= 16'b1111111111110000;
        weights1[20754] <= 16'b1111111111111010;
        weights1[20755] <= 16'b1111111111010110;
        weights1[20756] <= 16'b0000000000000100;
        weights1[20757] <= 16'b0000000000000011;
        weights1[20758] <= 16'b0000000000000001;
        weights1[20759] <= 16'b1111111111101101;
        weights1[20760] <= 16'b1111111111111000;
        weights1[20761] <= 16'b1111111111101110;
        weights1[20762] <= 16'b1111111111101101;
        weights1[20763] <= 16'b1111111111011111;
        weights1[20764] <= 16'b1111111111010111;
        weights1[20765] <= 16'b1111111111001001;
        weights1[20766] <= 16'b1111111110111110;
        weights1[20767] <= 16'b1111111111010000;
        weights1[20768] <= 16'b1111111110111111;
        weights1[20769] <= 16'b1111111110111001;
        weights1[20770] <= 16'b1111111110110101;
        weights1[20771] <= 16'b1111111110110011;
        weights1[20772] <= 16'b1111111111011000;
        weights1[20773] <= 16'b1111111110110111;
        weights1[20774] <= 16'b1111111111000100;
        weights1[20775] <= 16'b1111111111000100;
        weights1[20776] <= 16'b1111111111111011;
        weights1[20777] <= 16'b1111111111110101;
        weights1[20778] <= 16'b0000000000000100;
        weights1[20779] <= 16'b0000000000000111;
        weights1[20780] <= 16'b0000000000100010;
        weights1[20781] <= 16'b0000000000011011;
        weights1[20782] <= 16'b1111111111111110;
        weights1[20783] <= 16'b0000000000100001;
        weights1[20784] <= 16'b1111111111111011;
        weights1[20785] <= 16'b0000000000001010;
        weights1[20786] <= 16'b0000000000010000;
        weights1[20787] <= 16'b0000000000000001;
        weights1[20788] <= 16'b0000000000010100;
        weights1[20789] <= 16'b0000000000000010;
        weights1[20790] <= 16'b0000000000000011;
        weights1[20791] <= 16'b0000000000000111;
        weights1[20792] <= 16'b0000000000000111;
        weights1[20793] <= 16'b1111111111101101;
        weights1[20794] <= 16'b1111111111100001;
        weights1[20795] <= 16'b1111111111001000;
        weights1[20796] <= 16'b1111111111001111;
        weights1[20797] <= 16'b1111111111000001;
        weights1[20798] <= 16'b1111111111010101;
        weights1[20799] <= 16'b1111111110111101;
        weights1[20800] <= 16'b1111111110110001;
        weights1[20801] <= 16'b1111111110111000;
        weights1[20802] <= 16'b1111111111001000;
        weights1[20803] <= 16'b1111111111010000;
        weights1[20804] <= 16'b0000000000001011;
        weights1[20805] <= 16'b0000000000011010;
        weights1[20806] <= 16'b0000000000011010;
        weights1[20807] <= 16'b0000000000101111;
        weights1[20808] <= 16'b0000000000011011;
        weights1[20809] <= 16'b0000000000111001;
        weights1[20810] <= 16'b0000000000101110;
        weights1[20811] <= 16'b0000000000101111;
        weights1[20812] <= 16'b0000000000100001;
        weights1[20813] <= 16'b0000000000100100;
        weights1[20814] <= 16'b0000000000101010;
        weights1[20815] <= 16'b0000000000110011;
        weights1[20816] <= 16'b0000000000101010;
        weights1[20817] <= 16'b0000000000011011;
        weights1[20818] <= 16'b0000000000001010;
        weights1[20819] <= 16'b0000000000010000;
        weights1[20820] <= 16'b0000000000010011;
        weights1[20821] <= 16'b0000000000100011;
        weights1[20822] <= 16'b1111111111110100;
        weights1[20823] <= 16'b0000000000001100;
        weights1[20824] <= 16'b1111111111111001;
        weights1[20825] <= 16'b1111111111100101;
        weights1[20826] <= 16'b1111111111100100;
        weights1[20827] <= 16'b1111111111100000;
        weights1[20828] <= 16'b1111111111111100;
        weights1[20829] <= 16'b1111111111100111;
        weights1[20830] <= 16'b1111111111011111;
        weights1[20831] <= 16'b1111111111011010;
        weights1[20832] <= 16'b0000000000010011;
        weights1[20833] <= 16'b0000000000100010;
        weights1[20834] <= 16'b0000000000100110;
        weights1[20835] <= 16'b0000000001001001;
        weights1[20836] <= 16'b0000000000110111;
        weights1[20837] <= 16'b0000000000101011;
        weights1[20838] <= 16'b0000000000110110;
        weights1[20839] <= 16'b0000000000100111;
        weights1[20840] <= 16'b0000000000101111;
        weights1[20841] <= 16'b0000000000110110;
        weights1[20842] <= 16'b0000000000110100;
        weights1[20843] <= 16'b0000000000111000;
        weights1[20844] <= 16'b0000000000101010;
        weights1[20845] <= 16'b0000000000100111;
        weights1[20846] <= 16'b0000000000101100;
        weights1[20847] <= 16'b0000000000101111;
        weights1[20848] <= 16'b0000000000100001;
        weights1[20849] <= 16'b0000000000101010;
        weights1[20850] <= 16'b0000000000100001;
        weights1[20851] <= 16'b0000000000011010;
        weights1[20852] <= 16'b0000000000101011;
        weights1[20853] <= 16'b0000000001010001;
        weights1[20854] <= 16'b0000000000100110;
        weights1[20855] <= 16'b0000000000010101;
        weights1[20856] <= 16'b0000000000010110;
        weights1[20857] <= 16'b0000000000010010;
        weights1[20858] <= 16'b1111111111111100;
        weights1[20859] <= 16'b1111111111111101;
        weights1[20860] <= 16'b0000000000011110;
        weights1[20861] <= 16'b0000000000110011;
        weights1[20862] <= 16'b0000000000101100;
        weights1[20863] <= 16'b0000000000110111;
        weights1[20864] <= 16'b0000000000011111;
        weights1[20865] <= 16'b0000000000110010;
        weights1[20866] <= 16'b0000000001000000;
        weights1[20867] <= 16'b0000000000100110;
        weights1[20868] <= 16'b0000000001001001;
        weights1[20869] <= 16'b0000000000100110;
        weights1[20870] <= 16'b0000000000101111;
        weights1[20871] <= 16'b0000000000101010;
        weights1[20872] <= 16'b0000000000110010;
        weights1[20873] <= 16'b0000000000110011;
        weights1[20874] <= 16'b0000000000110101;
        weights1[20875] <= 16'b0000000000111010;
        weights1[20876] <= 16'b0000000000110111;
        weights1[20877] <= 16'b0000000000110110;
        weights1[20878] <= 16'b0000000000111010;
        weights1[20879] <= 16'b0000000000101010;
        weights1[20880] <= 16'b0000000000101100;
        weights1[20881] <= 16'b0000000000011011;
        weights1[20882] <= 16'b0000000000011110;
        weights1[20883] <= 16'b0000000001000000;
        weights1[20884] <= 16'b0000000000110111;
        weights1[20885] <= 16'b0000000001001110;
        weights1[20886] <= 16'b0000000000100001;
        weights1[20887] <= 16'b0000000000011001;
        weights1[20888] <= 16'b0000000000100101;
        weights1[20889] <= 16'b0000000000101100;
        weights1[20890] <= 16'b0000000000010110;
        weights1[20891] <= 16'b0000000000011110;
        weights1[20892] <= 16'b0000000000101001;
        weights1[20893] <= 16'b0000000000101110;
        weights1[20894] <= 16'b0000000000011101;
        weights1[20895] <= 16'b0000000000011010;
        weights1[20896] <= 16'b0000000000011000;
        weights1[20897] <= 16'b0000000000010001;
        weights1[20898] <= 16'b0000000000001100;
        weights1[20899] <= 16'b0000000000010110;
        weights1[20900] <= 16'b0000000000010111;
        weights1[20901] <= 16'b0000000000011001;
        weights1[20902] <= 16'b0000000000011011;
        weights1[20903] <= 16'b0000000000101010;
        weights1[20904] <= 16'b0000000001000110;
        weights1[20905] <= 16'b0000000000111111;
        weights1[20906] <= 16'b0000000000100101;
        weights1[20907] <= 16'b0000000000101101;
        weights1[20908] <= 16'b0000000000111100;
        weights1[20909] <= 16'b0000000000101001;
        weights1[20910] <= 16'b0000000000100110;
        weights1[20911] <= 16'b0000000001001101;
        weights1[20912] <= 16'b0000000001100001;
        weights1[20913] <= 16'b0000000001001000;
        weights1[20914] <= 16'b0000000001000011;
        weights1[20915] <= 16'b0000000000111100;
        weights1[20916] <= 16'b0000000000100001;
        weights1[20917] <= 16'b0000000000011101;
        weights1[20918] <= 16'b0000000000000111;
        weights1[20919] <= 16'b0000000000010011;
        weights1[20920] <= 16'b0000000000011100;
        weights1[20921] <= 16'b0000000000000111;
        weights1[20922] <= 16'b0000000000001101;
        weights1[20923] <= 16'b0000000000000011;
        weights1[20924] <= 16'b0000000000011000;
        weights1[20925] <= 16'b0000000000011010;
        weights1[20926] <= 16'b0000000000100000;
        weights1[20927] <= 16'b1111111111110111;
        weights1[20928] <= 16'b0000000000001011;
        weights1[20929] <= 16'b0000000000110011;
        weights1[20930] <= 16'b0000000000011010;
        weights1[20931] <= 16'b0000000000110011;
        weights1[20932] <= 16'b0000000000101111;
        weights1[20933] <= 16'b0000000001000101;
        weights1[20934] <= 16'b0000000000110111;
        weights1[20935] <= 16'b0000000001001001;
        weights1[20936] <= 16'b0000000000110000;
        weights1[20937] <= 16'b0000000001000011;
        weights1[20938] <= 16'b0000000000111111;
        weights1[20939] <= 16'b0000000000111000;
        weights1[20940] <= 16'b0000000001000100;
        weights1[20941] <= 16'b0000000001010110;
        weights1[20942] <= 16'b0000000001010100;
        weights1[20943] <= 16'b0000000001000000;
        weights1[20944] <= 16'b0000000000001001;
        weights1[20945] <= 16'b0000000000001100;
        weights1[20946] <= 16'b1111111111111101;
        weights1[20947] <= 16'b0000000000000010;
        weights1[20948] <= 16'b0000000000010010;
        weights1[20949] <= 16'b1111111111100000;
        weights1[20950] <= 16'b0000000000011000;
        weights1[20951] <= 16'b0000000000010000;
        weights1[20952] <= 16'b0000000000001011;
        weights1[20953] <= 16'b0000000000011011;
        weights1[20954] <= 16'b0000000000001000;
        weights1[20955] <= 16'b0000000000100001;
        weights1[20956] <= 16'b1111111111110101;
        weights1[20957] <= 16'b0000000000000100;
        weights1[20958] <= 16'b0000000000010000;
        weights1[20959] <= 16'b0000000000001010;
        weights1[20960] <= 16'b0000000000010101;
        weights1[20961] <= 16'b0000000000100000;
        weights1[20962] <= 16'b0000000000111101;
        weights1[20963] <= 16'b0000000001000001;
        weights1[20964] <= 16'b0000000001010110;
        weights1[20965] <= 16'b0000000001000000;
        weights1[20966] <= 16'b0000000000110001;
        weights1[20967] <= 16'b0000000000110111;
        weights1[20968] <= 16'b0000000001000110;
        weights1[20969] <= 16'b0000000000110110;
        weights1[20970] <= 16'b0000000001000100;
        weights1[20971] <= 16'b0000000000101000;
        weights1[20972] <= 16'b1111111111110100;
        weights1[20973] <= 16'b0000000000000111;
        weights1[20974] <= 16'b1111111111110001;
        weights1[20975] <= 16'b1111111111101011;
        weights1[20976] <= 16'b1111111111101110;
        weights1[20977] <= 16'b0000000000100101;
        weights1[20978] <= 16'b0000000000001110;
        weights1[20979] <= 16'b1111111111111011;
        weights1[20980] <= 16'b0000000000000101;
        weights1[20981] <= 16'b0000000000000111;
        weights1[20982] <= 16'b0000000000000110;
        weights1[20983] <= 16'b0000000000000010;
        weights1[20984] <= 16'b0000000000001000;
        weights1[20985] <= 16'b0000000000000011;
        weights1[20986] <= 16'b1111111111111011;
        weights1[20987] <= 16'b1111111111110011;
        weights1[20988] <= 16'b0000000000000010;
        weights1[20989] <= 16'b0000000000000001;
        weights1[20990] <= 16'b1111111111100000;
        weights1[20991] <= 16'b0000000000000110;
        weights1[20992] <= 16'b0000000000101100;
        weights1[20993] <= 16'b0000000000001101;
        weights1[20994] <= 16'b0000000000100011;
        weights1[20995] <= 16'b0000000000101001;
        weights1[20996] <= 16'b0000000000011101;
        weights1[20997] <= 16'b0000000000011010;
        weights1[20998] <= 16'b0000000000011010;
        weights1[20999] <= 16'b0000000000001001;
        weights1[21000] <= 16'b1111111111111000;
        weights1[21001] <= 16'b1111111111110111;
        weights1[21002] <= 16'b1111111111110001;
        weights1[21003] <= 16'b1111111111101110;
        weights1[21004] <= 16'b1111111111111101;
        weights1[21005] <= 16'b0000000000001011;
        weights1[21006] <= 16'b1111111111011111;
        weights1[21007] <= 16'b1111111111111010;
        weights1[21008] <= 16'b0000000000001000;
        weights1[21009] <= 16'b1111111111110000;
        weights1[21010] <= 16'b1111111111111101;
        weights1[21011] <= 16'b0000000000001011;
        weights1[21012] <= 16'b1111111111101101;
        weights1[21013] <= 16'b0000000000001010;
        weights1[21014] <= 16'b1111111111110010;
        weights1[21015] <= 16'b1111111111101100;
        weights1[21016] <= 16'b1111111111101000;
        weights1[21017] <= 16'b1111111111100110;
        weights1[21018] <= 16'b1111111111011010;
        weights1[21019] <= 16'b1111111111101011;
        weights1[21020] <= 16'b0000000000001000;
        weights1[21021] <= 16'b1111111111110110;
        weights1[21022] <= 16'b0000000000010001;
        weights1[21023] <= 16'b1111111111101111;
        weights1[21024] <= 16'b1111111111100110;
        weights1[21025] <= 16'b1111111111111000;
        weights1[21026] <= 16'b1111111111111000;
        weights1[21027] <= 16'b1111111111110111;
        weights1[21028] <= 16'b1111111111111001;
        weights1[21029] <= 16'b1111111111101010;
        weights1[21030] <= 16'b1111111111101110;
        weights1[21031] <= 16'b1111111111101011;
        weights1[21032] <= 16'b1111111111100011;
        weights1[21033] <= 16'b0000000000000000;
        weights1[21034] <= 16'b1111111111101110;
        weights1[21035] <= 16'b1111111111110001;
        weights1[21036] <= 16'b1111111111110110;
        weights1[21037] <= 16'b1111111111101010;
        weights1[21038] <= 16'b1111111111111001;
        weights1[21039] <= 16'b0000000000001001;
        weights1[21040] <= 16'b0000000000000000;
        weights1[21041] <= 16'b1111111111110100;
        weights1[21042] <= 16'b1111111111110011;
        weights1[21043] <= 16'b1111111111111000;
        weights1[21044] <= 16'b1111111111100100;
        weights1[21045] <= 16'b1111111111011110;
        weights1[21046] <= 16'b1111111111100101;
        weights1[21047] <= 16'b1111111111100101;
        weights1[21048] <= 16'b1111111111010110;
        weights1[21049] <= 16'b1111111111100111;
        weights1[21050] <= 16'b1111111111011100;
        weights1[21051] <= 16'b1111111111011101;
        weights1[21052] <= 16'b1111111111001111;
        weights1[21053] <= 16'b1111111111011101;
        weights1[21054] <= 16'b1111111111110001;
        weights1[21055] <= 16'b1111111111110100;
        weights1[21056] <= 16'b1111111111111001;
        weights1[21057] <= 16'b1111111111110001;
        weights1[21058] <= 16'b1111111111101110;
        weights1[21059] <= 16'b1111111111100100;
        weights1[21060] <= 16'b1111111111101110;
        weights1[21061] <= 16'b1111111111101101;
        weights1[21062] <= 16'b1111111111010001;
        weights1[21063] <= 16'b1111111111110010;
        weights1[21064] <= 16'b1111111111100111;
        weights1[21065] <= 16'b1111111111111010;
        weights1[21066] <= 16'b0000000000010010;
        weights1[21067] <= 16'b1111111111110000;
        weights1[21068] <= 16'b1111111111111011;
        weights1[21069] <= 16'b1111111111110001;
        weights1[21070] <= 16'b1111111111110000;
        weights1[21071] <= 16'b0000000000001111;
        weights1[21072] <= 16'b1111111111101110;
        weights1[21073] <= 16'b1111111111111011;
        weights1[21074] <= 16'b1111111111101110;
        weights1[21075] <= 16'b1111111111001100;
        weights1[21076] <= 16'b1111111111010110;
        weights1[21077] <= 16'b1111111111001001;
        weights1[21078] <= 16'b1111111111001010;
        weights1[21079] <= 16'b1111111111000101;
        weights1[21080] <= 16'b1111111111011011;
        weights1[21081] <= 16'b1111111111100010;
        weights1[21082] <= 16'b1111111111100110;
        weights1[21083] <= 16'b1111111111110011;
        weights1[21084] <= 16'b1111111111111101;
        weights1[21085] <= 16'b1111111111111000;
        weights1[21086] <= 16'b1111111111110011;
        weights1[21087] <= 16'b1111111111101101;
        weights1[21088] <= 16'b1111111111101000;
        weights1[21089] <= 16'b1111111111101001;
        weights1[21090] <= 16'b1111111111010100;
        weights1[21091] <= 16'b1111111111011010;
        weights1[21092] <= 16'b1111111111100011;
        weights1[21093] <= 16'b1111111111011011;
        weights1[21094] <= 16'b1111111111100101;
        weights1[21095] <= 16'b1111111111011011;
        weights1[21096] <= 16'b1111111111110111;
        weights1[21097] <= 16'b1111111111101010;
        weights1[21098] <= 16'b1111111111100010;
        weights1[21099] <= 16'b1111111111011010;
        weights1[21100] <= 16'b1111111111011111;
        weights1[21101] <= 16'b1111111111100110;
        weights1[21102] <= 16'b1111111111101101;
        weights1[21103] <= 16'b1111111111000001;
        weights1[21104] <= 16'b1111111111001100;
        weights1[21105] <= 16'b1111111111001010;
        weights1[21106] <= 16'b1111111111000110;
        weights1[21107] <= 16'b1111111111001011;
        weights1[21108] <= 16'b1111111111000110;
        weights1[21109] <= 16'b1111111111011100;
        weights1[21110] <= 16'b1111111111101010;
        weights1[21111] <= 16'b1111111111111000;
        weights1[21112] <= 16'b1111111111111100;
        weights1[21113] <= 16'b1111111111111011;
        weights1[21114] <= 16'b1111111111110101;
        weights1[21115] <= 16'b1111111111110010;
        weights1[21116] <= 16'b1111111111101011;
        weights1[21117] <= 16'b1111111111100110;
        weights1[21118] <= 16'b1111111111011001;
        weights1[21119] <= 16'b1111111111101001;
        weights1[21120] <= 16'b1111111111011101;
        weights1[21121] <= 16'b1111111111100111;
        weights1[21122] <= 16'b1111111111100101;
        weights1[21123] <= 16'b1111111111100110;
        weights1[21124] <= 16'b1111111111101010;
        weights1[21125] <= 16'b1111111111100000;
        weights1[21126] <= 16'b1111111111101100;
        weights1[21127] <= 16'b1111111111110001;
        weights1[21128] <= 16'b1111111111010110;
        weights1[21129] <= 16'b1111111111100111;
        weights1[21130] <= 16'b1111111111100100;
        weights1[21131] <= 16'b1111111111011100;
        weights1[21132] <= 16'b1111111111100001;
        weights1[21133] <= 16'b1111111111010010;
        weights1[21134] <= 16'b1111111111010101;
        weights1[21135] <= 16'b1111111111011100;
        weights1[21136] <= 16'b1111111111011101;
        weights1[21137] <= 16'b1111111111100101;
        weights1[21138] <= 16'b1111111111110000;
        weights1[21139] <= 16'b1111111111111000;
        weights1[21140] <= 16'b1111111111111111;
        weights1[21141] <= 16'b1111111111111110;
        weights1[21142] <= 16'b1111111111111001;
        weights1[21143] <= 16'b1111111111111101;
        weights1[21144] <= 16'b1111111111101111;
        weights1[21145] <= 16'b1111111111101000;
        weights1[21146] <= 16'b1111111111100110;
        weights1[21147] <= 16'b1111111111011011;
        weights1[21148] <= 16'b1111111111011100;
        weights1[21149] <= 16'b1111111111100001;
        weights1[21150] <= 16'b1111111111011010;
        weights1[21151] <= 16'b1111111111110000;
        weights1[21152] <= 16'b1111111111100011;
        weights1[21153] <= 16'b1111111111001100;
        weights1[21154] <= 16'b1111111111001111;
        weights1[21155] <= 16'b1111111111010010;
        weights1[21156] <= 16'b1111111111010111;
        weights1[21157] <= 16'b1111111111100100;
        weights1[21158] <= 16'b1111111111010101;
        weights1[21159] <= 16'b1111111111010000;
        weights1[21160] <= 16'b1111111111100000;
        weights1[21161] <= 16'b1111111111010001;
        weights1[21162] <= 16'b1111111111011101;
        weights1[21163] <= 16'b1111111111100110;
        weights1[21164] <= 16'b1111111111100111;
        weights1[21165] <= 16'b1111111111110001;
        weights1[21166] <= 16'b1111111111110111;
        weights1[21167] <= 16'b1111111111111101;
        weights1[21168] <= 16'b0000000000000000;
        weights1[21169] <= 16'b0000000000000000;
        weights1[21170] <= 16'b1111111111111101;
        weights1[21171] <= 16'b0000000000000000;
        weights1[21172] <= 16'b0000000000000001;
        weights1[21173] <= 16'b0000000000000000;
        weights1[21174] <= 16'b1111111111111110;
        weights1[21175] <= 16'b1111111111111011;
        weights1[21176] <= 16'b1111111111111010;
        weights1[21177] <= 16'b1111111111111100;
        weights1[21178] <= 16'b0000000000001000;
        weights1[21179] <= 16'b1111111111111011;
        weights1[21180] <= 16'b0000000000000110;
        weights1[21181] <= 16'b1111111111110110;
        weights1[21182] <= 16'b1111111111101011;
        weights1[21183] <= 16'b1111111111110110;
        weights1[21184] <= 16'b1111111111111011;
        weights1[21185] <= 16'b0000000000010010;
        weights1[21186] <= 16'b0000000000001001;
        weights1[21187] <= 16'b1111111111110111;
        weights1[21188] <= 16'b1111111111111000;
        weights1[21189] <= 16'b0000000000001001;
        weights1[21190] <= 16'b0000000000001100;
        weights1[21191] <= 16'b0000000000001010;
        weights1[21192] <= 16'b0000000000001111;
        weights1[21193] <= 16'b0000000000001001;
        weights1[21194] <= 16'b0000000000000001;
        weights1[21195] <= 16'b0000000000000010;
        weights1[21196] <= 16'b0000000000000001;
        weights1[21197] <= 16'b0000000000000000;
        weights1[21198] <= 16'b0000000000000001;
        weights1[21199] <= 16'b1111111111111110;
        weights1[21200] <= 16'b0000000000000011;
        weights1[21201] <= 16'b0000000000000011;
        weights1[21202] <= 16'b0000000000000001;
        weights1[21203] <= 16'b1111111111110100;
        weights1[21204] <= 16'b1111111111110011;
        weights1[21205] <= 16'b0000000000000110;
        weights1[21206] <= 16'b1111111111110011;
        weights1[21207] <= 16'b1111111111110001;
        weights1[21208] <= 16'b0000000000000000;
        weights1[21209] <= 16'b1111111111111100;
        weights1[21210] <= 16'b0000000000000001;
        weights1[21211] <= 16'b1111111111111110;
        weights1[21212] <= 16'b0000000000000011;
        weights1[21213] <= 16'b1111111111111111;
        weights1[21214] <= 16'b0000000000000011;
        weights1[21215] <= 16'b1111111111110111;
        weights1[21216] <= 16'b1111111111111011;
        weights1[21217] <= 16'b0000000000000010;
        weights1[21218] <= 16'b0000000000001100;
        weights1[21219] <= 16'b0000000000000011;
        weights1[21220] <= 16'b0000000000001000;
        weights1[21221] <= 16'b0000000000001010;
        weights1[21222] <= 16'b0000000000000001;
        weights1[21223] <= 16'b0000000000000100;
        weights1[21224] <= 16'b0000000000000000;
        weights1[21225] <= 16'b0000000000000010;
        weights1[21226] <= 16'b1111111111111110;
        weights1[21227] <= 16'b0000000000001010;
        weights1[21228] <= 16'b0000000000001011;
        weights1[21229] <= 16'b0000000000001111;
        weights1[21230] <= 16'b0000000000011101;
        weights1[21231] <= 16'b0000000000001001;
        weights1[21232] <= 16'b0000000000000001;
        weights1[21233] <= 16'b1111111111101101;
        weights1[21234] <= 16'b1111111111110101;
        weights1[21235] <= 16'b1111111111111001;
        weights1[21236] <= 16'b0000000000000011;
        weights1[21237] <= 16'b1111111111111001;
        weights1[21238] <= 16'b1111111111111100;
        weights1[21239] <= 16'b0000000000001100;
        weights1[21240] <= 16'b1111111111111000;
        weights1[21241] <= 16'b1111111111110110;
        weights1[21242] <= 16'b0000000000010000;
        weights1[21243] <= 16'b0000000000000110;
        weights1[21244] <= 16'b0000000000001101;
        weights1[21245] <= 16'b0000000000001100;
        weights1[21246] <= 16'b0000000000001000;
        weights1[21247] <= 16'b0000000000000111;
        weights1[21248] <= 16'b0000000000000011;
        weights1[21249] <= 16'b0000000000000110;
        weights1[21250] <= 16'b0000000000001011;
        weights1[21251] <= 16'b0000000000001000;
        weights1[21252] <= 16'b0000000000000010;
        weights1[21253] <= 16'b0000000000000011;
        weights1[21254] <= 16'b0000000000000111;
        weights1[21255] <= 16'b0000000000001111;
        weights1[21256] <= 16'b0000000000011111;
        weights1[21257] <= 16'b0000000000100111;
        weights1[21258] <= 16'b0000000000010111;
        weights1[21259] <= 16'b0000000000011011;
        weights1[21260] <= 16'b0000000000001000;
        weights1[21261] <= 16'b1111111111111111;
        weights1[21262] <= 16'b1111111111111100;
        weights1[21263] <= 16'b0000000000000011;
        weights1[21264] <= 16'b1111111111111100;
        weights1[21265] <= 16'b1111111111110011;
        weights1[21266] <= 16'b0000000000000010;
        weights1[21267] <= 16'b0000000000000111;
        weights1[21268] <= 16'b1111111111110101;
        weights1[21269] <= 16'b1111111111101111;
        weights1[21270] <= 16'b0000000000001011;
        weights1[21271] <= 16'b1111111111111010;
        weights1[21272] <= 16'b1111111111110101;
        weights1[21273] <= 16'b1111111111101000;
        weights1[21274] <= 16'b0000000000000001;
        weights1[21275] <= 16'b1111111111111110;
        weights1[21276] <= 16'b0000000000001011;
        weights1[21277] <= 16'b0000000000000001;
        weights1[21278] <= 16'b0000000000001010;
        weights1[21279] <= 16'b0000000000001010;
        weights1[21280] <= 16'b0000000000000001;
        weights1[21281] <= 16'b0000000000001000;
        weights1[21282] <= 16'b0000000000010001;
        weights1[21283] <= 16'b0000000000011101;
        weights1[21284] <= 16'b0000000000110010;
        weights1[21285] <= 16'b0000000000110011;
        weights1[21286] <= 16'b0000000000010101;
        weights1[21287] <= 16'b0000000000101100;
        weights1[21288] <= 16'b0000000000100111;
        weights1[21289] <= 16'b0000000000010000;
        weights1[21290] <= 16'b0000000000001010;
        weights1[21291] <= 16'b0000000000010100;
        weights1[21292] <= 16'b0000000000001101;
        weights1[21293] <= 16'b1111111111111101;
        weights1[21294] <= 16'b1111111111110101;
        weights1[21295] <= 16'b0000000000000001;
        weights1[21296] <= 16'b0000000000001110;
        weights1[21297] <= 16'b0000000000000010;
        weights1[21298] <= 16'b0000000000000001;
        weights1[21299] <= 16'b1111111111101000;
        weights1[21300] <= 16'b0000000000000011;
        weights1[21301] <= 16'b1111111111111101;
        weights1[21302] <= 16'b1111111111110001;
        weights1[21303] <= 16'b1111111111111100;
        weights1[21304] <= 16'b0000000000001010;
        weights1[21305] <= 16'b1111111111111000;
        weights1[21306] <= 16'b1111111111111101;
        weights1[21307] <= 16'b0000000000000001;
        weights1[21308] <= 16'b0000000000000101;
        weights1[21309] <= 16'b0000000000001111;
        weights1[21310] <= 16'b0000000000011011;
        weights1[21311] <= 16'b0000000000101001;
        weights1[21312] <= 16'b0000000000100010;
        weights1[21313] <= 16'b0000000000110011;
        weights1[21314] <= 16'b0000000000100000;
        weights1[21315] <= 16'b0000000000101000;
        weights1[21316] <= 16'b0000000000011001;
        weights1[21317] <= 16'b0000000000000110;
        weights1[21318] <= 16'b0000000000011011;
        weights1[21319] <= 16'b0000000000001000;
        weights1[21320] <= 16'b0000000000001001;
        weights1[21321] <= 16'b0000000000001000;
        weights1[21322] <= 16'b0000000000001100;
        weights1[21323] <= 16'b0000000000000101;
        weights1[21324] <= 16'b0000000000000100;
        weights1[21325] <= 16'b0000000000000100;
        weights1[21326] <= 16'b1111111111110011;
        weights1[21327] <= 16'b1111111111111110;
        weights1[21328] <= 16'b0000000000000111;
        weights1[21329] <= 16'b1111111111110001;
        weights1[21330] <= 16'b1111111111110101;
        weights1[21331] <= 16'b0000000000000010;
        weights1[21332] <= 16'b1111111111110110;
        weights1[21333] <= 16'b1111111111101111;
        weights1[21334] <= 16'b0000000000000000;
        weights1[21335] <= 16'b1111111111111101;
        weights1[21336] <= 16'b0000000000001011;
        weights1[21337] <= 16'b0000000000011100;
        weights1[21338] <= 16'b0000000000011000;
        weights1[21339] <= 16'b0000000000011111;
        weights1[21340] <= 16'b0000000000110000;
        weights1[21341] <= 16'b0000000000101110;
        weights1[21342] <= 16'b0000000000011110;
        weights1[21343] <= 16'b0000000000001011;
        weights1[21344] <= 16'b0000000000100111;
        weights1[21345] <= 16'b0000000000101101;
        weights1[21346] <= 16'b0000000000101100;
        weights1[21347] <= 16'b0000000000011100;
        weights1[21348] <= 16'b0000000000011110;
        weights1[21349] <= 16'b0000000000010011;
        weights1[21350] <= 16'b0000000000010010;
        weights1[21351] <= 16'b1111111111111011;
        weights1[21352] <= 16'b1111111111111100;
        weights1[21353] <= 16'b1111111111111101;
        weights1[21354] <= 16'b0000000000001001;
        weights1[21355] <= 16'b0000000000000110;
        weights1[21356] <= 16'b1111111111101101;
        weights1[21357] <= 16'b0000000000001001;
        weights1[21358] <= 16'b0000000000000010;
        weights1[21359] <= 16'b1111111111111110;
        weights1[21360] <= 16'b0000000000001000;
        weights1[21361] <= 16'b0000000000001101;
        weights1[21362] <= 16'b0000000000001010;
        weights1[21363] <= 16'b1111111111111000;
        weights1[21364] <= 16'b0000000000010011;
        weights1[21365] <= 16'b0000000000001111;
        weights1[21366] <= 16'b0000000000010000;
        weights1[21367] <= 16'b0000000000011010;
        weights1[21368] <= 16'b0000000000100100;
        weights1[21369] <= 16'b0000000000100011;
        weights1[21370] <= 16'b0000000000100110;
        weights1[21371] <= 16'b0000000000110010;
        weights1[21372] <= 16'b0000000000110011;
        weights1[21373] <= 16'b0000000000110000;
        weights1[21374] <= 16'b1111111111111100;
        weights1[21375] <= 16'b0000000000001111;
        weights1[21376] <= 16'b0000000000001001;
        weights1[21377] <= 16'b1111111111111001;
        weights1[21378] <= 16'b1111111111111101;
        weights1[21379] <= 16'b0000000000001011;
        weights1[21380] <= 16'b1111111111111010;
        weights1[21381] <= 16'b1111111111111011;
        weights1[21382] <= 16'b0000000000001111;
        weights1[21383] <= 16'b1111111111111011;
        weights1[21384] <= 16'b1111111111111101;
        weights1[21385] <= 16'b1111111111111000;
        weights1[21386] <= 16'b0000000000000011;
        weights1[21387] <= 16'b1111111111111100;
        weights1[21388] <= 16'b0000000000000010;
        weights1[21389] <= 16'b1111111111111001;
        weights1[21390] <= 16'b1111111111111000;
        weights1[21391] <= 16'b1111111111111110;
        weights1[21392] <= 16'b0000000000001110;
        weights1[21393] <= 16'b0000000000001001;
        weights1[21394] <= 16'b1111111111110000;
        weights1[21395] <= 16'b1111111111111011;
        weights1[21396] <= 16'b0000000000000011;
        weights1[21397] <= 16'b1111111111001111;
        weights1[21398] <= 16'b0000000000000111;
        weights1[21399] <= 16'b1111111111110110;
        weights1[21400] <= 16'b1111111111001111;
        weights1[21401] <= 16'b1111111111010011;
        weights1[21402] <= 16'b1111111111111111;
        weights1[21403] <= 16'b1111111111100001;
        weights1[21404] <= 16'b0000000000001010;
        weights1[21405] <= 16'b1111111111110011;
        weights1[21406] <= 16'b1111111111111011;
        weights1[21407] <= 16'b1111111111111000;
        weights1[21408] <= 16'b1111111111111001;
        weights1[21409] <= 16'b1111111111111000;
        weights1[21410] <= 16'b1111111111110001;
        weights1[21411] <= 16'b1111111111111001;
        weights1[21412] <= 16'b1111111111111111;
        weights1[21413] <= 16'b1111111111111111;
        weights1[21414] <= 16'b0000000000001000;
        weights1[21415] <= 16'b1111111111111101;
        weights1[21416] <= 16'b0000000000010011;
        weights1[21417] <= 16'b1111111111111011;
        weights1[21418] <= 16'b1111111111111110;
        weights1[21419] <= 16'b1111111111111110;
        weights1[21420] <= 16'b0000000000001001;
        weights1[21421] <= 16'b1111111111101010;
        weights1[21422] <= 16'b1111111111010010;
        weights1[21423] <= 16'b1111111111001110;
        weights1[21424] <= 16'b1111111111000111;
        weights1[21425] <= 16'b1111111110110010;
        weights1[21426] <= 16'b1111111110010101;
        weights1[21427] <= 16'b1111111110010111;
        weights1[21428] <= 16'b1111111110100101;
        weights1[21429] <= 16'b1111111110101001;
        weights1[21430] <= 16'b1111111111000100;
        weights1[21431] <= 16'b1111111111101100;
        weights1[21432] <= 16'b1111111111100111;
        weights1[21433] <= 16'b1111111111110100;
        weights1[21434] <= 16'b1111111111110001;
        weights1[21435] <= 16'b0000000000000100;
        weights1[21436] <= 16'b1111111111111101;
        weights1[21437] <= 16'b0000000000000110;
        weights1[21438] <= 16'b0000000000000000;
        weights1[21439] <= 16'b0000000000010011;
        weights1[21440] <= 16'b0000000000010010;
        weights1[21441] <= 16'b0000000000000101;
        weights1[21442] <= 16'b1111111111110110;
        weights1[21443] <= 16'b1111111111111010;
        weights1[21444] <= 16'b1111111111111011;
        weights1[21445] <= 16'b1111111111100101;
        weights1[21446] <= 16'b1111111111110100;
        weights1[21447] <= 16'b1111111111101011;
        weights1[21448] <= 16'b1111111111110010;
        weights1[21449] <= 16'b1111111111011011;
        weights1[21450] <= 16'b1111111111000010;
        weights1[21451] <= 16'b1111111110101111;
        weights1[21452] <= 16'b1111111110011000;
        weights1[21453] <= 16'b1111111110010100;
        weights1[21454] <= 16'b1111111110110010;
        weights1[21455] <= 16'b1111111111001010;
        weights1[21456] <= 16'b1111111111010010;
        weights1[21457] <= 16'b1111111111111110;
        weights1[21458] <= 16'b1111111111110010;
        weights1[21459] <= 16'b1111111111111000;
        weights1[21460] <= 16'b0000000000001010;
        weights1[21461] <= 16'b1111111111111100;
        weights1[21462] <= 16'b0000000000000101;
        weights1[21463] <= 16'b0000000000000001;
        weights1[21464] <= 16'b0000000000001101;
        weights1[21465] <= 16'b0000000000000110;
        weights1[21466] <= 16'b1111111111111011;
        weights1[21467] <= 16'b1111111111111111;
        weights1[21468] <= 16'b1111111111110000;
        weights1[21469] <= 16'b1111111111111011;
        weights1[21470] <= 16'b1111111111110101;
        weights1[21471] <= 16'b0000000000001100;
        weights1[21472] <= 16'b1111111111111010;
        weights1[21473] <= 16'b0000000000000010;
        weights1[21474] <= 16'b1111111111111111;
        weights1[21475] <= 16'b1111111111100111;
        weights1[21476] <= 16'b1111111111100111;
        weights1[21477] <= 16'b1111111111010111;
        weights1[21478] <= 16'b1111111111001110;
        weights1[21479] <= 16'b1111111111000000;
        weights1[21480] <= 16'b1111111111001101;
        weights1[21481] <= 16'b1111111111011100;
        weights1[21482] <= 16'b1111111111111011;
        weights1[21483] <= 16'b0000000000011000;
        weights1[21484] <= 16'b1111111111111011;
        weights1[21485] <= 16'b0000000000001100;
        weights1[21486] <= 16'b0000000000011000;
        weights1[21487] <= 16'b0000000000010010;
        weights1[21488] <= 16'b0000000000011101;
        weights1[21489] <= 16'b0000000000100010;
        weights1[21490] <= 16'b0000000000001011;
        weights1[21491] <= 16'b0000000000010101;
        weights1[21492] <= 16'b1111111111110000;
        weights1[21493] <= 16'b1111111111111011;
        weights1[21494] <= 16'b1111111111110100;
        weights1[21495] <= 16'b0000000000000001;
        weights1[21496] <= 16'b1111111111110011;
        weights1[21497] <= 16'b1111111111110100;
        weights1[21498] <= 16'b1111111111111100;
        weights1[21499] <= 16'b1111111111110000;
        weights1[21500] <= 16'b1111111111110100;
        weights1[21501] <= 16'b1111111111101010;
        weights1[21502] <= 16'b0000000000000010;
        weights1[21503] <= 16'b1111111111101000;
        weights1[21504] <= 16'b1111111111100100;
        weights1[21505] <= 16'b1111111111010010;
        weights1[21506] <= 16'b1111111111100101;
        weights1[21507] <= 16'b1111111111110101;
        weights1[21508] <= 16'b0000000000000100;
        weights1[21509] <= 16'b0000000000101010;
        weights1[21510] <= 16'b0000000000001001;
        weights1[21511] <= 16'b0000000000101100;
        weights1[21512] <= 16'b0000000000111100;
        weights1[21513] <= 16'b0000000000110000;
        weights1[21514] <= 16'b0000000000100100;
        weights1[21515] <= 16'b0000000000011011;
        weights1[21516] <= 16'b0000000000100011;
        weights1[21517] <= 16'b0000000000010101;
        weights1[21518] <= 16'b0000000000010010;
        weights1[21519] <= 16'b1111111111111000;
        weights1[21520] <= 16'b0000000000001010;
        weights1[21521] <= 16'b1111111111111001;
        weights1[21522] <= 16'b1111111111110010;
        weights1[21523] <= 16'b1111111111110001;
        weights1[21524] <= 16'b1111111111101111;
        weights1[21525] <= 16'b1111111111111100;
        weights1[21526] <= 16'b1111111111111000;
        weights1[21527] <= 16'b1111111111110000;
        weights1[21528] <= 16'b0000000000001100;
        weights1[21529] <= 16'b1111111111100111;
        weights1[21530] <= 16'b1111111111111000;
        weights1[21531] <= 16'b1111111111101011;
        weights1[21532] <= 16'b1111111111011100;
        weights1[21533] <= 16'b1111111111011001;
        weights1[21534] <= 16'b1111111111101100;
        weights1[21535] <= 16'b1111111111110110;
        weights1[21536] <= 16'b0000000000011101;
        weights1[21537] <= 16'b0000000000110110;
        weights1[21538] <= 16'b0000000000010100;
        weights1[21539] <= 16'b0000000000111011;
        weights1[21540] <= 16'b0000000000101010;
        weights1[21541] <= 16'b0000000000001001;
        weights1[21542] <= 16'b0000000000100100;
        weights1[21543] <= 16'b0000000000100010;
        weights1[21544] <= 16'b0000000000100000;
        weights1[21545] <= 16'b0000000000001100;
        weights1[21546] <= 16'b0000000000000101;
        weights1[21547] <= 16'b1111111111101010;
        weights1[21548] <= 16'b1111111111011011;
        weights1[21549] <= 16'b1111111111110111;
        weights1[21550] <= 16'b0000000000000000;
        weights1[21551] <= 16'b1111111111110110;
        weights1[21552] <= 16'b1111111111110101;
        weights1[21553] <= 16'b1111111111101111;
        weights1[21554] <= 16'b1111111111110001;
        weights1[21555] <= 16'b0000000000000101;
        weights1[21556] <= 16'b1111111111101100;
        weights1[21557] <= 16'b1111111111101001;
        weights1[21558] <= 16'b0000000000000000;
        weights1[21559] <= 16'b1111111111110001;
        weights1[21560] <= 16'b1111111111011011;
        weights1[21561] <= 16'b1111111111010101;
        weights1[21562] <= 16'b1111111111010011;
        weights1[21563] <= 16'b1111111111011111;
        weights1[21564] <= 16'b1111111111010111;
        weights1[21565] <= 16'b1111111111101110;
        weights1[21566] <= 16'b0000000000001101;
        weights1[21567] <= 16'b0000000000010100;
        weights1[21568] <= 16'b0000000000000001;
        weights1[21569] <= 16'b0000000000100100;
        weights1[21570] <= 16'b0000000000001101;
        weights1[21571] <= 16'b0000000000001100;
        weights1[21572] <= 16'b1111111111111000;
        weights1[21573] <= 16'b1111111111101110;
        weights1[21574] <= 16'b1111111111101000;
        weights1[21575] <= 16'b1111111111101110;
        weights1[21576] <= 16'b1111111111011111;
        weights1[21577] <= 16'b1111111111110101;
        weights1[21578] <= 16'b1111111111110011;
        weights1[21579] <= 16'b1111111111111010;
        weights1[21580] <= 16'b1111111111110101;
        weights1[21581] <= 16'b0000000000001101;
        weights1[21582] <= 16'b0000000000001101;
        weights1[21583] <= 16'b0000000000001001;
        weights1[21584] <= 16'b0000000000010000;
        weights1[21585] <= 16'b1111111111111101;
        weights1[21586] <= 16'b1111111111110001;
        weights1[21587] <= 16'b1111111111110010;
        weights1[21588] <= 16'b1111111111011100;
        weights1[21589] <= 16'b1111111110111011;
        weights1[21590] <= 16'b1111111110110110;
        weights1[21591] <= 16'b1111111110010100;
        weights1[21592] <= 16'b1111111110010000;
        weights1[21593] <= 16'b1111111101101110;
        weights1[21594] <= 16'b1111111110100010;
        weights1[21595] <= 16'b1111111111010011;
        weights1[21596] <= 16'b1111111111101111;
        weights1[21597] <= 16'b0000000000000110;
        weights1[21598] <= 16'b0000000000011100;
        weights1[21599] <= 16'b1111111111101001;
        weights1[21600] <= 16'b1111111111100100;
        weights1[21601] <= 16'b1111111111001110;
        weights1[21602] <= 16'b1111111111001011;
        weights1[21603] <= 16'b1111111111011010;
        weights1[21604] <= 16'b1111111111110010;
        weights1[21605] <= 16'b1111111111101010;
        weights1[21606] <= 16'b1111111111110000;
        weights1[21607] <= 16'b0000000000001010;
        weights1[21608] <= 16'b1111111111110100;
        weights1[21609] <= 16'b1111111111111000;
        weights1[21610] <= 16'b1111111111110111;
        weights1[21611] <= 16'b1111111111100110;
        weights1[21612] <= 16'b0000000000001011;
        weights1[21613] <= 16'b1111111111111110;
        weights1[21614] <= 16'b1111111111111100;
        weights1[21615] <= 16'b1111111111110111;
        weights1[21616] <= 16'b1111111111010000;
        weights1[21617] <= 16'b1111111110110111;
        weights1[21618] <= 16'b1111111110010110;
        weights1[21619] <= 16'b1111111101110010;
        weights1[21620] <= 16'b1111111101001101;
        weights1[21621] <= 16'b1111111100100101;
        weights1[21622] <= 16'b1111111100100001;
        weights1[21623] <= 16'b1111111100011100;
        weights1[21624] <= 16'b1111111100001101;
        weights1[21625] <= 16'b1111111101010111;
        weights1[21626] <= 16'b1111111101010101;
        weights1[21627] <= 16'b1111111101111101;
        weights1[21628] <= 16'b1111111110010101;
        weights1[21629] <= 16'b1111111110101011;
        weights1[21630] <= 16'b1111111111000110;
        weights1[21631] <= 16'b1111111111100111;
        weights1[21632] <= 16'b1111111111100111;
        weights1[21633] <= 16'b1111111111101010;
        weights1[21634] <= 16'b1111111111100110;
        weights1[21635] <= 16'b0000000000001001;
        weights1[21636] <= 16'b1111111111111101;
        weights1[21637] <= 16'b0000000000001010;
        weights1[21638] <= 16'b1111111111110100;
        weights1[21639] <= 16'b0000000000000001;
        weights1[21640] <= 16'b0000000000000010;
        weights1[21641] <= 16'b0000000000001001;
        weights1[21642] <= 16'b1111111111111100;
        weights1[21643] <= 16'b1111111111111001;
        weights1[21644] <= 16'b1111111111011100;
        weights1[21645] <= 16'b1111111110111000;
        weights1[21646] <= 16'b1111111110101011;
        weights1[21647] <= 16'b1111111110100111;
        weights1[21648] <= 16'b1111111101111101;
        weights1[21649] <= 16'b1111111101011111;
        weights1[21650] <= 16'b1111111101100100;
        weights1[21651] <= 16'b1111111100110000;
        weights1[21652] <= 16'b1111111100101100;
        weights1[21653] <= 16'b1111111100011111;
        weights1[21654] <= 16'b1111111101011110;
        weights1[21655] <= 16'b1111111110000100;
        weights1[21656] <= 16'b1111111110110010;
        weights1[21657] <= 16'b1111111111001110;
        weights1[21658] <= 16'b1111111111100101;
        weights1[21659] <= 16'b1111111111101010;
        weights1[21660] <= 16'b1111111111110100;
        weights1[21661] <= 16'b0000000000001001;
        weights1[21662] <= 16'b1111111111111010;
        weights1[21663] <= 16'b0000000000000110;
        weights1[21664] <= 16'b1111111111111000;
        weights1[21665] <= 16'b0000000000001011;
        weights1[21666] <= 16'b0000000000000110;
        weights1[21667] <= 16'b0000000000000100;
        weights1[21668] <= 16'b1111111111110100;
        weights1[21669] <= 16'b0000000000000011;
        weights1[21670] <= 16'b0000000000001001;
        weights1[21671] <= 16'b1111111111110111;
        weights1[21672] <= 16'b1111111111110011;
        weights1[21673] <= 16'b1111111111011001;
        weights1[21674] <= 16'b1111111111011111;
        weights1[21675] <= 16'b1111111111100110;
        weights1[21676] <= 16'b1111111111100000;
        weights1[21677] <= 16'b1111111111100000;
        weights1[21678] <= 16'b1111111111100010;
        weights1[21679] <= 16'b1111111111000101;
        weights1[21680] <= 16'b1111111111100100;
        weights1[21681] <= 16'b0000000000010001;
        weights1[21682] <= 16'b0000000000001111;
        weights1[21683] <= 16'b1111111111111111;
        weights1[21684] <= 16'b0000000000011001;
        weights1[21685] <= 16'b0000000000010001;
        weights1[21686] <= 16'b1111111111111111;
        weights1[21687] <= 16'b0000000000001100;
        weights1[21688] <= 16'b0000000000001100;
        weights1[21689] <= 16'b1111111111111110;
        weights1[21690] <= 16'b0000000000000111;
        weights1[21691] <= 16'b0000000000010010;
        weights1[21692] <= 16'b0000000000001110;
        weights1[21693] <= 16'b0000000000010111;
        weights1[21694] <= 16'b0000000000001100;
        weights1[21695] <= 16'b0000000000001111;
        weights1[21696] <= 16'b0000000000000100;
        weights1[21697] <= 16'b1111111111110111;
        weights1[21698] <= 16'b1111111111111011;
        weights1[21699] <= 16'b0000000000000101;
        weights1[21700] <= 16'b0000000000000010;
        weights1[21701] <= 16'b1111111111111010;
        weights1[21702] <= 16'b0000000000000011;
        weights1[21703] <= 16'b0000000000101000;
        weights1[21704] <= 16'b0000000000010100;
        weights1[21705] <= 16'b0000000000110101;
        weights1[21706] <= 16'b0000000000110101;
        weights1[21707] <= 16'b0000000001000111;
        weights1[21708] <= 16'b0000000001001110;
        weights1[21709] <= 16'b0000000000111111;
        weights1[21710] <= 16'b0000000000101010;
        weights1[21711] <= 16'b0000000000101011;
        weights1[21712] <= 16'b0000000000110001;
        weights1[21713] <= 16'b0000000000011011;
        weights1[21714] <= 16'b0000000000011001;
        weights1[21715] <= 16'b0000000000000010;
        weights1[21716] <= 16'b0000000000000011;
        weights1[21717] <= 16'b0000000000010101;
        weights1[21718] <= 16'b0000000000001100;
        weights1[21719] <= 16'b0000000000000010;
        weights1[21720] <= 16'b0000000000001010;
        weights1[21721] <= 16'b0000000000010000;
        weights1[21722] <= 16'b0000000000010000;
        weights1[21723] <= 16'b0000000000000100;
        weights1[21724] <= 16'b1111111111111111;
        weights1[21725] <= 16'b0000000000000111;
        weights1[21726] <= 16'b0000000000001001;
        weights1[21727] <= 16'b0000000000000101;
        weights1[21728] <= 16'b0000000000010010;
        weights1[21729] <= 16'b0000000000010100;
        weights1[21730] <= 16'b0000000000000111;
        weights1[21731] <= 16'b0000000001000101;
        weights1[21732] <= 16'b0000000001000011;
        weights1[21733] <= 16'b0000000000110101;
        weights1[21734] <= 16'b0000000000101101;
        weights1[21735] <= 16'b0000000000111011;
        weights1[21736] <= 16'b0000000001001000;
        weights1[21737] <= 16'b0000000000100101;
        weights1[21738] <= 16'b0000000000001101;
        weights1[21739] <= 16'b0000000000100000;
        weights1[21740] <= 16'b0000000000001111;
        weights1[21741] <= 16'b0000000000001010;
        weights1[21742] <= 16'b0000000000010100;
        weights1[21743] <= 16'b0000000000010011;
        weights1[21744] <= 16'b1111111111111101;
        weights1[21745] <= 16'b0000000000001101;
        weights1[21746] <= 16'b1111111111110001;
        weights1[21747] <= 16'b1111111111111100;
        weights1[21748] <= 16'b0000000000011001;
        weights1[21749] <= 16'b1111111111111010;
        weights1[21750] <= 16'b1111111111111110;
        weights1[21751] <= 16'b1111111111111110;
        weights1[21752] <= 16'b0000000000001000;
        weights1[21753] <= 16'b0000000000001110;
        weights1[21754] <= 16'b0000000000001101;
        weights1[21755] <= 16'b0000000000001110;
        weights1[21756] <= 16'b0000000000010100;
        weights1[21757] <= 16'b0000000000011011;
        weights1[21758] <= 16'b0000000000100011;
        weights1[21759] <= 16'b0000000000100011;
        weights1[21760] <= 16'b0000000000110001;
        weights1[21761] <= 16'b0000000000100010;
        weights1[21762] <= 16'b0000000000001111;
        weights1[21763] <= 16'b0000000000100110;
        weights1[21764] <= 16'b0000000000001001;
        weights1[21765] <= 16'b0000000000010010;
        weights1[21766] <= 16'b0000000000010001;
        weights1[21767] <= 16'b0000000000010001;
        weights1[21768] <= 16'b1111111111110100;
        weights1[21769] <= 16'b0000000000011100;
        weights1[21770] <= 16'b0000000000000011;
        weights1[21771] <= 16'b0000000000000011;
        weights1[21772] <= 16'b0000000000010001;
        weights1[21773] <= 16'b1111111111110111;
        weights1[21774] <= 16'b0000000000001111;
        weights1[21775] <= 16'b1111111111111100;
        weights1[21776] <= 16'b0000000000000101;
        weights1[21777] <= 16'b1111111111111010;
        weights1[21778] <= 16'b0000000000010111;
        weights1[21779] <= 16'b1111111111111111;
        weights1[21780] <= 16'b0000000000011101;
        weights1[21781] <= 16'b0000000000001101;
        weights1[21782] <= 16'b0000000000010110;
        weights1[21783] <= 16'b0000000000010100;
        weights1[21784] <= 16'b0000000000000110;
        weights1[21785] <= 16'b0000000000010000;
        weights1[21786] <= 16'b0000000000010010;
        weights1[21787] <= 16'b0000000000011011;
        weights1[21788] <= 16'b0000000000100011;
        weights1[21789] <= 16'b1111111111111101;
        weights1[21790] <= 16'b0000000000010011;
        weights1[21791] <= 16'b0000000000010101;
        weights1[21792] <= 16'b0000000000010111;
        weights1[21793] <= 16'b0000000000010101;
        weights1[21794] <= 16'b0000000000000101;
        weights1[21795] <= 16'b0000000000001010;
        weights1[21796] <= 16'b0000000000010111;
        weights1[21797] <= 16'b1111111111111101;
        weights1[21798] <= 16'b1111111111111100;
        weights1[21799] <= 16'b1111111111111110;
        weights1[21800] <= 16'b0000000000001100;
        weights1[21801] <= 16'b0000000000001101;
        weights1[21802] <= 16'b0000000000000000;
        weights1[21803] <= 16'b0000000000101010;
        weights1[21804] <= 16'b0000000000000111;
        weights1[21805] <= 16'b1111111111111000;
        weights1[21806] <= 16'b1111111111111110;
        weights1[21807] <= 16'b0000000000010011;
        weights1[21808] <= 16'b1111111111110010;
        weights1[21809] <= 16'b0000000000001010;
        weights1[21810] <= 16'b0000000000010100;
        weights1[21811] <= 16'b0000000000001101;
        weights1[21812] <= 16'b0000000000000101;
        weights1[21813] <= 16'b0000000000000111;
        weights1[21814] <= 16'b0000000000010010;
        weights1[21815] <= 16'b0000000000011000;
        weights1[21816] <= 16'b0000000000001011;
        weights1[21817] <= 16'b0000000000100101;
        weights1[21818] <= 16'b0000000000000101;
        weights1[21819] <= 16'b0000000000010111;
        weights1[21820] <= 16'b1111111111111101;
        weights1[21821] <= 16'b0000000000100100;
        weights1[21822] <= 16'b0000000000001000;
        weights1[21823] <= 16'b0000000000000111;
        weights1[21824] <= 16'b0000000000001011;
        weights1[21825] <= 16'b0000000000000110;
        weights1[21826] <= 16'b0000000000001100;
        weights1[21827] <= 16'b0000000000001100;
        weights1[21828] <= 16'b0000000000000100;
        weights1[21829] <= 16'b1111111111111101;
        weights1[21830] <= 16'b1111111111110110;
        weights1[21831] <= 16'b1111111111110101;
        weights1[21832] <= 16'b0000000000000001;
        weights1[21833] <= 16'b0000000000000011;
        weights1[21834] <= 16'b1111111111110111;
        weights1[21835] <= 16'b1111111111111111;
        weights1[21836] <= 16'b0000000000001000;
        weights1[21837] <= 16'b0000000000001110;
        weights1[21838] <= 16'b0000000000011010;
        weights1[21839] <= 16'b0000000000001111;
        weights1[21840] <= 16'b0000000000000011;
        weights1[21841] <= 16'b0000000000000010;
        weights1[21842] <= 16'b1111111111111101;
        weights1[21843] <= 16'b0000000000010011;
        weights1[21844] <= 16'b0000000000001010;
        weights1[21845] <= 16'b1111111111111101;
        weights1[21846] <= 16'b0000000000010111;
        weights1[21847] <= 16'b1111111111101010;
        weights1[21848] <= 16'b1111111111111010;
        weights1[21849] <= 16'b1111111111101111;
        weights1[21850] <= 16'b1111111111111000;
        weights1[21851] <= 16'b0000000000000011;
        weights1[21852] <= 16'b1111111111111010;
        weights1[21853] <= 16'b0000000000010000;
        weights1[21854] <= 16'b1111111111111000;
        weights1[21855] <= 16'b1111111111101011;
        weights1[21856] <= 16'b1111111111110100;
        weights1[21857] <= 16'b1111111111110001;
        weights1[21858] <= 16'b1111111111110110;
        weights1[21859] <= 16'b0000000000000110;
        weights1[21860] <= 16'b0000000000000101;
        weights1[21861] <= 16'b1111111111111001;
        weights1[21862] <= 16'b0000000000001101;
        weights1[21863] <= 16'b0000000000001110;
        weights1[21864] <= 16'b1111111111111101;
        weights1[21865] <= 16'b0000000000001001;
        weights1[21866] <= 16'b0000000000010110;
        weights1[21867] <= 16'b0000000000001000;
        weights1[21868] <= 16'b0000000000000100;
        weights1[21869] <= 16'b0000000000001010;
        weights1[21870] <= 16'b1111111111111100;
        weights1[21871] <= 16'b1111111111110110;
        weights1[21872] <= 16'b1111111111111011;
        weights1[21873] <= 16'b1111111111101110;
        weights1[21874] <= 16'b1111111111111000;
        weights1[21875] <= 16'b1111111111110110;
        weights1[21876] <= 16'b1111111111111010;
        weights1[21877] <= 16'b1111111111101001;
        weights1[21878] <= 16'b0000000000010010;
        weights1[21879] <= 16'b0000000000010011;
        weights1[21880] <= 16'b1111111111110111;
        weights1[21881] <= 16'b1111111111101011;
        weights1[21882] <= 16'b0000000000000101;
        weights1[21883] <= 16'b1111111111111101;
        weights1[21884] <= 16'b0000000000000011;
        weights1[21885] <= 16'b1111111111111110;
        weights1[21886] <= 16'b0000000000001110;
        weights1[21887] <= 16'b0000000000000011;
        weights1[21888] <= 16'b1111111111111101;
        weights1[21889] <= 16'b0000000000001010;
        weights1[21890] <= 16'b1111111111110100;
        weights1[21891] <= 16'b1111111111111000;
        weights1[21892] <= 16'b0000000000001011;
        weights1[21893] <= 16'b0000000000001000;
        weights1[21894] <= 16'b0000000000000000;
        weights1[21895] <= 16'b0000000000000111;
        weights1[21896] <= 16'b0000000000000111;
        weights1[21897] <= 16'b0000000000001001;
        weights1[21898] <= 16'b0000000000000011;
        weights1[21899] <= 16'b1111111111111010;
        weights1[21900] <= 16'b1111111111111000;
        weights1[21901] <= 16'b1111111111100101;
        weights1[21902] <= 16'b1111111111110100;
        weights1[21903] <= 16'b1111111111101001;
        weights1[21904] <= 16'b1111111111111100;
        weights1[21905] <= 16'b1111111111110011;
        weights1[21906] <= 16'b1111111111110000;
        weights1[21907] <= 16'b1111111111111101;
        weights1[21908] <= 16'b1111111111101101;
        weights1[21909] <= 16'b0000000000001100;
        weights1[21910] <= 16'b1111111111111110;
        weights1[21911] <= 16'b0000000000001001;
        weights1[21912] <= 16'b1111111111111110;
        weights1[21913] <= 16'b0000000000000110;
        weights1[21914] <= 16'b0000000000000111;
        weights1[21915] <= 16'b0000000000000110;
        weights1[21916] <= 16'b0000000000001010;
        weights1[21917] <= 16'b0000000000011000;
        weights1[21918] <= 16'b0000000000001111;
        weights1[21919] <= 16'b1111111111111001;
        weights1[21920] <= 16'b0000000000000101;
        weights1[21921] <= 16'b0000000000001000;
        weights1[21922] <= 16'b0000000000000100;
        weights1[21923] <= 16'b0000000000000001;
        weights1[21924] <= 16'b0000000000000010;
        weights1[21925] <= 16'b0000000000001010;
        weights1[21926] <= 16'b0000000000001011;
        weights1[21927] <= 16'b0000000000001000;
        weights1[21928] <= 16'b0000000000000111;
        weights1[21929] <= 16'b1111111111111111;
        weights1[21930] <= 16'b0000000000001101;
        weights1[21931] <= 16'b1111111111111111;
        weights1[21932] <= 16'b0000000000000110;
        weights1[21933] <= 16'b0000000000000100;
        weights1[21934] <= 16'b0000000000000111;
        weights1[21935] <= 16'b0000000000001110;
        weights1[21936] <= 16'b0000000000010010;
        weights1[21937] <= 16'b0000000000100011;
        weights1[21938] <= 16'b0000000000011001;
        weights1[21939] <= 16'b0000000000011000;
        weights1[21940] <= 16'b0000000000001101;
        weights1[21941] <= 16'b0000000000010100;
        weights1[21942] <= 16'b0000000000000011;
        weights1[21943] <= 16'b0000000000001101;
        weights1[21944] <= 16'b0000000000001110;
        weights1[21945] <= 16'b0000000000010001;
        weights1[21946] <= 16'b1111111111111110;
        weights1[21947] <= 16'b0000000000000000;
        weights1[21948] <= 16'b1111111111111001;
        weights1[21949] <= 16'b0000000000000011;
        weights1[21950] <= 16'b0000000000000101;
        weights1[21951] <= 16'b0000000000000000;
        weights1[21952] <= 16'b0000000000000000;
        weights1[21953] <= 16'b0000000000000000;
        weights1[21954] <= 16'b0000000000000000;
        weights1[21955] <= 16'b0000000000000000;
        weights1[21956] <= 16'b0000000000000000;
        weights1[21957] <= 16'b0000000000000000;
        weights1[21958] <= 16'b1111111111111011;
        weights1[21959] <= 16'b1111111111111100;
        weights1[21960] <= 16'b1111111111111010;
        weights1[21961] <= 16'b1111111111111010;
        weights1[21962] <= 16'b1111111111111100;
        weights1[21963] <= 16'b1111111111110101;
        weights1[21964] <= 16'b1111111111110000;
        weights1[21965] <= 16'b1111111111101111;
        weights1[21966] <= 16'b1111111111101100;
        weights1[21967] <= 16'b1111111111110101;
        weights1[21968] <= 16'b1111111111101000;
        weights1[21969] <= 16'b1111111111101010;
        weights1[21970] <= 16'b1111111111110110;
        weights1[21971] <= 16'b1111111111111010;
        weights1[21972] <= 16'b1111111111111001;
        weights1[21973] <= 16'b1111111111111000;
        weights1[21974] <= 16'b0000000000000000;
        weights1[21975] <= 16'b0000000000000011;
        weights1[21976] <= 16'b0000000000000100;
        weights1[21977] <= 16'b0000000000000110;
        weights1[21978] <= 16'b0000000000000001;
        weights1[21979] <= 16'b1111111111111111;
        weights1[21980] <= 16'b0000000000000000;
        weights1[21981] <= 16'b0000000000000000;
        weights1[21982] <= 16'b0000000000000001;
        weights1[21983] <= 16'b0000000000000001;
        weights1[21984] <= 16'b1111111111111100;
        weights1[21985] <= 16'b0000000000000010;
        weights1[21986] <= 16'b0000000000000000;
        weights1[21987] <= 16'b0000000000000001;
        weights1[21988] <= 16'b0000000000000000;
        weights1[21989] <= 16'b1111111111111111;
        weights1[21990] <= 16'b1111111111111011;
        weights1[21991] <= 16'b1111111111101111;
        weights1[21992] <= 16'b1111111111101100;
        weights1[21993] <= 16'b1111111111101100;
        weights1[21994] <= 16'b1111111111100011;
        weights1[21995] <= 16'b1111111111100110;
        weights1[21996] <= 16'b1111111111100100;
        weights1[21997] <= 16'b1111111111010101;
        weights1[21998] <= 16'b1111111111100101;
        weights1[21999] <= 16'b1111111111100011;
        weights1[22000] <= 16'b1111111111101001;
        weights1[22001] <= 16'b1111111111101111;
        weights1[22002] <= 16'b1111111111111000;
        weights1[22003] <= 16'b1111111111111010;
        weights1[22004] <= 16'b1111111111111100;
        weights1[22005] <= 16'b0000000000000000;
        weights1[22006] <= 16'b0000000000000011;
        weights1[22007] <= 16'b0000000000000011;
        weights1[22008] <= 16'b0000000000000000;
        weights1[22009] <= 16'b0000000000000000;
        weights1[22010] <= 16'b0000000000000000;
        weights1[22011] <= 16'b1111111111111101;
        weights1[22012] <= 16'b1111111111111011;
        weights1[22013] <= 16'b1111111111111101;
        weights1[22014] <= 16'b1111111111111011;
        weights1[22015] <= 16'b0000000000000100;
        weights1[22016] <= 16'b1111111111111111;
        weights1[22017] <= 16'b0000000000000001;
        weights1[22018] <= 16'b1111111111110101;
        weights1[22019] <= 16'b1111111111101101;
        weights1[22020] <= 16'b1111111111010010;
        weights1[22021] <= 16'b1111111111011011;
        weights1[22022] <= 16'b1111111111110011;
        weights1[22023] <= 16'b1111111111101001;
        weights1[22024] <= 16'b1111111111101010;
        weights1[22025] <= 16'b1111111111100011;
        weights1[22026] <= 16'b0000000000000011;
        weights1[22027] <= 16'b0000000000000010;
        weights1[22028] <= 16'b1111111111101100;
        weights1[22029] <= 16'b1111111111111111;
        weights1[22030] <= 16'b1111111111101100;
        weights1[22031] <= 16'b1111111111111100;
        weights1[22032] <= 16'b1111111111110100;
        weights1[22033] <= 16'b0000000000000110;
        weights1[22034] <= 16'b0000000000000011;
        weights1[22035] <= 16'b0000000000000101;
        weights1[22036] <= 16'b0000000000000000;
        weights1[22037] <= 16'b0000000000000000;
        weights1[22038] <= 16'b1111111111111101;
        weights1[22039] <= 16'b1111111111111101;
        weights1[22040] <= 16'b1111111111111010;
        weights1[22041] <= 16'b1111111111110111;
        weights1[22042] <= 16'b1111111111111101;
        weights1[22043] <= 16'b1111111111110111;
        weights1[22044] <= 16'b1111111111110001;
        weights1[22045] <= 16'b1111111111101011;
        weights1[22046] <= 16'b1111111111011000;
        weights1[22047] <= 16'b1111111111011110;
        weights1[22048] <= 16'b1111111111001011;
        weights1[22049] <= 16'b1111111111110010;
        weights1[22050] <= 16'b1111111111010101;
        weights1[22051] <= 16'b1111111111100010;
        weights1[22052] <= 16'b1111111111101111;
        weights1[22053] <= 16'b0000000000001001;
        weights1[22054] <= 16'b0000000000000110;
        weights1[22055] <= 16'b1111111111111110;
        weights1[22056] <= 16'b1111111111110100;
        weights1[22057] <= 16'b1111111111111110;
        weights1[22058] <= 16'b0000000000000110;
        weights1[22059] <= 16'b1111111111111110;
        weights1[22060] <= 16'b1111111111111000;
        weights1[22061] <= 16'b1111111111110011;
        weights1[22062] <= 16'b1111111111110101;
        weights1[22063] <= 16'b0000000000000001;
        weights1[22064] <= 16'b1111111111111110;
        weights1[22065] <= 16'b0000000000000000;
        weights1[22066] <= 16'b1111111111111110;
        weights1[22067] <= 16'b1111111111111101;
        weights1[22068] <= 16'b1111111111111101;
        weights1[22069] <= 16'b1111111111110100;
        weights1[22070] <= 16'b1111111111100000;
        weights1[22071] <= 16'b1111111111011111;
        weights1[22072] <= 16'b1111111111011111;
        weights1[22073] <= 16'b1111111111111011;
        weights1[22074] <= 16'b1111111111110111;
        weights1[22075] <= 16'b1111111111111101;
        weights1[22076] <= 16'b1111111111110000;
        weights1[22077] <= 16'b0000000000000100;
        weights1[22078] <= 16'b1111111111101110;
        weights1[22079] <= 16'b1111111111101000;
        weights1[22080] <= 16'b1111111111110110;
        weights1[22081] <= 16'b1111111111111001;
        weights1[22082] <= 16'b1111111111101111;
        weights1[22083] <= 16'b1111111111111000;
        weights1[22084] <= 16'b1111111111100010;
        weights1[22085] <= 16'b0000000000000111;
        weights1[22086] <= 16'b1111111111110000;
        weights1[22087] <= 16'b0000000000000000;
        weights1[22088] <= 16'b1111111111111000;
        weights1[22089] <= 16'b0000000000001010;
        weights1[22090] <= 16'b1111111111111001;
        weights1[22091] <= 16'b1111111111111100;
        weights1[22092] <= 16'b1111111111111110;
        weights1[22093] <= 16'b1111111111111100;
        weights1[22094] <= 16'b1111111111111100;
        weights1[22095] <= 16'b1111111111111000;
        weights1[22096] <= 16'b1111111111111111;
        weights1[22097] <= 16'b0000000000010010;
        weights1[22098] <= 16'b1111111111110110;
        weights1[22099] <= 16'b1111111111011011;
        weights1[22100] <= 16'b1111111111100111;
        weights1[22101] <= 16'b0000000000000110;
        weights1[22102] <= 16'b1111111111110001;
        weights1[22103] <= 16'b0000000000001001;
        weights1[22104] <= 16'b1111111111110001;
        weights1[22105] <= 16'b1111111111101011;
        weights1[22106] <= 16'b1111111111111000;
        weights1[22107] <= 16'b0000000000000011;
        weights1[22108] <= 16'b0000000000000010;
        weights1[22109] <= 16'b0000000000001100;
        weights1[22110] <= 16'b1111111111101111;
        weights1[22111] <= 16'b0000000000001010;
        weights1[22112] <= 16'b0000000000000001;
        weights1[22113] <= 16'b1111111111111110;
        weights1[22114] <= 16'b1111111111111111;
        weights1[22115] <= 16'b1111111111111010;
        weights1[22116] <= 16'b0000000000000110;
        weights1[22117] <= 16'b0000000000000011;
        weights1[22118] <= 16'b0000000000001001;
        weights1[22119] <= 16'b0000000000000011;
        weights1[22120] <= 16'b1111111111111100;
        weights1[22121] <= 16'b1111111111110110;
        weights1[22122] <= 16'b1111111111101111;
        weights1[22123] <= 16'b1111111111110111;
        weights1[22124] <= 16'b0000000000000000;
        weights1[22125] <= 16'b0000000000001101;
        weights1[22126] <= 16'b1111111111110110;
        weights1[22127] <= 16'b1111111111101101;
        weights1[22128] <= 16'b1111111111100011;
        weights1[22129] <= 16'b1111111111100100;
        weights1[22130] <= 16'b1111111111110111;
        weights1[22131] <= 16'b0000000000000001;
        weights1[22132] <= 16'b0000000000000101;
        weights1[22133] <= 16'b1111111111110011;
        weights1[22134] <= 16'b0000000000000000;
        weights1[22135] <= 16'b1111111111110111;
        weights1[22136] <= 16'b1111111111111110;
        weights1[22137] <= 16'b0000000000000111;
        weights1[22138] <= 16'b0000000000001101;
        weights1[22139] <= 16'b0000000000010000;
        weights1[22140] <= 16'b0000000000011100;
        weights1[22141] <= 16'b0000000000001110;
        weights1[22142] <= 16'b0000000000000111;
        weights1[22143] <= 16'b0000000000000100;
        weights1[22144] <= 16'b0000000000101111;
        weights1[22145] <= 16'b0000000000010111;
        weights1[22146] <= 16'b0000000000010101;
        weights1[22147] <= 16'b0000000000010001;
        weights1[22148] <= 16'b1111111111111100;
        weights1[22149] <= 16'b1111111111110111;
        weights1[22150] <= 16'b1111111111101111;
        weights1[22151] <= 16'b1111111111110110;
        weights1[22152] <= 16'b1111111111111001;
        weights1[22153] <= 16'b1111111111100011;
        weights1[22154] <= 16'b0000000000000011;
        weights1[22155] <= 16'b1111111111101101;
        weights1[22156] <= 16'b1111111111111100;
        weights1[22157] <= 16'b1111111111111011;
        weights1[22158] <= 16'b1111111111110110;
        weights1[22159] <= 16'b1111111111111000;
        weights1[22160] <= 16'b1111111111111110;
        weights1[22161] <= 16'b0000000000010000;
        weights1[22162] <= 16'b1111111111110010;
        weights1[22163] <= 16'b0000000000001000;
        weights1[22164] <= 16'b1111111111110100;
        weights1[22165] <= 16'b0000000000001110;
        weights1[22166] <= 16'b0000000000000010;
        weights1[22167] <= 16'b1111111111110011;
        weights1[22168] <= 16'b0000000000001101;
        weights1[22169] <= 16'b0000000000100101;
        weights1[22170] <= 16'b0000000000101110;
        weights1[22171] <= 16'b0000000000011011;
        weights1[22172] <= 16'b1111111111111100;
        weights1[22173] <= 16'b0000000000011001;
        weights1[22174] <= 16'b0000000000011000;
        weights1[22175] <= 16'b0000000000011110;
        weights1[22176] <= 16'b1111111111111010;
        weights1[22177] <= 16'b1111111111110101;
        weights1[22178] <= 16'b1111111111110101;
        weights1[22179] <= 16'b1111111111111000;
        weights1[22180] <= 16'b1111111111110010;
        weights1[22181] <= 16'b1111111111101011;
        weights1[22182] <= 16'b0000000000000001;
        weights1[22183] <= 16'b1111111111011101;
        weights1[22184] <= 16'b0000000000000010;
        weights1[22185] <= 16'b1111111111110001;
        weights1[22186] <= 16'b0000000000001001;
        weights1[22187] <= 16'b1111111111111110;
        weights1[22188] <= 16'b1111111111111001;
        weights1[22189] <= 16'b1111111111110101;
        weights1[22190] <= 16'b0000000000001000;
        weights1[22191] <= 16'b0000000000010101;
        weights1[22192] <= 16'b0000000000011011;
        weights1[22193] <= 16'b0000000000000001;
        weights1[22194] <= 16'b0000000000010010;
        weights1[22195] <= 16'b0000000000000100;
        weights1[22196] <= 16'b0000000000010010;
        weights1[22197] <= 16'b0000000000011110;
        weights1[22198] <= 16'b0000000000010111;
        weights1[22199] <= 16'b0000000000010110;
        weights1[22200] <= 16'b0000000000110110;
        weights1[22201] <= 16'b0000000000101010;
        weights1[22202] <= 16'b0000000000011110;
        weights1[22203] <= 16'b0000000000110101;
        weights1[22204] <= 16'b1111111111110101;
        weights1[22205] <= 16'b1111111111111101;
        weights1[22206] <= 16'b1111111111111001;
        weights1[22207] <= 16'b1111111111110100;
        weights1[22208] <= 16'b1111111111111111;
        weights1[22209] <= 16'b1111111111110101;
        weights1[22210] <= 16'b1111111111101110;
        weights1[22211] <= 16'b1111111111011111;
        weights1[22212] <= 16'b0000000000000011;
        weights1[22213] <= 16'b1111111111110010;
        weights1[22214] <= 16'b1111111111101110;
        weights1[22215] <= 16'b1111111111111010;
        weights1[22216] <= 16'b1111111111111111;
        weights1[22217] <= 16'b0000000000001000;
        weights1[22218] <= 16'b0000000000000101;
        weights1[22219] <= 16'b0000000000010100;
        weights1[22220] <= 16'b0000000000010000;
        weights1[22221] <= 16'b0000000000100010;
        weights1[22222] <= 16'b0000000000100110;
        weights1[22223] <= 16'b0000000000111001;
        weights1[22224] <= 16'b0000000000101100;
        weights1[22225] <= 16'b0000000000100100;
        weights1[22226] <= 16'b0000000000101110;
        weights1[22227] <= 16'b0000000000111000;
        weights1[22228] <= 16'b0000000001000001;
        weights1[22229] <= 16'b0000000000110101;
        weights1[22230] <= 16'b0000000000000101;
        weights1[22231] <= 16'b0000000000101100;
        weights1[22232] <= 16'b1111111111110010;
        weights1[22233] <= 16'b1111111111111100;
        weights1[22234] <= 16'b0000000000010101;
        weights1[22235] <= 16'b1111111111110100;
        weights1[22236] <= 16'b1111111111100110;
        weights1[22237] <= 16'b1111111111101110;
        weights1[22238] <= 16'b1111111111111000;
        weights1[22239] <= 16'b1111111111110101;
        weights1[22240] <= 16'b1111111111110101;
        weights1[22241] <= 16'b1111111111101000;
        weights1[22242] <= 16'b0000000000000000;
        weights1[22243] <= 16'b1111111111110100;
        weights1[22244] <= 16'b1111111111111000;
        weights1[22245] <= 16'b0000000000001000;
        weights1[22246] <= 16'b1111111111110110;
        weights1[22247] <= 16'b1111111111111011;
        weights1[22248] <= 16'b0000000000010010;
        weights1[22249] <= 16'b0000000000011100;
        weights1[22250] <= 16'b0000000000100111;
        weights1[22251] <= 16'b0000000000011000;
        weights1[22252] <= 16'b0000000000110011;
        weights1[22253] <= 16'b0000000000110000;
        weights1[22254] <= 16'b0000000000111000;
        weights1[22255] <= 16'b0000000001001111;
        weights1[22256] <= 16'b0000000000100110;
        weights1[22257] <= 16'b0000000001000011;
        weights1[22258] <= 16'b0000000000001101;
        weights1[22259] <= 16'b1111111111111100;
        weights1[22260] <= 16'b1111111111110001;
        weights1[22261] <= 16'b1111111111110000;
        weights1[22262] <= 16'b0000000000000011;
        weights1[22263] <= 16'b1111111111101110;
        weights1[22264] <= 16'b1111111111111110;
        weights1[22265] <= 16'b1111111111110111;
        weights1[22266] <= 16'b1111111111110011;
        weights1[22267] <= 16'b0000000000000101;
        weights1[22268] <= 16'b1111111111110110;
        weights1[22269] <= 16'b0000000000000111;
        weights1[22270] <= 16'b1111111111110100;
        weights1[22271] <= 16'b1111111111100111;
        weights1[22272] <= 16'b1111111111110100;
        weights1[22273] <= 16'b1111111111011100;
        weights1[22274] <= 16'b1111111111010001;
        weights1[22275] <= 16'b1111111111000011;
        weights1[22276] <= 16'b1111111110110111;
        weights1[22277] <= 16'b1111111111001100;
        weights1[22278] <= 16'b1111111111001001;
        weights1[22279] <= 16'b1111111111100001;
        weights1[22280] <= 16'b1111111111100110;
        weights1[22281] <= 16'b0000000000011111;
        weights1[22282] <= 16'b0000000000010100;
        weights1[22283] <= 16'b0000000000000010;
        weights1[22284] <= 16'b1111111111110110;
        weights1[22285] <= 16'b1111111111111100;
        weights1[22286] <= 16'b1111111111101001;
        weights1[22287] <= 16'b1111111111101100;
        weights1[22288] <= 16'b1111111111111100;
        weights1[22289] <= 16'b1111111111110001;
        weights1[22290] <= 16'b0000000000001000;
        weights1[22291] <= 16'b1111111111111101;
        weights1[22292] <= 16'b1111111111110001;
        weights1[22293] <= 16'b0000000000000010;
        weights1[22294] <= 16'b1111111111111101;
        weights1[22295] <= 16'b1111111111101010;
        weights1[22296] <= 16'b1111111111111001;
        weights1[22297] <= 16'b1111111111100000;
        weights1[22298] <= 16'b1111111111111000;
        weights1[22299] <= 16'b1111111111101110;
        weights1[22300] <= 16'b1111111111011100;
        weights1[22301] <= 16'b1111111111101100;
        weights1[22302] <= 16'b1111111111010001;
        weights1[22303] <= 16'b1111111110111101;
        weights1[22304] <= 16'b1111111101110101;
        weights1[22305] <= 16'b1111111101000110;
        weights1[22306] <= 16'b1111111100011110;
        weights1[22307] <= 16'b1111111100100010;
        weights1[22308] <= 16'b1111111100010110;
        weights1[22309] <= 16'b1111111101000010;
        weights1[22310] <= 16'b1111111101010010;
        weights1[22311] <= 16'b1111111101100001;
        weights1[22312] <= 16'b1111111110001110;
        weights1[22313] <= 16'b1111111110011010;
        weights1[22314] <= 16'b1111111110101111;
        weights1[22315] <= 16'b1111111110110010;
        weights1[22316] <= 16'b0000000000001000;
        weights1[22317] <= 16'b1111111111111010;
        weights1[22318] <= 16'b0000000000010000;
        weights1[22319] <= 16'b0000000000001101;
        weights1[22320] <= 16'b1111111111111101;
        weights1[22321] <= 16'b1111111111111110;
        weights1[22322] <= 16'b1111111111110000;
        weights1[22323] <= 16'b1111111111110111;
        weights1[22324] <= 16'b0000000000000100;
        weights1[22325] <= 16'b1111111111110010;
        weights1[22326] <= 16'b1111111111101101;
        weights1[22327] <= 16'b1111111111111010;
        weights1[22328] <= 16'b0000000000001111;
        weights1[22329] <= 16'b1111111111111100;
        weights1[22330] <= 16'b1111111111111101;
        weights1[22331] <= 16'b1111111111101011;
        weights1[22332] <= 16'b1111111111101011;
        weights1[22333] <= 16'b1111111111001111;
        weights1[22334] <= 16'b1111111110001001;
        weights1[22335] <= 16'b1111111100010000;
        weights1[22336] <= 16'b1111111100001111;
        weights1[22337] <= 16'b1111111100011001;
        weights1[22338] <= 16'b1111111100111000;
        weights1[22339] <= 16'b1111111101000000;
        weights1[22340] <= 16'b1111111101011101;
        weights1[22341] <= 16'b1111111110000100;
        weights1[22342] <= 16'b1111111110101100;
        weights1[22343] <= 16'b1111111110110001;
        weights1[22344] <= 16'b0000000000000101;
        weights1[22345] <= 16'b1111111111111110;
        weights1[22346] <= 16'b1111111111111111;
        weights1[22347] <= 16'b0000000000010001;
        weights1[22348] <= 16'b0000000000010010;
        weights1[22349] <= 16'b1111111111111001;
        weights1[22350] <= 16'b0000000000001000;
        weights1[22351] <= 16'b1111111111110101;
        weights1[22352] <= 16'b0000000000000011;
        weights1[22353] <= 16'b0000000000001100;
        weights1[22354] <= 16'b0000000000000010;
        weights1[22355] <= 16'b1111111111111110;
        weights1[22356] <= 16'b1111111111110011;
        weights1[22357] <= 16'b1111111111110101;
        weights1[22358] <= 16'b0000000000010010;
        weights1[22359] <= 16'b0000000000001010;
        weights1[22360] <= 16'b0000000000011101;
        weights1[22361] <= 16'b0000000000000111;
        weights1[22362] <= 16'b0000000000001010;
        weights1[22363] <= 16'b1111111111011111;
        weights1[22364] <= 16'b1111111110100110;
        weights1[22365] <= 16'b1111111101010111;
        weights1[22366] <= 16'b1111111101010010;
        weights1[22367] <= 16'b1111111101100101;
        weights1[22368] <= 16'b1111111101110100;
        weights1[22369] <= 16'b1111111110001101;
        weights1[22370] <= 16'b1111111110101001;
        weights1[22371] <= 16'b1111111110101000;
        weights1[22372] <= 16'b0000000000000101;
        weights1[22373] <= 16'b0000000000000011;
        weights1[22374] <= 16'b0000000000001001;
        weights1[22375] <= 16'b0000000000000010;
        weights1[22376] <= 16'b1111111111111001;
        weights1[22377] <= 16'b0000000000001011;
        weights1[22378] <= 16'b0000000000010111;
        weights1[22379] <= 16'b1111111111111110;
        weights1[22380] <= 16'b0000000000001011;
        weights1[22381] <= 16'b0000000000001010;
        weights1[22382] <= 16'b1111111111110100;
        weights1[22383] <= 16'b0000000000000001;
        weights1[22384] <= 16'b1111111111111011;
        weights1[22385] <= 16'b1111111111111001;
        weights1[22386] <= 16'b1111111111111111;
        weights1[22387] <= 16'b0000000000000001;
        weights1[22388] <= 16'b0000000000000100;
        weights1[22389] <= 16'b0000000000011110;
        weights1[22390] <= 16'b0000000000101100;
        weights1[22391] <= 16'b0000000000001000;
        weights1[22392] <= 16'b0000000000010010;
        weights1[22393] <= 16'b1111111111011111;
        weights1[22394] <= 16'b1111111110101000;
        weights1[22395] <= 16'b1111111110010101;
        weights1[22396] <= 16'b1111111101110010;
        weights1[22397] <= 16'b1111111110011001;
        weights1[22398] <= 16'b1111111110111100;
        weights1[22399] <= 16'b1111111110011101;
        weights1[22400] <= 16'b0000000000010000;
        weights1[22401] <= 16'b0000000000010110;
        weights1[22402] <= 16'b1111111111101111;
        weights1[22403] <= 16'b1111111111111001;
        weights1[22404] <= 16'b1111111111110111;
        weights1[22405] <= 16'b0000000000010000;
        weights1[22406] <= 16'b1111111111111111;
        weights1[22407] <= 16'b0000000000001001;
        weights1[22408] <= 16'b1111111111111011;
        weights1[22409] <= 16'b0000000000001100;
        weights1[22410] <= 16'b1111111111110111;
        weights1[22411] <= 16'b0000000000000000;
        weights1[22412] <= 16'b0000000000001000;
        weights1[22413] <= 16'b1111111111111011;
        weights1[22414] <= 16'b1111111111110110;
        weights1[22415] <= 16'b1111111111111101;
        weights1[22416] <= 16'b0000000000010000;
        weights1[22417] <= 16'b0000000000000010;
        weights1[22418] <= 16'b0000000000001100;
        weights1[22419] <= 16'b0000000000001111;
        weights1[22420] <= 16'b0000000000010100;
        weights1[22421] <= 16'b0000000000011100;
        weights1[22422] <= 16'b0000000000011110;
        weights1[22423] <= 16'b1111111111101011;
        weights1[22424] <= 16'b1111111110110100;
        weights1[22425] <= 16'b1111111110100111;
        weights1[22426] <= 16'b1111111110111110;
        weights1[22427] <= 16'b1111111110111011;
        weights1[22428] <= 16'b0000000000001101;
        weights1[22429] <= 16'b0000000000000101;
        weights1[22430] <= 16'b1111111111101111;
        weights1[22431] <= 16'b1111111111111000;
        weights1[22432] <= 16'b0000000000001001;
        weights1[22433] <= 16'b0000000000000100;
        weights1[22434] <= 16'b0000000000000001;
        weights1[22435] <= 16'b0000000000010001;
        weights1[22436] <= 16'b1111111111111110;
        weights1[22437] <= 16'b1111111111111000;
        weights1[22438] <= 16'b0000000000000111;
        weights1[22439] <= 16'b1111111111101001;
        weights1[22440] <= 16'b1111111111111111;
        weights1[22441] <= 16'b1111111111111100;
        weights1[22442] <= 16'b1111111111111101;
        weights1[22443] <= 16'b0000000000001101;
        weights1[22444] <= 16'b0000000000000111;
        weights1[22445] <= 16'b0000000000001010;
        weights1[22446] <= 16'b0000000000001000;
        weights1[22447] <= 16'b0000000000010111;
        weights1[22448] <= 16'b0000000000011110;
        weights1[22449] <= 16'b1111111111111000;
        weights1[22450] <= 16'b0000000000011100;
        weights1[22451] <= 16'b0000000000011011;
        weights1[22452] <= 16'b1111111111110110;
        weights1[22453] <= 16'b1111111111100111;
        weights1[22454] <= 16'b1111111111001110;
        weights1[22455] <= 16'b1111111111001010;
        weights1[22456] <= 16'b0000000000000001;
        weights1[22457] <= 16'b0000000000000101;
        weights1[22458] <= 16'b0000000000001100;
        weights1[22459] <= 16'b0000000000000110;
        weights1[22460] <= 16'b0000000000000010;
        weights1[22461] <= 16'b0000000000000101;
        weights1[22462] <= 16'b1111111111111111;
        weights1[22463] <= 16'b0000000000001111;
        weights1[22464] <= 16'b0000000000000000;
        weights1[22465] <= 16'b1111111111111011;
        weights1[22466] <= 16'b0000000000000111;
        weights1[22467] <= 16'b0000000000000011;
        weights1[22468] <= 16'b0000000000000000;
        weights1[22469] <= 16'b1111111111111001;
        weights1[22470] <= 16'b0000000000001000;
        weights1[22471] <= 16'b1111111111111110;
        weights1[22472] <= 16'b0000000000001100;
        weights1[22473] <= 16'b0000000000001000;
        weights1[22474] <= 16'b0000000000010011;
        weights1[22475] <= 16'b1111111111111111;
        weights1[22476] <= 16'b0000000000011110;
        weights1[22477] <= 16'b1111111111111110;
        weights1[22478] <= 16'b0000000000001000;
        weights1[22479] <= 16'b0000000000001000;
        weights1[22480] <= 16'b1111111111110101;
        weights1[22481] <= 16'b1111111111101001;
        weights1[22482] <= 16'b1111111111011011;
        weights1[22483] <= 16'b1111111111010001;
        weights1[22484] <= 16'b1111111111111101;
        weights1[22485] <= 16'b0000000000001010;
        weights1[22486] <= 16'b1111111111111111;
        weights1[22487] <= 16'b0000000000001001;
        weights1[22488] <= 16'b1111111111110100;
        weights1[22489] <= 16'b1111111111111011;
        weights1[22490] <= 16'b0000000000000111;
        weights1[22491] <= 16'b0000000000001111;
        weights1[22492] <= 16'b0000000000000101;
        weights1[22493] <= 16'b0000000000000011;
        weights1[22494] <= 16'b1111111111110101;
        weights1[22495] <= 16'b0000000000001110;
        weights1[22496] <= 16'b0000000000000011;
        weights1[22497] <= 16'b1111111111111100;
        weights1[22498] <= 16'b0000000000000001;
        weights1[22499] <= 16'b0000000000001011;
        weights1[22500] <= 16'b0000000000001100;
        weights1[22501] <= 16'b0000000000000101;
        weights1[22502] <= 16'b0000000000000010;
        weights1[22503] <= 16'b0000000000000101;
        weights1[22504] <= 16'b0000000000010110;
        weights1[22505] <= 16'b0000000000000101;
        weights1[22506] <= 16'b0000000000100000;
        weights1[22507] <= 16'b0000000000011000;
        weights1[22508] <= 16'b0000000000001110;
        weights1[22509] <= 16'b1111111111110100;
        weights1[22510] <= 16'b1111111111100101;
        weights1[22511] <= 16'b1111111111011111;
        weights1[22512] <= 16'b1111111111111010;
        weights1[22513] <= 16'b1111111111111001;
        weights1[22514] <= 16'b0000000000010010;
        weights1[22515] <= 16'b1111111111111101;
        weights1[22516] <= 16'b1111111111111110;
        weights1[22517] <= 16'b0000000000001010;
        weights1[22518] <= 16'b0000000000000000;
        weights1[22519] <= 16'b1111111111110111;
        weights1[22520] <= 16'b0000000000001010;
        weights1[22521] <= 16'b1111111111111000;
        weights1[22522] <= 16'b0000000000000110;
        weights1[22523] <= 16'b0000000000000101;
        weights1[22524] <= 16'b0000000000000101;
        weights1[22525] <= 16'b1111111111111010;
        weights1[22526] <= 16'b0000000000000100;
        weights1[22527] <= 16'b0000000000000110;
        weights1[22528] <= 16'b0000000000000101;
        weights1[22529] <= 16'b1111111111111011;
        weights1[22530] <= 16'b0000000000011101;
        weights1[22531] <= 16'b1111111111110110;
        weights1[22532] <= 16'b0000000000011000;
        weights1[22533] <= 16'b0000000000000111;
        weights1[22534] <= 16'b0000000000000001;
        weights1[22535] <= 16'b0000000000010010;
        weights1[22536] <= 16'b0000000000000100;
        weights1[22537] <= 16'b0000000000000111;
        weights1[22538] <= 16'b1111111111111001;
        weights1[22539] <= 16'b1111111111101101;
        weights1[22540] <= 16'b0000000000000010;
        weights1[22541] <= 16'b1111111111110100;
        weights1[22542] <= 16'b0000000000001000;
        weights1[22543] <= 16'b0000000000000010;
        weights1[22544] <= 16'b1111111111111001;
        weights1[22545] <= 16'b1111111111111001;
        weights1[22546] <= 16'b1111111111101000;
        weights1[22547] <= 16'b0000000000000111;
        weights1[22548] <= 16'b0000000000001010;
        weights1[22549] <= 16'b0000000000000100;
        weights1[22550] <= 16'b0000000000001100;
        weights1[22551] <= 16'b1111111111110100;
        weights1[22552] <= 16'b0000000000010010;
        weights1[22553] <= 16'b0000000000000111;
        weights1[22554] <= 16'b0000000000001010;
        weights1[22555] <= 16'b0000000000000101;
        weights1[22556] <= 16'b0000000000001001;
        weights1[22557] <= 16'b0000000000001100;
        weights1[22558] <= 16'b0000000000001110;
        weights1[22559] <= 16'b0000000000000110;
        weights1[22560] <= 16'b0000000000001110;
        weights1[22561] <= 16'b0000000000010011;
        weights1[22562] <= 16'b0000000000001110;
        weights1[22563] <= 16'b0000000000001110;
        weights1[22564] <= 16'b0000000000000001;
        weights1[22565] <= 16'b0000000000010000;
        weights1[22566] <= 16'b0000000000000111;
        weights1[22567] <= 16'b1111111111111001;
        weights1[22568] <= 16'b1111111111111100;
        weights1[22569] <= 16'b0000000000000110;
        weights1[22570] <= 16'b0000000000001101;
        weights1[22571] <= 16'b0000000000000101;
        weights1[22572] <= 16'b1111111111110110;
        weights1[22573] <= 16'b0000000000000001;
        weights1[22574] <= 16'b1111111111111010;
        weights1[22575] <= 16'b1111111111111001;
        weights1[22576] <= 16'b1111111111101010;
        weights1[22577] <= 16'b0000000000010001;
        weights1[22578] <= 16'b0000000000000001;
        weights1[22579] <= 16'b0000000000001100;
        weights1[22580] <= 16'b0000000000010001;
        weights1[22581] <= 16'b0000000000000101;
        weights1[22582] <= 16'b0000000000001000;
        weights1[22583] <= 16'b0000000000010010;
        weights1[22584] <= 16'b0000000000001011;
        weights1[22585] <= 16'b0000000000001010;
        weights1[22586] <= 16'b0000000000010010;
        weights1[22587] <= 16'b1111111111111010;
        weights1[22588] <= 16'b0000000000010100;
        weights1[22589] <= 16'b0000000000011001;
        weights1[22590] <= 16'b0000000000000110;
        weights1[22591] <= 16'b0000000000000100;
        weights1[22592] <= 16'b0000000000100100;
        weights1[22593] <= 16'b0000000000010100;
        weights1[22594] <= 16'b0000000000001100;
        weights1[22595] <= 16'b0000000000000010;
        weights1[22596] <= 16'b0000000000000000;
        weights1[22597] <= 16'b0000000000001100;
        weights1[22598] <= 16'b0000000000000101;
        weights1[22599] <= 16'b0000000000001101;
        weights1[22600] <= 16'b0000000000000011;
        weights1[22601] <= 16'b1111111111111111;
        weights1[22602] <= 16'b0000000000010001;
        weights1[22603] <= 16'b1111111111111100;
        weights1[22604] <= 16'b1111111111111001;
        weights1[22605] <= 16'b1111111111111001;
        weights1[22606] <= 16'b0000000000000110;
        weights1[22607] <= 16'b0000000000000110;
        weights1[22608] <= 16'b1111111111111111;
        weights1[22609] <= 16'b1111111111111111;
        weights1[22610] <= 16'b0000000000001000;
        weights1[22611] <= 16'b1111111111111101;
        weights1[22612] <= 16'b0000000000000001;
        weights1[22613] <= 16'b1111111111110111;
        weights1[22614] <= 16'b0000000000001001;
        weights1[22615] <= 16'b1111111111110010;
        weights1[22616] <= 16'b0000000000001101;
        weights1[22617] <= 16'b0000000000010001;
        weights1[22618] <= 16'b0000000000000111;
        weights1[22619] <= 16'b0000000000010110;
        weights1[22620] <= 16'b0000000000100100;
        weights1[22621] <= 16'b0000000000011101;
        weights1[22622] <= 16'b0000000000011011;
        weights1[22623] <= 16'b0000000000000001;
        weights1[22624] <= 16'b0000000000000000;
        weights1[22625] <= 16'b0000000000000010;
        weights1[22626] <= 16'b0000000000001110;
        weights1[22627] <= 16'b1111111111111101;
        weights1[22628] <= 16'b1111111111111000;
        weights1[22629] <= 16'b0000000000000010;
        weights1[22630] <= 16'b0000000000000011;
        weights1[22631] <= 16'b0000000000000100;
        weights1[22632] <= 16'b0000000000001000;
        weights1[22633] <= 16'b0000000000001000;
        weights1[22634] <= 16'b0000000000000100;
        weights1[22635] <= 16'b1111111111111101;
        weights1[22636] <= 16'b0000000000000011;
        weights1[22637] <= 16'b0000000000000100;
        weights1[22638] <= 16'b0000000000000000;
        weights1[22639] <= 16'b0000000000010001;
        weights1[22640] <= 16'b0000000000000101;
        weights1[22641] <= 16'b0000000000011010;
        weights1[22642] <= 16'b0000000000001101;
        weights1[22643] <= 16'b0000000000000001;
        weights1[22644] <= 16'b0000000000000101;
        weights1[22645] <= 16'b0000000000010011;
        weights1[22646] <= 16'b1111111111111110;
        weights1[22647] <= 16'b1111111111110100;
        weights1[22648] <= 16'b0000000000001011;
        weights1[22649] <= 16'b1111111111110111;
        weights1[22650] <= 16'b0000000000000011;
        weights1[22651] <= 16'b1111111111111111;
        weights1[22652] <= 16'b0000000000000000;
        weights1[22653] <= 16'b0000000000000110;
        weights1[22654] <= 16'b1111111111111100;
        weights1[22655] <= 16'b0000000000000011;
        weights1[22656] <= 16'b0000000000000100;
        weights1[22657] <= 16'b0000000000000000;
        weights1[22658] <= 16'b0000000000000010;
        weights1[22659] <= 16'b0000000000000110;
        weights1[22660] <= 16'b0000000000010101;
        weights1[22661] <= 16'b1111111111111011;
        weights1[22662] <= 16'b0000000000010001;
        weights1[22663] <= 16'b0000000000000001;
        weights1[22664] <= 16'b0000000000011001;
        weights1[22665] <= 16'b0000000000001000;
        weights1[22666] <= 16'b0000000000001001;
        weights1[22667] <= 16'b1111111111110111;
        weights1[22668] <= 16'b1111111111111001;
        weights1[22669] <= 16'b0000000000000000;
        weights1[22670] <= 16'b1111111111111101;
        weights1[22671] <= 16'b0000000000000001;
        weights1[22672] <= 16'b0000000000010000;
        weights1[22673] <= 16'b0000000000001100;
        weights1[22674] <= 16'b1111111111111111;
        weights1[22675] <= 16'b0000000000000010;
        weights1[22676] <= 16'b0000000000010011;
        weights1[22677] <= 16'b0000000000000011;
        weights1[22678] <= 16'b0000000000000010;
        weights1[22679] <= 16'b1111111111111100;
        weights1[22680] <= 16'b1111111111111111;
        weights1[22681] <= 16'b1111111111110110;
        weights1[22682] <= 16'b1111111111110110;
        weights1[22683] <= 16'b0000000000000011;
        weights1[22684] <= 16'b0000000000001001;
        weights1[22685] <= 16'b1111111111111111;
        weights1[22686] <= 16'b0000000000000001;
        weights1[22687] <= 16'b0000000000000001;
        weights1[22688] <= 16'b0000000000000001;
        weights1[22689] <= 16'b0000000000000000;
        weights1[22690] <= 16'b1111111111110011;
        weights1[22691] <= 16'b1111111111111111;
        weights1[22692] <= 16'b0000000000000001;
        weights1[22693] <= 16'b0000000000000100;
        weights1[22694] <= 16'b1111111111110101;
        weights1[22695] <= 16'b0000000000000110;
        weights1[22696] <= 16'b0000000000010011;
        weights1[22697] <= 16'b0000000000000100;
        weights1[22698] <= 16'b0000000000010011;
        weights1[22699] <= 16'b1111111111111010;
        weights1[22700] <= 16'b0000000000001010;
        weights1[22701] <= 16'b0000000000010111;
        weights1[22702] <= 16'b1111111111111000;
        weights1[22703] <= 16'b0000000000000100;
        weights1[22704] <= 16'b0000000000001110;
        weights1[22705] <= 16'b0000000000001001;
        weights1[22706] <= 16'b0000000000000010;
        weights1[22707] <= 16'b0000000000000000;
        weights1[22708] <= 16'b1111111111111110;
        weights1[22709] <= 16'b1111111111111100;
        weights1[22710] <= 16'b1111111111111101;
        weights1[22711] <= 16'b1111111111110111;
        weights1[22712] <= 16'b1111111111111000;
        weights1[22713] <= 16'b0000000000001100;
        weights1[22714] <= 16'b0000000000001001;
        weights1[22715] <= 16'b0000000000001100;
        weights1[22716] <= 16'b0000000000001000;
        weights1[22717] <= 16'b0000000000001110;
        weights1[22718] <= 16'b0000000000001010;
        weights1[22719] <= 16'b0000000000010111;
        weights1[22720] <= 16'b0000000000010001;
        weights1[22721] <= 16'b0000000000000000;
        weights1[22722] <= 16'b0000000000011000;
        weights1[22723] <= 16'b0000000000001010;
        weights1[22724] <= 16'b1111111111111000;
        weights1[22725] <= 16'b0000000000000000;
        weights1[22726] <= 16'b0000000000010010;
        weights1[22727] <= 16'b0000000000000111;
        weights1[22728] <= 16'b0000000000011010;
        weights1[22729] <= 16'b0000000000010000;
        weights1[22730] <= 16'b0000000000000110;
        weights1[22731] <= 16'b0000000000000100;
        weights1[22732] <= 16'b0000000000000101;
        weights1[22733] <= 16'b0000000000001001;
        weights1[22734] <= 16'b1111111111111111;
        weights1[22735] <= 16'b1111111111111111;
        weights1[22736] <= 16'b0000000000000000;
        weights1[22737] <= 16'b0000000000000000;
        weights1[22738] <= 16'b1111111111111110;
        weights1[22739] <= 16'b1111111111110011;
        weights1[22740] <= 16'b1111111111101011;
        weights1[22741] <= 16'b1111111111100011;
        weights1[22742] <= 16'b1111111111110000;
        weights1[22743] <= 16'b0000000000000001;
        weights1[22744] <= 16'b0000000000011001;
        weights1[22745] <= 16'b0000000000111011;
        weights1[22746] <= 16'b0000000001010000;
        weights1[22747] <= 16'b0000000001010111;
        weights1[22748] <= 16'b0000000001000101;
        weights1[22749] <= 16'b0000000000101000;
        weights1[22750] <= 16'b0000000000100010;
        weights1[22751] <= 16'b0000000000010001;
        weights1[22752] <= 16'b0000000000001100;
        weights1[22753] <= 16'b1111111111110011;
        weights1[22754] <= 16'b1111111111101010;
        weights1[22755] <= 16'b1111111111101110;
        weights1[22756] <= 16'b1111111111100101;
        weights1[22757] <= 16'b1111111111100111;
        weights1[22758] <= 16'b1111111111101100;
        weights1[22759] <= 16'b1111111111111110;
        weights1[22760] <= 16'b1111111111111011;
        weights1[22761] <= 16'b0000000000000001;
        weights1[22762] <= 16'b0000000000000010;
        weights1[22763] <= 16'b0000000000000001;
        weights1[22764] <= 16'b0000000000000000;
        weights1[22765] <= 16'b1111111111111110;
        weights1[22766] <= 16'b1111111111110111;
        weights1[22767] <= 16'b1111111111100111;
        weights1[22768] <= 16'b1111111111011110;
        weights1[22769] <= 16'b1111111111011101;
        weights1[22770] <= 16'b1111111111100011;
        weights1[22771] <= 16'b0000000000001110;
        weights1[22772] <= 16'b0000000000010110;
        weights1[22773] <= 16'b0000000000110010;
        weights1[22774] <= 16'b0000000001000101;
        weights1[22775] <= 16'b0000000000111110;
        weights1[22776] <= 16'b0000000000100111;
        weights1[22777] <= 16'b0000000000010010;
        weights1[22778] <= 16'b1111111111111010;
        weights1[22779] <= 16'b1111111111111110;
        weights1[22780] <= 16'b1111111111111111;
        weights1[22781] <= 16'b1111111111101001;
        weights1[22782] <= 16'b1111111111010010;
        weights1[22783] <= 16'b1111111111000100;
        weights1[22784] <= 16'b1111111110111111;
        weights1[22785] <= 16'b1111111111011001;
        weights1[22786] <= 16'b1111111111100011;
        weights1[22787] <= 16'b1111111111110010;
        weights1[22788] <= 16'b1111111111111001;
        weights1[22789] <= 16'b0000000000000100;
        weights1[22790] <= 16'b0000000000001010;
        weights1[22791] <= 16'b0000000000000000;
        weights1[22792] <= 16'b1111111111111100;
        weights1[22793] <= 16'b1111111111111000;
        weights1[22794] <= 16'b1111111111110000;
        weights1[22795] <= 16'b1111111111011101;
        weights1[22796] <= 16'b1111111111001011;
        weights1[22797] <= 16'b1111111111001111;
        weights1[22798] <= 16'b1111111111101110;
        weights1[22799] <= 16'b0000000000101111;
        weights1[22800] <= 16'b0000000000111010;
        weights1[22801] <= 16'b0000000001001010;
        weights1[22802] <= 16'b0000000000101110;
        weights1[22803] <= 16'b0000000000011111;
        weights1[22804] <= 16'b0000000000101110;
        weights1[22805] <= 16'b0000000000011101;
        weights1[22806] <= 16'b0000000000000111;
        weights1[22807] <= 16'b1111111111110011;
        weights1[22808] <= 16'b1111111111011100;
        weights1[22809] <= 16'b1111111110111001;
        weights1[22810] <= 16'b1111111110100011;
        weights1[22811] <= 16'b1111111110011110;
        weights1[22812] <= 16'b1111111110101100;
        weights1[22813] <= 16'b1111111111010101;
        weights1[22814] <= 16'b1111111111101100;
        weights1[22815] <= 16'b1111111111111010;
        weights1[22816] <= 16'b1111111111111010;
        weights1[22817] <= 16'b0000000000000001;
        weights1[22818] <= 16'b0000000000000110;
        weights1[22819] <= 16'b1111111111111101;
        weights1[22820] <= 16'b1111111111110110;
        weights1[22821] <= 16'b1111111111101111;
        weights1[22822] <= 16'b1111111111011110;
        weights1[22823] <= 16'b1111111111000111;
        weights1[22824] <= 16'b1111111111000001;
        weights1[22825] <= 16'b1111111111011110;
        weights1[22826] <= 16'b1111111111110101;
        weights1[22827] <= 16'b0000000000011111;
        weights1[22828] <= 16'b0000000000111110;
        weights1[22829] <= 16'b0000000001001001;
        weights1[22830] <= 16'b0000000000110011;
        weights1[22831] <= 16'b0000000000101101;
        weights1[22832] <= 16'b0000000000100110;
        weights1[22833] <= 16'b0000000000000111;
        weights1[22834] <= 16'b1111111111100101;
        weights1[22835] <= 16'b1111111111000001;
        weights1[22836] <= 16'b1111111110010111;
        weights1[22837] <= 16'b1111111101110110;
        weights1[22838] <= 16'b1111111110000100;
        weights1[22839] <= 16'b1111111110011001;
        weights1[22840] <= 16'b1111111111000010;
        weights1[22841] <= 16'b1111111111100101;
        weights1[22842] <= 16'b0000000000000010;
        weights1[22843] <= 16'b0000000000000010;
        weights1[22844] <= 16'b1111111111111101;
        weights1[22845] <= 16'b0000000000000100;
        weights1[22846] <= 16'b0000000000001110;
        weights1[22847] <= 16'b0000000000001000;
        weights1[22848] <= 16'b1111111111110101;
        weights1[22849] <= 16'b1111111111100111;
        weights1[22850] <= 16'b1111111111010100;
        weights1[22851] <= 16'b1111111110111010;
        weights1[22852] <= 16'b1111111111001100;
        weights1[22853] <= 16'b1111111111111100;
        weights1[22854] <= 16'b0000000000000011;
        weights1[22855] <= 16'b0000000000110100;
        weights1[22856] <= 16'b0000000001000111;
        weights1[22857] <= 16'b0000000000111001;
        weights1[22858] <= 16'b0000000000100101;
        weights1[22859] <= 16'b0000000000110101;
        weights1[22860] <= 16'b0000000000001001;
        weights1[22861] <= 16'b1111111111011110;
        weights1[22862] <= 16'b1111111110100100;
        weights1[22863] <= 16'b1111111101111110;
        weights1[22864] <= 16'b1111111101010111;
        weights1[22865] <= 16'b1111111101100010;
        weights1[22866] <= 16'b1111111110000111;
        weights1[22867] <= 16'b1111111111000111;
        weights1[22868] <= 16'b1111111111101000;
        weights1[22869] <= 16'b1111111111101010;
        weights1[22870] <= 16'b1111111111111111;
        weights1[22871] <= 16'b1111111111111111;
        weights1[22872] <= 16'b1111111111111011;
        weights1[22873] <= 16'b1111111111111010;
        weights1[22874] <= 16'b1111111111111110;
        weights1[22875] <= 16'b0000000000001001;
        weights1[22876] <= 16'b1111111111110100;
        weights1[22877] <= 16'b1111111111100110;
        weights1[22878] <= 16'b1111111111001100;
        weights1[22879] <= 16'b1111111110111110;
        weights1[22880] <= 16'b1111111111100000;
        weights1[22881] <= 16'b0000000000001100;
        weights1[22882] <= 16'b0000000000001010;
        weights1[22883] <= 16'b0000000000011001;
        weights1[22884] <= 16'b0000000000001000;
        weights1[22885] <= 16'b0000000000100000;
        weights1[22886] <= 16'b0000000000111110;
        weights1[22887] <= 16'b0000000000011100;
        weights1[22888] <= 16'b1111111111001100;
        weights1[22889] <= 16'b1111111110010011;
        weights1[22890] <= 16'b1111111110001010;
        weights1[22891] <= 16'b1111111101100010;
        weights1[22892] <= 16'b1111111110001000;
        weights1[22893] <= 16'b1111111111000111;
        weights1[22894] <= 16'b1111111111010100;
        weights1[22895] <= 16'b1111111111101111;
        weights1[22896] <= 16'b1111111111111111;
        weights1[22897] <= 16'b0000000000000101;
        weights1[22898] <= 16'b1111111111111100;
        weights1[22899] <= 16'b1111111111100111;
        weights1[22900] <= 16'b1111111111111000;
        weights1[22901] <= 16'b0000000000000001;
        weights1[22902] <= 16'b0000000000011100;
        weights1[22903] <= 16'b0000000000010001;
        weights1[22904] <= 16'b1111111111110110;
        weights1[22905] <= 16'b1111111111100000;
        weights1[22906] <= 16'b1111111111001010;
        weights1[22907] <= 16'b1111111111000011;
        weights1[22908] <= 16'b1111111111110010;
        weights1[22909] <= 16'b0000000000010010;
        weights1[22910] <= 16'b0000000000011000;
        weights1[22911] <= 16'b0000000000001100;
        weights1[22912] <= 16'b0000000000010100;
        weights1[22913] <= 16'b0000000000110111;
        weights1[22914] <= 16'b0000000000111011;
        weights1[22915] <= 16'b0000000000000111;
        weights1[22916] <= 16'b1111111110101000;
        weights1[22917] <= 16'b1111111110010000;
        weights1[22918] <= 16'b1111111101110001;
        weights1[22919] <= 16'b1111111101111011;
        weights1[22920] <= 16'b1111111110101011;
        weights1[22921] <= 16'b1111111111101111;
        weights1[22922] <= 16'b1111111111111000;
        weights1[22923] <= 16'b0000000000000111;
        weights1[22924] <= 16'b0000000000000111;
        weights1[22925] <= 16'b0000000000001101;
        weights1[22926] <= 16'b1111111111110111;
        weights1[22927] <= 16'b0000000000010101;
        weights1[22928] <= 16'b1111111111111011;
        weights1[22929] <= 16'b0000000000001101;
        weights1[22930] <= 16'b0000000000010101;
        weights1[22931] <= 16'b0000000000010000;
        weights1[22932] <= 16'b1111111111101110;
        weights1[22933] <= 16'b1111111111011100;
        weights1[22934] <= 16'b1111111111001001;
        weights1[22935] <= 16'b1111111111010110;
        weights1[22936] <= 16'b1111111111110111;
        weights1[22937] <= 16'b0000000000011100;
        weights1[22938] <= 16'b0000000000010110;
        weights1[22939] <= 16'b0000000000101100;
        weights1[22940] <= 16'b0000000000010011;
        weights1[22941] <= 16'b0000000000010110;
        weights1[22942] <= 16'b0000000000100111;
        weights1[22943] <= 16'b1111111111101011;
        weights1[22944] <= 16'b1111111101111011;
        weights1[22945] <= 16'b1111111110001001;
        weights1[22946] <= 16'b1111111110100111;
        weights1[22947] <= 16'b1111111110111000;
        weights1[22948] <= 16'b1111111111101110;
        weights1[22949] <= 16'b1111111111111010;
        weights1[22950] <= 16'b1111111111010011;
        weights1[22951] <= 16'b0000000000000010;
        weights1[22952] <= 16'b0000000000010000;
        weights1[22953] <= 16'b0000000000011110;
        weights1[22954] <= 16'b1111111111111101;
        weights1[22955] <= 16'b0000000000010111;
        weights1[22956] <= 16'b0000000000000110;
        weights1[22957] <= 16'b1111111111111101;
        weights1[22958] <= 16'b0000000000010000;
        weights1[22959] <= 16'b0000000000001110;
        weights1[22960] <= 16'b1111111111110100;
        weights1[22961] <= 16'b1111111111100010;
        weights1[22962] <= 16'b1111111111011001;
        weights1[22963] <= 16'b1111111111010100;
        weights1[22964] <= 16'b1111111111111100;
        weights1[22965] <= 16'b0000000000010001;
        weights1[22966] <= 16'b0000000000000000;
        weights1[22967] <= 16'b0000000000011110;
        weights1[22968] <= 16'b0000000000010111;
        weights1[22969] <= 16'b0000000000100001;
        weights1[22970] <= 16'b0000000000110001;
        weights1[22971] <= 16'b1111111111010000;
        weights1[22972] <= 16'b1111111110010000;
        weights1[22973] <= 16'b1111111111000010;
        weights1[22974] <= 16'b1111111111000100;
        weights1[22975] <= 16'b1111111111100100;
        weights1[22976] <= 16'b1111111111110111;
        weights1[22977] <= 16'b0000000000011011;
        weights1[22978] <= 16'b0000000000011011;
        weights1[22979] <= 16'b0000000000011101;
        weights1[22980] <= 16'b0000000000001010;
        weights1[22981] <= 16'b0000000000011001;
        weights1[22982] <= 16'b0000000000001110;
        weights1[22983] <= 16'b0000000000100100;
        weights1[22984] <= 16'b0000000000001110;
        weights1[22985] <= 16'b0000000000011010;
        weights1[22986] <= 16'b0000000000001001;
        weights1[22987] <= 16'b0000000000000101;
        weights1[22988] <= 16'b1111111111111000;
        weights1[22989] <= 16'b1111111111101110;
        weights1[22990] <= 16'b1111111111101010;
        weights1[22991] <= 16'b1111111111010111;
        weights1[22992] <= 16'b1111111111110011;
        weights1[22993] <= 16'b1111111111111100;
        weights1[22994] <= 16'b0000000000001000;
        weights1[22995] <= 16'b0000000000001011;
        weights1[22996] <= 16'b0000000000010000;
        weights1[22997] <= 16'b0000000000001100;
        weights1[22998] <= 16'b0000000000010100;
        weights1[22999] <= 16'b1111111111001111;
        weights1[23000] <= 16'b1111111110011100;
        weights1[23001] <= 16'b1111111111000001;
        weights1[23002] <= 16'b1111111111001101;
        weights1[23003] <= 16'b1111111111111010;
        weights1[23004] <= 16'b0000000000010101;
        weights1[23005] <= 16'b0000000000001011;
        weights1[23006] <= 16'b0000000000011011;
        weights1[23007] <= 16'b0000000000001100;
        weights1[23008] <= 16'b0000000000001000;
        weights1[23009] <= 16'b0000000000011110;
        weights1[23010] <= 16'b0000000000001011;
        weights1[23011] <= 16'b0000000000000111;
        weights1[23012] <= 16'b1111111111111110;
        weights1[23013] <= 16'b0000000000001101;
        weights1[23014] <= 16'b0000000000010011;
        weights1[23015] <= 16'b0000000000001011;
        weights1[23016] <= 16'b1111111111110111;
        weights1[23017] <= 16'b1111111111110101;
        weights1[23018] <= 16'b1111111111100001;
        weights1[23019] <= 16'b1111111111011110;
        weights1[23020] <= 16'b0000000000000000;
        weights1[23021] <= 16'b1111111111110011;
        weights1[23022] <= 16'b1111111111110010;
        weights1[23023] <= 16'b0000000000001010;
        weights1[23024] <= 16'b0000000000001111;
        weights1[23025] <= 16'b0000000000001101;
        weights1[23026] <= 16'b0000000000001001;
        weights1[23027] <= 16'b1111111110110011;
        weights1[23028] <= 16'b1111111110110010;
        weights1[23029] <= 16'b1111111111100100;
        weights1[23030] <= 16'b0000000000000110;
        weights1[23031] <= 16'b1111111111111110;
        weights1[23032] <= 16'b0000000000011110;
        weights1[23033] <= 16'b0000000000011111;
        weights1[23034] <= 16'b0000000000010001;
        weights1[23035] <= 16'b0000000000011011;
        weights1[23036] <= 16'b0000000000010011;
        weights1[23037] <= 16'b0000000000010001;
        weights1[23038] <= 16'b1111111111111011;
        weights1[23039] <= 16'b0000000000000010;
        weights1[23040] <= 16'b0000000000011010;
        weights1[23041] <= 16'b0000000000001010;
        weights1[23042] <= 16'b0000000000011101;
        weights1[23043] <= 16'b0000000000001100;
        weights1[23044] <= 16'b0000000000000001;
        weights1[23045] <= 16'b1111111111111001;
        weights1[23046] <= 16'b1111111111100000;
        weights1[23047] <= 16'b1111111111101101;
        weights1[23048] <= 16'b1111111111110000;
        weights1[23049] <= 16'b1111111111110010;
        weights1[23050] <= 16'b1111111111111101;
        weights1[23051] <= 16'b0000000000010000;
        weights1[23052] <= 16'b0000000000010000;
        weights1[23053] <= 16'b0000000000100000;
        weights1[23054] <= 16'b1111111111101000;
        weights1[23055] <= 16'b1111111111010000;
        weights1[23056] <= 16'b1111111111001010;
        weights1[23057] <= 16'b1111111111110001;
        weights1[23058] <= 16'b0000000000000000;
        weights1[23059] <= 16'b0000000000001000;
        weights1[23060] <= 16'b0000000000100000;
        weights1[23061] <= 16'b0000000000001111;
        weights1[23062] <= 16'b0000000000101001;
        weights1[23063] <= 16'b0000000000000100;
        weights1[23064] <= 16'b0000000000010010;
        weights1[23065] <= 16'b0000000000001100;
        weights1[23066] <= 16'b0000000000001000;
        weights1[23067] <= 16'b0000000000010011;
        weights1[23068] <= 16'b0000000000000011;
        weights1[23069] <= 16'b1111111111110100;
        weights1[23070] <= 16'b0000000000000011;
        weights1[23071] <= 16'b0000000000010101;
        weights1[23072] <= 16'b1111111111111111;
        weights1[23073] <= 16'b1111111111110111;
        weights1[23074] <= 16'b1111111111101111;
        weights1[23075] <= 16'b1111111111100100;
        weights1[23076] <= 16'b0000000000000011;
        weights1[23077] <= 16'b0000000000001001;
        weights1[23078] <= 16'b0000000000000011;
        weights1[23079] <= 16'b0000000000001110;
        weights1[23080] <= 16'b1111111111110100;
        weights1[23081] <= 16'b0000000000010000;
        weights1[23082] <= 16'b1111111111101001;
        weights1[23083] <= 16'b1111111111001000;
        weights1[23084] <= 16'b1111111111010001;
        weights1[23085] <= 16'b1111111111110000;
        weights1[23086] <= 16'b0000000000000110;
        weights1[23087] <= 16'b0000000000001101;
        weights1[23088] <= 16'b0000000000001110;
        weights1[23089] <= 16'b0000000000000101;
        weights1[23090] <= 16'b0000000000010000;
        weights1[23091] <= 16'b0000000000010011;
        weights1[23092] <= 16'b1111111111111000;
        weights1[23093] <= 16'b1111111111010101;
        weights1[23094] <= 16'b1111111111000110;
        weights1[23095] <= 16'b1111111111000001;
        weights1[23096] <= 16'b1111111111001111;
        weights1[23097] <= 16'b1111111111000010;
        weights1[23098] <= 16'b1111111111011100;
        weights1[23099] <= 16'b1111111111101000;
        weights1[23100] <= 16'b1111111111111010;
        weights1[23101] <= 16'b0000000000000000;
        weights1[23102] <= 16'b0000000000000010;
        weights1[23103] <= 16'b1111111111111111;
        weights1[23104] <= 16'b1111111111111100;
        weights1[23105] <= 16'b1111111111111000;
        weights1[23106] <= 16'b1111111111111100;
        weights1[23107] <= 16'b1111111111111000;
        weights1[23108] <= 16'b0000000000001110;
        weights1[23109] <= 16'b0000000000010001;
        weights1[23110] <= 16'b0000000000001000;
        weights1[23111] <= 16'b1111111111100101;
        weights1[23112] <= 16'b1111111111110001;
        weights1[23113] <= 16'b1111111111110101;
        weights1[23114] <= 16'b0000000000001010;
        weights1[23115] <= 16'b0000000000000010;
        weights1[23116] <= 16'b0000000000001111;
        weights1[23117] <= 16'b1111111111111110;
        weights1[23118] <= 16'b0000000000000011;
        weights1[23119] <= 16'b1111111111101001;
        weights1[23120] <= 16'b1111111111011011;
        weights1[23121] <= 16'b1111111111001110;
        weights1[23122] <= 16'b1111111111001110;
        weights1[23123] <= 16'b1111111111000000;
        weights1[23124] <= 16'b1111111111000111;
        weights1[23125] <= 16'b1111111111000000;
        weights1[23126] <= 16'b1111111111001001;
        weights1[23127] <= 16'b1111111111011100;
        weights1[23128] <= 16'b1111111111111000;
        weights1[23129] <= 16'b1111111111111111;
        weights1[23130] <= 16'b1111111111111110;
        weights1[23131] <= 16'b0000000000000111;
        weights1[23132] <= 16'b0000000000000011;
        weights1[23133] <= 16'b1111111111111100;
        weights1[23134] <= 16'b0000000000010011;
        weights1[23135] <= 16'b1111111111111100;
        weights1[23136] <= 16'b0000000000000100;
        weights1[23137] <= 16'b1111111111110111;
        weights1[23138] <= 16'b0000000000010101;
        weights1[23139] <= 16'b1111111111111110;
        weights1[23140] <= 16'b1111111111101001;
        weights1[23141] <= 16'b1111111111111110;
        weights1[23142] <= 16'b1111111111111110;
        weights1[23143] <= 16'b0000000000010011;
        weights1[23144] <= 16'b0000000000000011;
        weights1[23145] <= 16'b1111111111111110;
        weights1[23146] <= 16'b1111111111110000;
        weights1[23147] <= 16'b1111111111101100;
        weights1[23148] <= 16'b1111111111110110;
        weights1[23149] <= 16'b1111111111110010;
        weights1[23150] <= 16'b0000000000000100;
        weights1[23151] <= 16'b1111111111110100;
        weights1[23152] <= 16'b1111111111100100;
        weights1[23153] <= 16'b1111111111010110;
        weights1[23154] <= 16'b1111111111011001;
        weights1[23155] <= 16'b1111111111100100;
        weights1[23156] <= 16'b1111111111111011;
        weights1[23157] <= 16'b1111111111111000;
        weights1[23158] <= 16'b1111111111111100;
        weights1[23159] <= 16'b1111111111110111;
        weights1[23160] <= 16'b1111111111110100;
        weights1[23161] <= 16'b0000000000000010;
        weights1[23162] <= 16'b1111111111111110;
        weights1[23163] <= 16'b0000000000010000;
        weights1[23164] <= 16'b1111111111111001;
        weights1[23165] <= 16'b0000000000011101;
        weights1[23166] <= 16'b0000000000000101;
        weights1[23167] <= 16'b0000000000000010;
        weights1[23168] <= 16'b1111111111111001;
        weights1[23169] <= 16'b0000000000000000;
        weights1[23170] <= 16'b1111111111110100;
        weights1[23171] <= 16'b0000000000000101;
        weights1[23172] <= 16'b0000000000000101;
        weights1[23173] <= 16'b1111111111101000;
        weights1[23174] <= 16'b1111111111101100;
        weights1[23175] <= 16'b1111111111101100;
        weights1[23176] <= 16'b0000000000000000;
        weights1[23177] <= 16'b0000000000000100;
        weights1[23178] <= 16'b1111111111111110;
        weights1[23179] <= 16'b0000000000001000;
        weights1[23180] <= 16'b1111111111111101;
        weights1[23181] <= 16'b1111111111110111;
        weights1[23182] <= 16'b1111111111110000;
        weights1[23183] <= 16'b1111111111101001;
        weights1[23184] <= 16'b1111111111110011;
        weights1[23185] <= 16'b1111111111111101;
        weights1[23186] <= 16'b0000000000000001;
        weights1[23187] <= 16'b0000000000000111;
        weights1[23188] <= 16'b0000000000000001;
        weights1[23189] <= 16'b0000000000001100;
        weights1[23190] <= 16'b0000000000010111;
        weights1[23191] <= 16'b0000000000001001;
        weights1[23192] <= 16'b0000000000001111;
        weights1[23193] <= 16'b0000000000010010;
        weights1[23194] <= 16'b1111111111111110;
        weights1[23195] <= 16'b0000000000001100;
        weights1[23196] <= 16'b1111111111111000;
        weights1[23197] <= 16'b0000000000001100;
        weights1[23198] <= 16'b1111111111101101;
        weights1[23199] <= 16'b1111111111111100;
        weights1[23200] <= 16'b1111111111111100;
        weights1[23201] <= 16'b0000000000000000;
        weights1[23202] <= 16'b1111111111101010;
        weights1[23203] <= 16'b1111111111110111;
        weights1[23204] <= 16'b1111111111011101;
        weights1[23205] <= 16'b1111111111101111;
        weights1[23206] <= 16'b1111111111110011;
        weights1[23207] <= 16'b0000000000001100;
        weights1[23208] <= 16'b0000000000001010;
        weights1[23209] <= 16'b0000000000001111;
        weights1[23210] <= 16'b0000000000001001;
        weights1[23211] <= 16'b1111111111111001;
        weights1[23212] <= 16'b1111111111110100;
        weights1[23213] <= 16'b0000000000001010;
        weights1[23214] <= 16'b0000000000001100;
        weights1[23215] <= 16'b1111111111111011;
        weights1[23216] <= 16'b1111111111110110;
        weights1[23217] <= 16'b0000000000001110;
        weights1[23218] <= 16'b0000000000000101;
        weights1[23219] <= 16'b0000000000000010;
        weights1[23220] <= 16'b1111111111111100;
        weights1[23221] <= 16'b0000000000001101;
        weights1[23222] <= 16'b1111111111111100;
        weights1[23223] <= 16'b0000000000010000;
        weights1[23224] <= 16'b0000000000000000;
        weights1[23225] <= 16'b0000000000000101;
        weights1[23226] <= 16'b1111111111101100;
        weights1[23227] <= 16'b1111111111111011;
        weights1[23228] <= 16'b1111111111111001;
        weights1[23229] <= 16'b1111111111110111;
        weights1[23230] <= 16'b0000000000001000;
        weights1[23231] <= 16'b1111111111101101;
        weights1[23232] <= 16'b1111111111111110;
        weights1[23233] <= 16'b1111111111111110;
        weights1[23234] <= 16'b0000000000010001;
        weights1[23235] <= 16'b1111111111111101;
        weights1[23236] <= 16'b0000000000000010;
        weights1[23237] <= 16'b0000000000001101;
        weights1[23238] <= 16'b0000000000000100;
        weights1[23239] <= 16'b1111111111111010;
        weights1[23240] <= 16'b1111111111110111;
        weights1[23241] <= 16'b0000000000010001;
        weights1[23242] <= 16'b0000000000001010;
        weights1[23243] <= 16'b1111111111111010;
        weights1[23244] <= 16'b1111111111010111;
        weights1[23245] <= 16'b0000000000000011;
        weights1[23246] <= 16'b1111111111110100;
        weights1[23247] <= 16'b0000000000001001;
        weights1[23248] <= 16'b1111111111111000;
        weights1[23249] <= 16'b0000000000000001;
        weights1[23250] <= 16'b0000000000000011;
        weights1[23251] <= 16'b0000000000001010;
        weights1[23252] <= 16'b0000000000001001;
        weights1[23253] <= 16'b1111111111101110;
        weights1[23254] <= 16'b1111111111111101;
        weights1[23255] <= 16'b1111111111110001;
        weights1[23256] <= 16'b1111111111110101;
        weights1[23257] <= 16'b1111111111110101;
        weights1[23258] <= 16'b1111111111111101;
        weights1[23259] <= 16'b1111111111111011;
        weights1[23260] <= 16'b1111111111110011;
        weights1[23261] <= 16'b1111111111110111;
        weights1[23262] <= 16'b0000000000001010;
        weights1[23263] <= 16'b0000000000011010;
        weights1[23264] <= 16'b0000000000000000;
        weights1[23265] <= 16'b0000000000000001;
        weights1[23266] <= 16'b0000000000001001;
        weights1[23267] <= 16'b1111111111110011;
        weights1[23268] <= 16'b1111111111111000;
        weights1[23269] <= 16'b0000000000001011;
        weights1[23270] <= 16'b0000000000010011;
        weights1[23271] <= 16'b0000000000001100;
        weights1[23272] <= 16'b1111111111110000;
        weights1[23273] <= 16'b1111111111111110;
        weights1[23274] <= 16'b0000000000011000;
        weights1[23275] <= 16'b1111111111111111;
        weights1[23276] <= 16'b1111111111110011;
        weights1[23277] <= 16'b0000000000010101;
        weights1[23278] <= 16'b0000000000000001;
        weights1[23279] <= 16'b0000000000001011;
        weights1[23280] <= 16'b0000000000000000;
        weights1[23281] <= 16'b0000000000001101;
        weights1[23282] <= 16'b0000000000001001;
        weights1[23283] <= 16'b1111111111111110;
        weights1[23284] <= 16'b1111111111111010;
        weights1[23285] <= 16'b1111111111111001;
        weights1[23286] <= 16'b1111111111111011;
        weights1[23287] <= 16'b1111111111100011;
        weights1[23288] <= 16'b0000000000001101;
        weights1[23289] <= 16'b0000000000000011;
        weights1[23290] <= 16'b0000000000010011;
        weights1[23291] <= 16'b0000000000000000;
        weights1[23292] <= 16'b1111111111111100;
        weights1[23293] <= 16'b0000000000000000;
        weights1[23294] <= 16'b0000000000000001;
        weights1[23295] <= 16'b0000000000000100;
        weights1[23296] <= 16'b0000000000000001;
        weights1[23297] <= 16'b1111111111111001;
        weights1[23298] <= 16'b0000000000001001;
        weights1[23299] <= 16'b0000000000001000;
        weights1[23300] <= 16'b0000000000001101;
        weights1[23301] <= 16'b1111111111110110;
        weights1[23302] <= 16'b0000000000000101;
        weights1[23303] <= 16'b1111111111111100;
        weights1[23304] <= 16'b0000000000000000;
        weights1[23305] <= 16'b0000000000001110;
        weights1[23306] <= 16'b0000000000010010;
        weights1[23307] <= 16'b1111111111111011;
        weights1[23308] <= 16'b0000000000010110;
        weights1[23309] <= 16'b0000000000000000;
        weights1[23310] <= 16'b0000000000000011;
        weights1[23311] <= 16'b1111111111111001;
        weights1[23312] <= 16'b1111111111110011;
        weights1[23313] <= 16'b1111111111111101;
        weights1[23314] <= 16'b1111111111110101;
        weights1[23315] <= 16'b0000000000000001;
        weights1[23316] <= 16'b1111111111111000;
        weights1[23317] <= 16'b1111111111111101;
        weights1[23318] <= 16'b1111111111111000;
        weights1[23319] <= 16'b1111111111111001;
        weights1[23320] <= 16'b0000000000010010;
        weights1[23321] <= 16'b1111111111111110;
        weights1[23322] <= 16'b0000000000000110;
        weights1[23323] <= 16'b0000000000000101;
        weights1[23324] <= 16'b0000000000000010;
        weights1[23325] <= 16'b1111111111111011;
        weights1[23326] <= 16'b1111111111111111;
        weights1[23327] <= 16'b0000000000000001;
        weights1[23328] <= 16'b0000000000010110;
        weights1[23329] <= 16'b0000000000001101;
        weights1[23330] <= 16'b0000000000000111;
        weights1[23331] <= 16'b1111111111111100;
        weights1[23332] <= 16'b0000000000010101;
        weights1[23333] <= 16'b1111111111110000;
        weights1[23334] <= 16'b1111111111111110;
        weights1[23335] <= 16'b1111111111111001;
        weights1[23336] <= 16'b1111111111111101;
        weights1[23337] <= 16'b1111111111110011;
        weights1[23338] <= 16'b1111111111111101;
        weights1[23339] <= 16'b0000000000001100;
        weights1[23340] <= 16'b1111111111111110;
        weights1[23341] <= 16'b1111111111110001;
        weights1[23342] <= 16'b1111111111110111;
        weights1[23343] <= 16'b1111111111110001;
        weights1[23344] <= 16'b0000000000000101;
        weights1[23345] <= 16'b0000000000010000;
        weights1[23346] <= 16'b1111111111111001;
        weights1[23347] <= 16'b0000000000000110;
        weights1[23348] <= 16'b0000000000010110;
        weights1[23349] <= 16'b1111111111110010;
        weights1[23350] <= 16'b0000000000000000;
        weights1[23351] <= 16'b1111111111110101;
        weights1[23352] <= 16'b0000000000000001;
        weights1[23353] <= 16'b1111111111111101;
        weights1[23354] <= 16'b1111111111111111;
        weights1[23355] <= 16'b1111111111110100;
        weights1[23356] <= 16'b0000000000001010;
        weights1[23357] <= 16'b0000000000000100;
        weights1[23358] <= 16'b0000000000001101;
        weights1[23359] <= 16'b1111111111101111;
        weights1[23360] <= 16'b1111111111111001;
        weights1[23361] <= 16'b0000000000000110;
        weights1[23362] <= 16'b0000000000010100;
        weights1[23363] <= 16'b0000000000000011;
        weights1[23364] <= 16'b0000000000001000;
        weights1[23365] <= 16'b0000000000000011;
        weights1[23366] <= 16'b1111111111111001;
        weights1[23367] <= 16'b1111111111111010;
        weights1[23368] <= 16'b1111111111111000;
        weights1[23369] <= 16'b1111111111110110;
        weights1[23370] <= 16'b0000000000001001;
        weights1[23371] <= 16'b1111111111111100;
        weights1[23372] <= 16'b1111111111111101;
        weights1[23373] <= 16'b1111111111101111;
        weights1[23374] <= 16'b0000000000000010;
        weights1[23375] <= 16'b0000000000001010;
        weights1[23376] <= 16'b0000000000010100;
        weights1[23377] <= 16'b1111111111111101;
        weights1[23378] <= 16'b1111111111111111;
        weights1[23379] <= 16'b1111111111111101;
        weights1[23380] <= 16'b1111111111111001;
        weights1[23381] <= 16'b1111111111111101;
        weights1[23382] <= 16'b1111111111111011;
        weights1[23383] <= 16'b0000000000000000;
        weights1[23384] <= 16'b1111111111111000;
        weights1[23385] <= 16'b0000000000000100;
        weights1[23386] <= 16'b0000000000000111;
        weights1[23387] <= 16'b1111111111111101;
        weights1[23388] <= 16'b0000000000000001;
        weights1[23389] <= 16'b0000000000000000;
        weights1[23390] <= 16'b0000000000001110;
        weights1[23391] <= 16'b0000000000000101;
        weights1[23392] <= 16'b0000000000001111;
        weights1[23393] <= 16'b0000000000000011;
        weights1[23394] <= 16'b0000000000001010;
        weights1[23395] <= 16'b0000000000010010;
        weights1[23396] <= 16'b0000000000000011;
        weights1[23397] <= 16'b0000000000000010;
        weights1[23398] <= 16'b0000000000000001;
        weights1[23399] <= 16'b1111111111110001;
        weights1[23400] <= 16'b0000000000000001;
        weights1[23401] <= 16'b0000000000001100;
        weights1[23402] <= 16'b0000000000010110;
        weights1[23403] <= 16'b1111111111111100;
        weights1[23404] <= 16'b1111111111110111;
        weights1[23405] <= 16'b0000000000000000;
        weights1[23406] <= 16'b0000000000000000;
        weights1[23407] <= 16'b1111111111110011;
        weights1[23408] <= 16'b1111111111111000;
        weights1[23409] <= 16'b1111111111111101;
        weights1[23410] <= 16'b0000000000000000;
        weights1[23411] <= 16'b1111111111101010;
        weights1[23412] <= 16'b1111111111111101;
        weights1[23413] <= 16'b0000000000000010;
        weights1[23414] <= 16'b1111111111110010;
        weights1[23415] <= 16'b1111111111110100;
        weights1[23416] <= 16'b1111111111110001;
        weights1[23417] <= 16'b1111111111111011;
        weights1[23418] <= 16'b1111111111110000;
        weights1[23419] <= 16'b0000000000000001;
        weights1[23420] <= 16'b0000000000000010;
        weights1[23421] <= 16'b1111111111111110;
        weights1[23422] <= 16'b0000000000000100;
        weights1[23423] <= 16'b1111111111111011;
        weights1[23424] <= 16'b1111111111111111;
        weights1[23425] <= 16'b0000000000001110;
        weights1[23426] <= 16'b0000000000000100;
        weights1[23427] <= 16'b0000000000001010;
        weights1[23428] <= 16'b0000000000001101;
        weights1[23429] <= 16'b0000000000001100;
        weights1[23430] <= 16'b0000000000000111;
        weights1[23431] <= 16'b0000000000000010;
        weights1[23432] <= 16'b1111111111111010;
        weights1[23433] <= 16'b1111111111111001;
        weights1[23434] <= 16'b1111111111111000;
        weights1[23435] <= 16'b1111111111110100;
        weights1[23436] <= 16'b1111111111111111;
        weights1[23437] <= 16'b1111111111110110;
        weights1[23438] <= 16'b1111111111110100;
        weights1[23439] <= 16'b1111111111111010;
        weights1[23440] <= 16'b1111111111111010;
        weights1[23441] <= 16'b0000000000001010;
        weights1[23442] <= 16'b1111111111110111;
        weights1[23443] <= 16'b1111111111111001;
        weights1[23444] <= 16'b0000000000001010;
        weights1[23445] <= 16'b1111111111111101;
        weights1[23446] <= 16'b1111111111111100;
        weights1[23447] <= 16'b0000000000001010;
        weights1[23448] <= 16'b1111111111101111;
        weights1[23449] <= 16'b1111111111111110;
        weights1[23450] <= 16'b1111111111111101;
        weights1[23451] <= 16'b0000000000000011;
        weights1[23452] <= 16'b0000000000010010;
        weights1[23453] <= 16'b1111111111111101;
        weights1[23454] <= 16'b0000000000010000;
        weights1[23455] <= 16'b1111111111110010;
        weights1[23456] <= 16'b1111111111110001;
        weights1[23457] <= 16'b0000000000001001;
        weights1[23458] <= 16'b0000000000001101;
        weights1[23459] <= 16'b0000000000000011;
        weights1[23460] <= 16'b1111111111100100;
        weights1[23461] <= 16'b1111111111111010;
        weights1[23462] <= 16'b0000000000000100;
        weights1[23463] <= 16'b1111111111111001;
        weights1[23464] <= 16'b1111111111111111;
        weights1[23465] <= 16'b1111111111111111;
        weights1[23466] <= 16'b1111111111110111;
        weights1[23467] <= 16'b1111111111111100;
        weights1[23468] <= 16'b0000000000000111;
        weights1[23469] <= 16'b1111111111110000;
        weights1[23470] <= 16'b1111111111110011;
        weights1[23471] <= 16'b1111111111110100;
        weights1[23472] <= 16'b1111111111110001;
        weights1[23473] <= 16'b1111111111111100;
        weights1[23474] <= 16'b0000000000001011;
        weights1[23475] <= 16'b1111111111110100;
        weights1[23476] <= 16'b1111111111111010;
        weights1[23477] <= 16'b1111111111110110;
        weights1[23478] <= 16'b1111111111111100;
        weights1[23479] <= 16'b1111111111101010;
        weights1[23480] <= 16'b1111111111110001;
        weights1[23481] <= 16'b1111111111110100;
        weights1[23482] <= 16'b1111111111111001;
        weights1[23483] <= 16'b1111111111101100;
        weights1[23484] <= 16'b0000000000001001;
        weights1[23485] <= 16'b1111111111011100;
        weights1[23486] <= 16'b1111111111111011;
        weights1[23487] <= 16'b1111111111111000;
        weights1[23488] <= 16'b1111111111101111;
        weights1[23489] <= 16'b1111111111111001;
        weights1[23490] <= 16'b1111111111110110;
        weights1[23491] <= 16'b1111111111111010;
        weights1[23492] <= 16'b0000000000000000;
        weights1[23493] <= 16'b0000000000000111;
        weights1[23494] <= 16'b0000000000000001;
        weights1[23495] <= 16'b1111111111111111;
        weights1[23496] <= 16'b0000000000000010;
        weights1[23497] <= 16'b1111111111110110;
        weights1[23498] <= 16'b1111111111101001;
        weights1[23499] <= 16'b1111111111111011;
        weights1[23500] <= 16'b0000000000000010;
        weights1[23501] <= 16'b1111111111111000;
        weights1[23502] <= 16'b1111111111110000;
        weights1[23503] <= 16'b1111111111110010;
        weights1[23504] <= 16'b1111111111111010;
        weights1[23505] <= 16'b1111111111110111;
        weights1[23506] <= 16'b1111111111110111;
        weights1[23507] <= 16'b1111111111110010;
        weights1[23508] <= 16'b1111111111111110;
        weights1[23509] <= 16'b1111111111111011;
        weights1[23510] <= 16'b0000000000000000;
        weights1[23511] <= 16'b1111111111111011;
        weights1[23512] <= 16'b1111111111111010;
        weights1[23513] <= 16'b1111111111100110;
        weights1[23514] <= 16'b1111111111111000;
        weights1[23515] <= 16'b1111111111101010;
        weights1[23516] <= 16'b1111111111101101;
        weights1[23517] <= 16'b1111111111111000;
        weights1[23518] <= 16'b1111111111111010;
        weights1[23519] <= 16'b1111111111111110;
        weights1[23520] <= 16'b0000000000000000;
        weights1[23521] <= 16'b0000000000000000;
        weights1[23522] <= 16'b0000000000000001;
        weights1[23523] <= 16'b0000000000000010;
        weights1[23524] <= 16'b0000000000000001;
        weights1[23525] <= 16'b0000000000000010;
        weights1[23526] <= 16'b1111111111111100;
        weights1[23527] <= 16'b0000000000000011;
        weights1[23528] <= 16'b1111111111111000;
        weights1[23529] <= 16'b1111111111111111;
        weights1[23530] <= 16'b1111111111111100;
        weights1[23531] <= 16'b0000000000000100;
        weights1[23532] <= 16'b0000000000010001;
        weights1[23533] <= 16'b0000000000010000;
        weights1[23534] <= 16'b0000000000011100;
        weights1[23535] <= 16'b0000000000001110;
        weights1[23536] <= 16'b0000000000000001;
        weights1[23537] <= 16'b1111111111110110;
        weights1[23538] <= 16'b1111111111110100;
        weights1[23539] <= 16'b1111111111111001;
        weights1[23540] <= 16'b1111111111110110;
        weights1[23541] <= 16'b1111111111110100;
        weights1[23542] <= 16'b1111111111111010;
        weights1[23543] <= 16'b1111111111111001;
        weights1[23544] <= 16'b1111111111111100;
        weights1[23545] <= 16'b1111111111111111;
        weights1[23546] <= 16'b0000000000000000;
        weights1[23547] <= 16'b0000000000000000;
        weights1[23548] <= 16'b0000000000000000;
        weights1[23549] <= 16'b0000000000000000;
        weights1[23550] <= 16'b0000000000000001;
        weights1[23551] <= 16'b0000000000000001;
        weights1[23552] <= 16'b0000000000000000;
        weights1[23553] <= 16'b1111111111111111;
        weights1[23554] <= 16'b1111111111111000;
        weights1[23555] <= 16'b1111111111101111;
        weights1[23556] <= 16'b1111111111101101;
        weights1[23557] <= 16'b1111111111110111;
        weights1[23558] <= 16'b0000000000000010;
        weights1[23559] <= 16'b0000000000000011;
        weights1[23560] <= 16'b1111111111111111;
        weights1[23561] <= 16'b1111111111111110;
        weights1[23562] <= 16'b0000000000010010;
        weights1[23563] <= 16'b0000000000010111;
        weights1[23564] <= 16'b1111111111111101;
        weights1[23565] <= 16'b0000000000000110;
        weights1[23566] <= 16'b0000000000001001;
        weights1[23567] <= 16'b1111111111111111;
        weights1[23568] <= 16'b1111111111101100;
        weights1[23569] <= 16'b1111111111110011;
        weights1[23570] <= 16'b1111111111110101;
        weights1[23571] <= 16'b1111111111101100;
        weights1[23572] <= 16'b1111111111111100;
        weights1[23573] <= 16'b0000000000000000;
        weights1[23574] <= 16'b0000000000000001;
        weights1[23575] <= 16'b0000000000000000;
        weights1[23576] <= 16'b0000000000000000;
        weights1[23577] <= 16'b0000000000000000;
        weights1[23578] <= 16'b0000000000000000;
        weights1[23579] <= 16'b0000000000000001;
        weights1[23580] <= 16'b1111111111110111;
        weights1[23581] <= 16'b1111111111110101;
        weights1[23582] <= 16'b1111111111110010;
        weights1[23583] <= 16'b1111111111100101;
        weights1[23584] <= 16'b1111111111011011;
        weights1[23585] <= 16'b1111111111100011;
        weights1[23586] <= 16'b1111111111011101;
        weights1[23587] <= 16'b1111111111100011;
        weights1[23588] <= 16'b1111111111100001;
        weights1[23589] <= 16'b1111111111111011;
        weights1[23590] <= 16'b0000000000000001;
        weights1[23591] <= 16'b1111111111111111;
        weights1[23592] <= 16'b1111111111110110;
        weights1[23593] <= 16'b1111111111110110;
        weights1[23594] <= 16'b1111111111111111;
        weights1[23595] <= 16'b0000000000000110;
        weights1[23596] <= 16'b1111111111101111;
        weights1[23597] <= 16'b1111111111110100;
        weights1[23598] <= 16'b1111111111101010;
        weights1[23599] <= 16'b1111111111101110;
        weights1[23600] <= 16'b1111111111110111;
        weights1[23601] <= 16'b1111111111111111;
        weights1[23602] <= 16'b0000000000000000;
        weights1[23603] <= 16'b0000000000000000;
        weights1[23604] <= 16'b0000000000000001;
        weights1[23605] <= 16'b0000000000000001;
        weights1[23606] <= 16'b0000000000000001;
        weights1[23607] <= 16'b1111111111111111;
        weights1[23608] <= 16'b1111111111110110;
        weights1[23609] <= 16'b1111111111110000;
        weights1[23610] <= 16'b1111111111101100;
        weights1[23611] <= 16'b1111111111011011;
        weights1[23612] <= 16'b1111111111000101;
        weights1[23613] <= 16'b1111111111000111;
        weights1[23614] <= 16'b1111111111001101;
        weights1[23615] <= 16'b1111111111100111;
        weights1[23616] <= 16'b1111111111101111;
        weights1[23617] <= 16'b1111111111111000;
        weights1[23618] <= 16'b1111111111111000;
        weights1[23619] <= 16'b1111111111110011;
        weights1[23620] <= 16'b1111111111110001;
        weights1[23621] <= 16'b1111111111110000;
        weights1[23622] <= 16'b1111111111110111;
        weights1[23623] <= 16'b1111111111110000;
        weights1[23624] <= 16'b1111111111100100;
        weights1[23625] <= 16'b1111111111100111;
        weights1[23626] <= 16'b1111111111111000;
        weights1[23627] <= 16'b1111111111110101;
        weights1[23628] <= 16'b1111111111110100;
        weights1[23629] <= 16'b1111111111111000;
        weights1[23630] <= 16'b1111111111111111;
        weights1[23631] <= 16'b0000000000000000;
        weights1[23632] <= 16'b1111111111111111;
        weights1[23633] <= 16'b0000000000000000;
        weights1[23634] <= 16'b0000000000000000;
        weights1[23635] <= 16'b1111111111110101;
        weights1[23636] <= 16'b1111111111111011;
        weights1[23637] <= 16'b1111111111110111;
        weights1[23638] <= 16'b1111111111101110;
        weights1[23639] <= 16'b1111111111010110;
        weights1[23640] <= 16'b1111111111101010;
        weights1[23641] <= 16'b1111111111101101;
        weights1[23642] <= 16'b1111111111111011;
        weights1[23643] <= 16'b0000000000000000;
        weights1[23644] <= 16'b1111111111101111;
        weights1[23645] <= 16'b0000000000010110;
        weights1[23646] <= 16'b1111111111111010;
        weights1[23647] <= 16'b0000000000001111;
        weights1[23648] <= 16'b0000000000001000;
        weights1[23649] <= 16'b0000000000001100;
        weights1[23650] <= 16'b0000000000010011;
        weights1[23651] <= 16'b1111111111111000;
        weights1[23652] <= 16'b1111111111111010;
        weights1[23653] <= 16'b1111111111110100;
        weights1[23654] <= 16'b1111111111010010;
        weights1[23655] <= 16'b1111111111100010;
        weights1[23656] <= 16'b1111111111110001;
        weights1[23657] <= 16'b1111111111110110;
        weights1[23658] <= 16'b1111111111111110;
        weights1[23659] <= 16'b1111111111111111;
        weights1[23660] <= 16'b1111111111111101;
        weights1[23661] <= 16'b0000000000000011;
        weights1[23662] <= 16'b1111111111111110;
        weights1[23663] <= 16'b1111111111111111;
        weights1[23664] <= 16'b0000000000000000;
        weights1[23665] <= 16'b1111111111111111;
        weights1[23666] <= 16'b0000000000000100;
        weights1[23667] <= 16'b0000000000000101;
        weights1[23668] <= 16'b1111111111110111;
        weights1[23669] <= 16'b0000000000010001;
        weights1[23670] <= 16'b1111111111111000;
        weights1[23671] <= 16'b1111111111111011;
        weights1[23672] <= 16'b0000000000000000;
        weights1[23673] <= 16'b0000000000100011;
        weights1[23674] <= 16'b0000000000000011;
        weights1[23675] <= 16'b0000000000001001;
        weights1[23676] <= 16'b0000000000010101;
        weights1[23677] <= 16'b1111111111111011;
        weights1[23678] <= 16'b0000000000000001;
        weights1[23679] <= 16'b0000000000001010;
        weights1[23680] <= 16'b1111111111111010;
        weights1[23681] <= 16'b1111111111010011;
        weights1[23682] <= 16'b1111111111000111;
        weights1[23683] <= 16'b1111111111000000;
        weights1[23684] <= 16'b1111111111101011;
        weights1[23685] <= 16'b1111111111110010;
        weights1[23686] <= 16'b1111111111111100;
        weights1[23687] <= 16'b0000000000000010;
        weights1[23688] <= 16'b1111111111111111;
        weights1[23689] <= 16'b0000000000000001;
        weights1[23690] <= 16'b1111111111111100;
        weights1[23691] <= 16'b0000000000000110;
        weights1[23692] <= 16'b0000000000001001;
        weights1[23693] <= 16'b0000000000010101;
        weights1[23694] <= 16'b0000000000010001;
        weights1[23695] <= 16'b0000000000011110;
        weights1[23696] <= 16'b0000000000011001;
        weights1[23697] <= 16'b0000000000011110;
        weights1[23698] <= 16'b0000000000011000;
        weights1[23699] <= 16'b0000000000000001;
        weights1[23700] <= 16'b1111111111111111;
        weights1[23701] <= 16'b0000000000011111;
        weights1[23702] <= 16'b0000000000010001;
        weights1[23703] <= 16'b0000000000001001;
        weights1[23704] <= 16'b0000000000000101;
        weights1[23705] <= 16'b0000000000000100;
        weights1[23706] <= 16'b0000000000000100;
        weights1[23707] <= 16'b1111111111111011;
        weights1[23708] <= 16'b0000000000010110;
        weights1[23709] <= 16'b1111111111001011;
        weights1[23710] <= 16'b1111111111010111;
        weights1[23711] <= 16'b1111111111001010;
        weights1[23712] <= 16'b1111111111101110;
        weights1[23713] <= 16'b1111111111110101;
        weights1[23714] <= 16'b1111111111111010;
        weights1[23715] <= 16'b1111111111111101;
        weights1[23716] <= 16'b0000000000000000;
        weights1[23717] <= 16'b0000000000000011;
        weights1[23718] <= 16'b0000000000001000;
        weights1[23719] <= 16'b0000000000001011;
        weights1[23720] <= 16'b0000000000010011;
        weights1[23721] <= 16'b0000000000001011;
        weights1[23722] <= 16'b0000000000100101;
        weights1[23723] <= 16'b0000000000111000;
        weights1[23724] <= 16'b0000000000100001;
        weights1[23725] <= 16'b0000000000100011;
        weights1[23726] <= 16'b0000000000101101;
        weights1[23727] <= 16'b0000000000010001;
        weights1[23728] <= 16'b0000000000110100;
        weights1[23729] <= 16'b0000000000011100;
        weights1[23730] <= 16'b0000000000101011;
        weights1[23731] <= 16'b0000000000001100;
        weights1[23732] <= 16'b0000000000000101;
        weights1[23733] <= 16'b0000000000101011;
        weights1[23734] <= 16'b0000000000000010;
        weights1[23735] <= 16'b1111111111110110;
        weights1[23736] <= 16'b0000000000001000;
        weights1[23737] <= 16'b1111111111110010;
        weights1[23738] <= 16'b1111111111101001;
        weights1[23739] <= 16'b1111111111010011;
        weights1[23740] <= 16'b1111111111100101;
        weights1[23741] <= 16'b1111111111110011;
        weights1[23742] <= 16'b1111111111111010;
        weights1[23743] <= 16'b1111111111111101;
        weights1[23744] <= 16'b0000000000000010;
        weights1[23745] <= 16'b0000000000001001;
        weights1[23746] <= 16'b0000000000001001;
        weights1[23747] <= 16'b0000000000001100;
        weights1[23748] <= 16'b0000000000011000;
        weights1[23749] <= 16'b0000000000011001;
        weights1[23750] <= 16'b0000000000010110;
        weights1[23751] <= 16'b0000000000100101;
        weights1[23752] <= 16'b0000000000011111;
        weights1[23753] <= 16'b0000000000111010;
        weights1[23754] <= 16'b0000000000111101;
        weights1[23755] <= 16'b0000000000011100;
        weights1[23756] <= 16'b1111111111111000;
        weights1[23757] <= 16'b0000000000010010;
        weights1[23758] <= 16'b0000000000001101;
        weights1[23759] <= 16'b0000000000100000;
        weights1[23760] <= 16'b0000000000010100;
        weights1[23761] <= 16'b0000000000010100;
        weights1[23762] <= 16'b0000000000001010;
        weights1[23763] <= 16'b0000000000000111;
        weights1[23764] <= 16'b1111111111100100;
        weights1[23765] <= 16'b1111111111110011;
        weights1[23766] <= 16'b1111111111011100;
        weights1[23767] <= 16'b1111111111000101;
        weights1[23768] <= 16'b1111111111001000;
        weights1[23769] <= 16'b1111111111101011;
        weights1[23770] <= 16'b1111111111110110;
        weights1[23771] <= 16'b1111111111111011;
        weights1[23772] <= 16'b0000000000000011;
        weights1[23773] <= 16'b0000000000001101;
        weights1[23774] <= 16'b1111111111111100;
        weights1[23775] <= 16'b0000000000000110;
        weights1[23776] <= 16'b0000000000101001;
        weights1[23777] <= 16'b0000000000001000;
        weights1[23778] <= 16'b0000000000101001;
        weights1[23779] <= 16'b0000000001000111;
        weights1[23780] <= 16'b0000000000111111;
        weights1[23781] <= 16'b0000000000111010;
        weights1[23782] <= 16'b1111111111111011;
        weights1[23783] <= 16'b1111111111011000;
        weights1[23784] <= 16'b1111111110000110;
        weights1[23785] <= 16'b1111111110111010;
        weights1[23786] <= 16'b1111111111110111;
        weights1[23787] <= 16'b0000000000000110;
        weights1[23788] <= 16'b0000000000001110;
        weights1[23789] <= 16'b0000000000001111;
        weights1[23790] <= 16'b1111111111111110;
        weights1[23791] <= 16'b0000000000001000;
        weights1[23792] <= 16'b1111111111101000;
        weights1[23793] <= 16'b1111111111111111;
        weights1[23794] <= 16'b1111111111011100;
        weights1[23795] <= 16'b1111111111011001;
        weights1[23796] <= 16'b1111111111100111;
        weights1[23797] <= 16'b1111111111110010;
        weights1[23798] <= 16'b1111111111110011;
        weights1[23799] <= 16'b1111111111111010;
        weights1[23800] <= 16'b0000000000000110;
        weights1[23801] <= 16'b0000000000000100;
        weights1[23802] <= 16'b1111111111110101;
        weights1[23803] <= 16'b1111111111111110;
        weights1[23804] <= 16'b0000000000010111;
        weights1[23805] <= 16'b0000000000011101;
        weights1[23806] <= 16'b0000000000001100;
        weights1[23807] <= 16'b1111111111110000;
        weights1[23808] <= 16'b1111111111000100;
        weights1[23809] <= 16'b1111111101110010;
        weights1[23810] <= 16'b1111111100011001;
        weights1[23811] <= 16'b1111111011111010;
        weights1[23812] <= 16'b1111111110100000;
        weights1[23813] <= 16'b1111111111011001;
        weights1[23814] <= 16'b1111111111111100;
        weights1[23815] <= 16'b0000000000001111;
        weights1[23816] <= 16'b0000000000010100;
        weights1[23817] <= 16'b0000000000011101;
        weights1[23818] <= 16'b0000000000000001;
        weights1[23819] <= 16'b1111111111101111;
        weights1[23820] <= 16'b1111111111100111;
        weights1[23821] <= 16'b1111111111011110;
        weights1[23822] <= 16'b1111111111011001;
        weights1[23823] <= 16'b1111111111100010;
        weights1[23824] <= 16'b1111111111110001;
        weights1[23825] <= 16'b1111111111110000;
        weights1[23826] <= 16'b1111111111111010;
        weights1[23827] <= 16'b1111111111110110;
        weights1[23828] <= 16'b1111111111111110;
        weights1[23829] <= 16'b1111111111110011;
        weights1[23830] <= 16'b1111111111101100;
        weights1[23831] <= 16'b1111111111100111;
        weights1[23832] <= 16'b1111111111111100;
        weights1[23833] <= 16'b1111111111100011;
        weights1[23834] <= 16'b1111111110111001;
        weights1[23835] <= 16'b1111111101100111;
        weights1[23836] <= 16'b1111111100011001;
        weights1[23837] <= 16'b1111111011011001;
        weights1[23838] <= 16'b1111111101011100;
        weights1[23839] <= 16'b1111111111100101;
        weights1[23840] <= 16'b1111111111101100;
        weights1[23841] <= 16'b0000000000000111;
        weights1[23842] <= 16'b0000000000011010;
        weights1[23843] <= 16'b0000000000010110;
        weights1[23844] <= 16'b0000000000011000;
        weights1[23845] <= 16'b1111111111111111;
        weights1[23846] <= 16'b0000000000001110;
        weights1[23847] <= 16'b1111111111110010;
        weights1[23848] <= 16'b1111111111111010;
        weights1[23849] <= 16'b1111111111011010;
        weights1[23850] <= 16'b1111111111011011;
        weights1[23851] <= 16'b1111111111110011;
        weights1[23852] <= 16'b1111111111110101;
        weights1[23853] <= 16'b1111111111111011;
        weights1[23854] <= 16'b1111111111111011;
        weights1[23855] <= 16'b1111111111111000;
        weights1[23856] <= 16'b1111111111110011;
        weights1[23857] <= 16'b1111111111100011;
        weights1[23858] <= 16'b1111111111010100;
        weights1[23859] <= 16'b1111111111000000;
        weights1[23860] <= 16'b1111111110101101;
        weights1[23861] <= 16'b1111111110011000;
        weights1[23862] <= 16'b1111111101101101;
        weights1[23863] <= 16'b1111111100110110;
        weights1[23864] <= 16'b1111111100110010;
        weights1[23865] <= 16'b1111111110111010;
        weights1[23866] <= 16'b0000000000001000;
        weights1[23867] <= 16'b0000000000100001;
        weights1[23868] <= 16'b0000000000010011;
        weights1[23869] <= 16'b0000000000001001;
        weights1[23870] <= 16'b0000000000010010;
        weights1[23871] <= 16'b0000000000001010;
        weights1[23872] <= 16'b0000000000011010;
        weights1[23873] <= 16'b0000000000010100;
        weights1[23874] <= 16'b0000000000001011;
        weights1[23875] <= 16'b1111111111101111;
        weights1[23876] <= 16'b1111111111011011;
        weights1[23877] <= 16'b1111111111101010;
        weights1[23878] <= 16'b1111111111101100;
        weights1[23879] <= 16'b1111111111111110;
        weights1[23880] <= 16'b1111111111111010;
        weights1[23881] <= 16'b1111111111111010;
        weights1[23882] <= 16'b1111111111111001;
        weights1[23883] <= 16'b0000000000000011;
        weights1[23884] <= 16'b1111111111100010;
        weights1[23885] <= 16'b1111111111010111;
        weights1[23886] <= 16'b1111111111000011;
        weights1[23887] <= 16'b1111111110101001;
        weights1[23888] <= 16'b1111111110100101;
        weights1[23889] <= 16'b1111111110000110;
        weights1[23890] <= 16'b1111111101101101;
        weights1[23891] <= 16'b1111111110001110;
        weights1[23892] <= 16'b1111111111000101;
        weights1[23893] <= 16'b0000000000000110;
        weights1[23894] <= 16'b0000000000101010;
        weights1[23895] <= 16'b0000000000011011;
        weights1[23896] <= 16'b0000000000010100;
        weights1[23897] <= 16'b0000000000001000;
        weights1[23898] <= 16'b0000000000100101;
        weights1[23899] <= 16'b0000000000001011;
        weights1[23900] <= 16'b0000000000000001;
        weights1[23901] <= 16'b0000000000001110;
        weights1[23902] <= 16'b0000000000000100;
        weights1[23903] <= 16'b1111111111101111;
        weights1[23904] <= 16'b1111111111101111;
        weights1[23905] <= 16'b1111111111111111;
        weights1[23906] <= 16'b1111111111110110;
        weights1[23907] <= 16'b1111111111111100;
        weights1[23908] <= 16'b1111111111110111;
        weights1[23909] <= 16'b1111111111111011;
        weights1[23910] <= 16'b0000000000000011;
        weights1[23911] <= 16'b0000000000000010;
        weights1[23912] <= 16'b1111111111100101;
        weights1[23913] <= 16'b1111111111001110;
        weights1[23914] <= 16'b1111111110110111;
        weights1[23915] <= 16'b1111111110100100;
        weights1[23916] <= 16'b1111111110100011;
        weights1[23917] <= 16'b1111111110000111;
        weights1[23918] <= 16'b1111111110101000;
        weights1[23919] <= 16'b1111111111101000;
        weights1[23920] <= 16'b0000000000100000;
        weights1[23921] <= 16'b1111111111110111;
        weights1[23922] <= 16'b0000000000000100;
        weights1[23923] <= 16'b0000000000000011;
        weights1[23924] <= 16'b0000000000001000;
        weights1[23925] <= 16'b0000000000000101;
        weights1[23926] <= 16'b0000000000010001;
        weights1[23927] <= 16'b0000000000010101;
        weights1[23928] <= 16'b0000000000000100;
        weights1[23929] <= 16'b0000000000001000;
        weights1[23930] <= 16'b1111111111110000;
        weights1[23931] <= 16'b1111111111111000;
        weights1[23932] <= 16'b1111111111111111;
        weights1[23933] <= 16'b1111111111111010;
        weights1[23934] <= 16'b1111111111110011;
        weights1[23935] <= 16'b1111111111111001;
        weights1[23936] <= 16'b0000000000000010;
        weights1[23937] <= 16'b0000000000000011;
        weights1[23938] <= 16'b0000000000001011;
        weights1[23939] <= 16'b0000000000000110;
        weights1[23940] <= 16'b1111111111100010;
        weights1[23941] <= 16'b1111111111001100;
        weights1[23942] <= 16'b1111111110111101;
        weights1[23943] <= 16'b1111111110111010;
        weights1[23944] <= 16'b1111111110110010;
        weights1[23945] <= 16'b1111111111011100;
        weights1[23946] <= 16'b1111111111111011;
        weights1[23947] <= 16'b1111111111110011;
        weights1[23948] <= 16'b1111111111100001;
        weights1[23949] <= 16'b0000000000010011;
        weights1[23950] <= 16'b1111111111110100;
        weights1[23951] <= 16'b0000000000000011;
        weights1[23952] <= 16'b1111111111111101;
        weights1[23953] <= 16'b1111111111111100;
        weights1[23954] <= 16'b0000000000001000;
        weights1[23955] <= 16'b0000000000000010;
        weights1[23956] <= 16'b1111111111110101;
        weights1[23957] <= 16'b1111111111111000;
        weights1[23958] <= 16'b1111111111101111;
        weights1[23959] <= 16'b1111111111101101;
        weights1[23960] <= 16'b1111111111101101;
        weights1[23961] <= 16'b1111111111111011;
        weights1[23962] <= 16'b0000000000001000;
        weights1[23963] <= 16'b0000000000000101;
        weights1[23964] <= 16'b1111111111111000;
        weights1[23965] <= 16'b0000000000001000;
        weights1[23966] <= 16'b0000000000000000;
        weights1[23967] <= 16'b0000000000000001;
        weights1[23968] <= 16'b1111111111101011;
        weights1[23969] <= 16'b1111111111010101;
        weights1[23970] <= 16'b1111111111010011;
        weights1[23971] <= 16'b1111111111011101;
        weights1[23972] <= 16'b1111111111100110;
        weights1[23973] <= 16'b1111111111101111;
        weights1[23974] <= 16'b1111111111111110;
        weights1[23975] <= 16'b1111111111110110;
        weights1[23976] <= 16'b0000000000000001;
        weights1[23977] <= 16'b0000000000010000;
        weights1[23978] <= 16'b1111111111110100;
        weights1[23979] <= 16'b1111111111111100;
        weights1[23980] <= 16'b0000000000000000;
        weights1[23981] <= 16'b0000000000000101;
        weights1[23982] <= 16'b0000000000000010;
        weights1[23983] <= 16'b1111111111101000;
        weights1[23984] <= 16'b1111111111111101;
        weights1[23985] <= 16'b1111111111110110;
        weights1[23986] <= 16'b0000000000000111;
        weights1[23987] <= 16'b0000000000011110;
        weights1[23988] <= 16'b1111111111111100;
        weights1[23989] <= 16'b0000000000000010;
        weights1[23990] <= 16'b1111111111111111;
        weights1[23991] <= 16'b1111111111111000;
        weights1[23992] <= 16'b0000000000010011;
        weights1[23993] <= 16'b0000000000010001;
        weights1[23994] <= 16'b0000000000001110;
        weights1[23995] <= 16'b0000000000000101;
        weights1[23996] <= 16'b1111111111111000;
        weights1[23997] <= 16'b1111111111100011;
        weights1[23998] <= 16'b1111111111101110;
        weights1[23999] <= 16'b1111111111101000;
        weights1[24000] <= 16'b1111111111101110;
        weights1[24001] <= 16'b1111111111110101;
        weights1[24002] <= 16'b1111111111100000;
        weights1[24003] <= 16'b1111111111110101;
        weights1[24004] <= 16'b1111111111101011;
        weights1[24005] <= 16'b1111111111100011;
        weights1[24006] <= 16'b1111111111010010;
        weights1[24007] <= 16'b1111111111111001;
        weights1[24008] <= 16'b1111111111101011;
        weights1[24009] <= 16'b1111111111111001;
        weights1[24010] <= 16'b1111111111111100;
        weights1[24011] <= 16'b1111111111111011;
        weights1[24012] <= 16'b1111111111110000;
        weights1[24013] <= 16'b1111111111110010;
        weights1[24014] <= 16'b1111111111101101;
        weights1[24015] <= 16'b0000000000000001;
        weights1[24016] <= 16'b0000000000000110;
        weights1[24017] <= 16'b0000000000000011;
        weights1[24018] <= 16'b0000000000001011;
        weights1[24019] <= 16'b0000000000011011;
        weights1[24020] <= 16'b0000000000001111;
        weights1[24021] <= 16'b0000000000000011;
        weights1[24022] <= 16'b0000000000000001;
        weights1[24023] <= 16'b1111111111111100;
        weights1[24024] <= 16'b1111111111111111;
        weights1[24025] <= 16'b1111111111111101;
        weights1[24026] <= 16'b1111111111110110;
        weights1[24027] <= 16'b1111111111110110;
        weights1[24028] <= 16'b1111111111101001;
        weights1[24029] <= 16'b0000000000000101;
        weights1[24030] <= 16'b1111111111100110;
        weights1[24031] <= 16'b1111111111111000;
        weights1[24032] <= 16'b1111111111011000;
        weights1[24033] <= 16'b1111111111110011;
        weights1[24034] <= 16'b1111111111010110;
        weights1[24035] <= 16'b1111111111001110;
        weights1[24036] <= 16'b1111111111001111;
        weights1[24037] <= 16'b1111111111111011;
        weights1[24038] <= 16'b1111111111110111;
        weights1[24039] <= 16'b1111111111110010;
        weights1[24040] <= 16'b1111111111100011;
        weights1[24041] <= 16'b1111111111111111;
        weights1[24042] <= 16'b1111111111101111;
        weights1[24043] <= 16'b0000000000001000;
        weights1[24044] <= 16'b1111111111101000;
        weights1[24045] <= 16'b0000000000001111;
        weights1[24046] <= 16'b1111111111110000;
        weights1[24047] <= 16'b1111111111110101;
        weights1[24048] <= 16'b1111111111110111;
        weights1[24049] <= 16'b0000000000010101;
        weights1[24050] <= 16'b0000000000001100;
        weights1[24051] <= 16'b0000000000001000;
        weights1[24052] <= 16'b0000000000010000;
        weights1[24053] <= 16'b0000000000000001;
        weights1[24054] <= 16'b0000000000000100;
        weights1[24055] <= 16'b0000000000011110;
        weights1[24056] <= 16'b1111111111011001;
        weights1[24057] <= 16'b1111111111111001;
        weights1[24058] <= 16'b0000000000001000;
        weights1[24059] <= 16'b1111111111110111;
        weights1[24060] <= 16'b1111111111101100;
        weights1[24061] <= 16'b1111111111111101;
        weights1[24062] <= 16'b1111111111110100;
        weights1[24063] <= 16'b1111111111110000;
        weights1[24064] <= 16'b0000000000000100;
        weights1[24065] <= 16'b0000000000000000;
        weights1[24066] <= 16'b1111111111111100;
        weights1[24067] <= 16'b1111111111110100;
        weights1[24068] <= 16'b0000000000001011;
        weights1[24069] <= 16'b1111111111011111;
        weights1[24070] <= 16'b1111111111101111;
        weights1[24071] <= 16'b1111111111100111;
        weights1[24072] <= 16'b1111111111101111;
        weights1[24073] <= 16'b0000000000001100;
        weights1[24074] <= 16'b0000000000000001;
        weights1[24075] <= 16'b1111111111111111;
        weights1[24076] <= 16'b1111111111111111;
        weights1[24077] <= 16'b0000000000010000;
        weights1[24078] <= 16'b0000000000000100;
        weights1[24079] <= 16'b0000000000001111;
        weights1[24080] <= 16'b0000000000010100;
        weights1[24081] <= 16'b0000000000001100;
        weights1[24082] <= 16'b0000000000001001;
        weights1[24083] <= 16'b0000000000010110;
        weights1[24084] <= 16'b0000000000001101;
        weights1[24085] <= 16'b1111111111101001;
        weights1[24086] <= 16'b0000000000001011;
        weights1[24087] <= 16'b1111111111111111;
        weights1[24088] <= 16'b1111111111111100;
        weights1[24089] <= 16'b0000000000001011;
        weights1[24090] <= 16'b1111111111110101;
        weights1[24091] <= 16'b1111111111111101;
        weights1[24092] <= 16'b0000000000001111;
        weights1[24093] <= 16'b1111111111111101;
        weights1[24094] <= 16'b0000000000001000;
        weights1[24095] <= 16'b1111111111110110;
        weights1[24096] <= 16'b1111111111110111;
        weights1[24097] <= 16'b1111111111101101;
        weights1[24098] <= 16'b0000000000010011;
        weights1[24099] <= 16'b0000000000000100;
        weights1[24100] <= 16'b1111111111110001;
        weights1[24101] <= 16'b0000000000010100;
        weights1[24102] <= 16'b1111111111111010;
        weights1[24103] <= 16'b1111111111111000;
        weights1[24104] <= 16'b0000000000000110;
        weights1[24105] <= 16'b0000000000001000;
        weights1[24106] <= 16'b0000000000000111;
        weights1[24107] <= 16'b0000000000000110;
        weights1[24108] <= 16'b0000000000010100;
        weights1[24109] <= 16'b0000000000001010;
        weights1[24110] <= 16'b0000000000000000;
        weights1[24111] <= 16'b0000000000011000;
        weights1[24112] <= 16'b0000000000001011;
        weights1[24113] <= 16'b1111111111111100;
        weights1[24114] <= 16'b0000000000001011;
        weights1[24115] <= 16'b1111111111100001;
        weights1[24116] <= 16'b0000000000001100;
        weights1[24117] <= 16'b1111111111100111;
        weights1[24118] <= 16'b0000000000001000;
        weights1[24119] <= 16'b0000000000000000;
        weights1[24120] <= 16'b1111111111101101;
        weights1[24121] <= 16'b0000000000000101;
        weights1[24122] <= 16'b0000000000010010;
        weights1[24123] <= 16'b1111111111101110;
        weights1[24124] <= 16'b0000000000010100;
        weights1[24125] <= 16'b1111111111111111;
        weights1[24126] <= 16'b1111111111100111;
        weights1[24127] <= 16'b1111111111101010;
        weights1[24128] <= 16'b0000000000000101;
        weights1[24129] <= 16'b1111111111101111;
        weights1[24130] <= 16'b1111111111100111;
        weights1[24131] <= 16'b0000000000001100;
        weights1[24132] <= 16'b0000000000010010;
        weights1[24133] <= 16'b1111111111110100;
        weights1[24134] <= 16'b1111111111111100;
        weights1[24135] <= 16'b0000000000000100;
        weights1[24136] <= 16'b0000000000000101;
        weights1[24137] <= 16'b0000000000001111;
        weights1[24138] <= 16'b0000000000000111;
        weights1[24139] <= 16'b0000000000000000;
        weights1[24140] <= 16'b0000000000010100;
        weights1[24141] <= 16'b0000000000010000;
        weights1[24142] <= 16'b0000000000010010;
        weights1[24143] <= 16'b0000000000010111;
        weights1[24144] <= 16'b1111111111111000;
        weights1[24145] <= 16'b0000000000100110;
        weights1[24146] <= 16'b0000000000000001;
        weights1[24147] <= 16'b1111111111111011;
        weights1[24148] <= 16'b1111111111110000;
        weights1[24149] <= 16'b1111111111111001;
        weights1[24150] <= 16'b0000000000010100;
        weights1[24151] <= 16'b0000000000001011;
        weights1[24152] <= 16'b0000000000000001;
        weights1[24153] <= 16'b1111111111111110;
        weights1[24154] <= 16'b1111111111111000;
        weights1[24155] <= 16'b1111111111111010;
        weights1[24156] <= 16'b1111111111011011;
        weights1[24157] <= 16'b1111111111100110;
        weights1[24158] <= 16'b1111111111100111;
        weights1[24159] <= 16'b1111111111101110;
        weights1[24160] <= 16'b1111111111111010;
        weights1[24161] <= 16'b1111111111101100;
        weights1[24162] <= 16'b1111111111111101;
        weights1[24163] <= 16'b1111111111111100;
        weights1[24164] <= 16'b0000000000001000;
        weights1[24165] <= 16'b0000000000001101;
        weights1[24166] <= 16'b0000000000001101;
        weights1[24167] <= 16'b0000000000001001;
        weights1[24168] <= 16'b1111111111111111;
        weights1[24169] <= 16'b0000000000000111;
        weights1[24170] <= 16'b1111111111111010;
        weights1[24171] <= 16'b0000000000010001;
        weights1[24172] <= 16'b0000000000011010;
        weights1[24173] <= 16'b0000000000000111;
        weights1[24174] <= 16'b1111111111111000;
        weights1[24175] <= 16'b0000000000001100;
        weights1[24176] <= 16'b0000000000001010;
        weights1[24177] <= 16'b1111111111111100;
        weights1[24178] <= 16'b1111111111111110;
        weights1[24179] <= 16'b1111111111111100;
        weights1[24180] <= 16'b0000000000000000;
        weights1[24181] <= 16'b0000000000000010;
        weights1[24182] <= 16'b1111111111111010;
        weights1[24183] <= 16'b1111111111110101;
        weights1[24184] <= 16'b0000000000000000;
        weights1[24185] <= 16'b1111111111011011;
        weights1[24186] <= 16'b1111111111101101;
        weights1[24187] <= 16'b1111111111110111;
        weights1[24188] <= 16'b1111111111110110;
        weights1[24189] <= 16'b1111111111110110;
        weights1[24190] <= 16'b1111111111111111;
        weights1[24191] <= 16'b1111111111111100;
        weights1[24192] <= 16'b0000000000001000;
        weights1[24193] <= 16'b0000000000010010;
        weights1[24194] <= 16'b0000000000001011;
        weights1[24195] <= 16'b0000000000010010;
        weights1[24196] <= 16'b0000000000001001;
        weights1[24197] <= 16'b0000000000000001;
        weights1[24198] <= 16'b0000000000000001;
        weights1[24199] <= 16'b0000000000010011;
        weights1[24200] <= 16'b0000000000000011;
        weights1[24201] <= 16'b0000000000001110;
        weights1[24202] <= 16'b1111111111111001;
        weights1[24203] <= 16'b0000000000000010;
        weights1[24204] <= 16'b1111111111110000;
        weights1[24205] <= 16'b1111111111101111;
        weights1[24206] <= 16'b0000000000001000;
        weights1[24207] <= 16'b1111111111110001;
        weights1[24208] <= 16'b1111111111100010;
        weights1[24209] <= 16'b1111111111111010;
        weights1[24210] <= 16'b1111111111111000;
        weights1[24211] <= 16'b1111111111110110;
        weights1[24212] <= 16'b1111111111110001;
        weights1[24213] <= 16'b1111111111110100;
        weights1[24214] <= 16'b1111111111110010;
        weights1[24215] <= 16'b1111111111110011;
        weights1[24216] <= 16'b1111111111110001;
        weights1[24217] <= 16'b0000000000000001;
        weights1[24218] <= 16'b1111111111111100;
        weights1[24219] <= 16'b1111111111111011;
        weights1[24220] <= 16'b0000000000001010;
        weights1[24221] <= 16'b0000000000001111;
        weights1[24222] <= 16'b0000000000010000;
        weights1[24223] <= 16'b1111111111111101;
        weights1[24224] <= 16'b0000000000000100;
        weights1[24225] <= 16'b0000000000001011;
        weights1[24226] <= 16'b0000000000010101;
        weights1[24227] <= 16'b0000000000001011;
        weights1[24228] <= 16'b1111111111111110;
        weights1[24229] <= 16'b1111111111101100;
        weights1[24230] <= 16'b1111111111111100;
        weights1[24231] <= 16'b1111111111111100;
        weights1[24232] <= 16'b0000000000001010;
        weights1[24233] <= 16'b1111111111110111;
        weights1[24234] <= 16'b1111111111111011;
        weights1[24235] <= 16'b1111111111100001;
        weights1[24236] <= 16'b0000000000010010;
        weights1[24237] <= 16'b0000000000001110;
        weights1[24238] <= 16'b0000000000001000;
        weights1[24239] <= 16'b0000000000000001;
        weights1[24240] <= 16'b0000000000001110;
        weights1[24241] <= 16'b1111111111111100;
        weights1[24242] <= 16'b0000000000000100;
        weights1[24243] <= 16'b1111111111111001;
        weights1[24244] <= 16'b1111111111111100;
        weights1[24245] <= 16'b0000000000000010;
        weights1[24246] <= 16'b1111111111111101;
        weights1[24247] <= 16'b1111111111111100;
        weights1[24248] <= 16'b0000000000000011;
        weights1[24249] <= 16'b0000000000001001;
        weights1[24250] <= 16'b0000000000010010;
        weights1[24251] <= 16'b0000000000001010;
        weights1[24252] <= 16'b1111111111110111;
        weights1[24253] <= 16'b1111111111110111;
        weights1[24254] <= 16'b0000000000001111;
        weights1[24255] <= 16'b0000000000010011;
        weights1[24256] <= 16'b1111111111110010;
        weights1[24257] <= 16'b1111111111100110;
        weights1[24258] <= 16'b1111111111111100;
        weights1[24259] <= 16'b1111111111111000;
        weights1[24260] <= 16'b1111111111110101;
        weights1[24261] <= 16'b0000000000000111;
        weights1[24262] <= 16'b0000000000000101;
        weights1[24263] <= 16'b0000000000001110;
        weights1[24264] <= 16'b0000000000000001;
        weights1[24265] <= 16'b1111111111111110;
        weights1[24266] <= 16'b0000000000000111;
        weights1[24267] <= 16'b0000000000000110;
        weights1[24268] <= 16'b0000000000001010;
        weights1[24269] <= 16'b0000000000000100;
        weights1[24270] <= 16'b0000000000000000;
        weights1[24271] <= 16'b1111111111111011;
        weights1[24272] <= 16'b1111111111111101;
        weights1[24273] <= 16'b0000000000000001;
        weights1[24274] <= 16'b1111111111111111;
        weights1[24275] <= 16'b1111111111111111;
        weights1[24276] <= 16'b0000000000000010;
        weights1[24277] <= 16'b0000000000000111;
        weights1[24278] <= 16'b0000000000001011;
        weights1[24279] <= 16'b0000000000011000;
        weights1[24280] <= 16'b0000000000010100;
        weights1[24281] <= 16'b0000000000011010;
        weights1[24282] <= 16'b0000000000100000;
        weights1[24283] <= 16'b0000000000010110;
        weights1[24284] <= 16'b0000000000010010;
        weights1[24285] <= 16'b0000000000001100;
        weights1[24286] <= 16'b0000000000000111;
        weights1[24287] <= 16'b0000000000000110;
        weights1[24288] <= 16'b0000000000001100;
        weights1[24289] <= 16'b0000000000000011;
        weights1[24290] <= 16'b1111111111110011;
        weights1[24291] <= 16'b0000000000001101;
        weights1[24292] <= 16'b0000000000010011;
        weights1[24293] <= 16'b1111111111111001;
        weights1[24294] <= 16'b1111111111111010;
        weights1[24295] <= 16'b0000000000010101;
        weights1[24296] <= 16'b0000000000001110;
        weights1[24297] <= 16'b0000000000000001;
        weights1[24298] <= 16'b1111111111111110;
        weights1[24299] <= 16'b0000000000000011;
        weights1[24300] <= 16'b0000000000000001;
        weights1[24301] <= 16'b0000000000000001;
        weights1[24302] <= 16'b0000000000000001;
        weights1[24303] <= 16'b0000000000000000;
        weights1[24304] <= 16'b0000000000000001;
        weights1[24305] <= 16'b0000000000000001;
        weights1[24306] <= 16'b0000000000000000;
        weights1[24307] <= 16'b1111111111111100;
        weights1[24308] <= 16'b0000000000000000;
        weights1[24309] <= 16'b1111111111111000;
        weights1[24310] <= 16'b1111111111110111;
        weights1[24311] <= 16'b1111111111111000;
        weights1[24312] <= 16'b1111111111111000;
        weights1[24313] <= 16'b1111111111110111;
        weights1[24314] <= 16'b1111111111111010;
        weights1[24315] <= 16'b0000000000000011;
        weights1[24316] <= 16'b1111111111111110;
        weights1[24317] <= 16'b1111111111110101;
        weights1[24318] <= 16'b1111111111111000;
        weights1[24319] <= 16'b1111111111101001;
        weights1[24320] <= 16'b1111111111110011;
        weights1[24321] <= 16'b1111111111110101;
        weights1[24322] <= 16'b1111111111111101;
        weights1[24323] <= 16'b1111111111101011;
        weights1[24324] <= 16'b1111111111110011;
        weights1[24325] <= 16'b1111111111111001;
        weights1[24326] <= 16'b1111111111111110;
        weights1[24327] <= 16'b0000000000000101;
        weights1[24328] <= 16'b0000000000000110;
        weights1[24329] <= 16'b0000000000000100;
        weights1[24330] <= 16'b0000000000000101;
        weights1[24331] <= 16'b0000000000000001;
        weights1[24332] <= 16'b0000000000000000;
        weights1[24333] <= 16'b1111111111111111;
        weights1[24334] <= 16'b1111111111111011;
        weights1[24335] <= 16'b1111111111111100;
        weights1[24336] <= 16'b1111111111111011;
        weights1[24337] <= 16'b1111111111110111;
        weights1[24338] <= 16'b1111111111110000;
        weights1[24339] <= 16'b1111111111101011;
        weights1[24340] <= 16'b1111111111111100;
        weights1[24341] <= 16'b1111111111111010;
        weights1[24342] <= 16'b0000000000000001;
        weights1[24343] <= 16'b0000000000001001;
        weights1[24344] <= 16'b1111111111111000;
        weights1[24345] <= 16'b1111111111111111;
        weights1[24346] <= 16'b1111111111111011;
        weights1[24347] <= 16'b1111111111110110;
        weights1[24348] <= 16'b1111111111110110;
        weights1[24349] <= 16'b1111111111111000;
        weights1[24350] <= 16'b1111111111111010;
        weights1[24351] <= 16'b1111111111110100;
        weights1[24352] <= 16'b0000000000000000;
        weights1[24353] <= 16'b0000000000000011;
        weights1[24354] <= 16'b0000000000000111;
        weights1[24355] <= 16'b0000000000000000;
        weights1[24356] <= 16'b1111111111111111;
        weights1[24357] <= 16'b0000000000000101;
        weights1[24358] <= 16'b0000000000000011;
        weights1[24359] <= 16'b0000000000000011;
        weights1[24360] <= 16'b0000000000000000;
        weights1[24361] <= 16'b1111111111111111;
        weights1[24362] <= 16'b1111111111110111;
        weights1[24363] <= 16'b1111111111111100;
        weights1[24364] <= 16'b1111111111111011;
        weights1[24365] <= 16'b1111111111110011;
        weights1[24366] <= 16'b1111111111110110;
        weights1[24367] <= 16'b1111111111101101;
        weights1[24368] <= 16'b1111111111111000;
        weights1[24369] <= 16'b1111111111111000;
        weights1[24370] <= 16'b0000000000000011;
        weights1[24371] <= 16'b1111111111111100;
        weights1[24372] <= 16'b1111111111111001;
        weights1[24373] <= 16'b0000000000000010;
        weights1[24374] <= 16'b0000000000000100;
        weights1[24375] <= 16'b1111111111111001;
        weights1[24376] <= 16'b1111111111110010;
        weights1[24377] <= 16'b1111111111111010;
        weights1[24378] <= 16'b1111111111110111;
        weights1[24379] <= 16'b1111111111110011;
        weights1[24380] <= 16'b1111111111111101;
        weights1[24381] <= 16'b0000000000000100;
        weights1[24382] <= 16'b0000000000001100;
        weights1[24383] <= 16'b0000000000000001;
        weights1[24384] <= 16'b1111111111111101;
        weights1[24385] <= 16'b1111111111111000;
        weights1[24386] <= 16'b0000000000000001;
        weights1[24387] <= 16'b1111111111111111;
        weights1[24388] <= 16'b0000000000000000;
        weights1[24389] <= 16'b1111111111111100;
        weights1[24390] <= 16'b1111111111111011;
        weights1[24391] <= 16'b1111111111111001;
        weights1[24392] <= 16'b1111111111111101;
        weights1[24393] <= 16'b1111111111111101;
        weights1[24394] <= 16'b0000000000000111;
        weights1[24395] <= 16'b1111111111110000;
        weights1[24396] <= 16'b0000000000001010;
        weights1[24397] <= 16'b1111111111101011;
        weights1[24398] <= 16'b1111111111110011;
        weights1[24399] <= 16'b1111111111110001;
        weights1[24400] <= 16'b0000000000000010;
        weights1[24401] <= 16'b1111111111110110;
        weights1[24402] <= 16'b0000000000001111;
        weights1[24403] <= 16'b0000000000001000;
        weights1[24404] <= 16'b0000000000000001;
        weights1[24405] <= 16'b1111111111110010;
        weights1[24406] <= 16'b1111111111111001;
        weights1[24407] <= 16'b1111111111111100;
        weights1[24408] <= 16'b0000000000001001;
        weights1[24409] <= 16'b0000000000010000;
        weights1[24410] <= 16'b1111111111111101;
        weights1[24411] <= 16'b1111111111111000;
        weights1[24412] <= 16'b0000000000001000;
        weights1[24413] <= 16'b0000000000000000;
        weights1[24414] <= 16'b0000000000000100;
        weights1[24415] <= 16'b1111111111111011;
        weights1[24416] <= 16'b1111111111111111;
        weights1[24417] <= 16'b1111111111111111;
        weights1[24418] <= 16'b0000000000000010;
        weights1[24419] <= 16'b1111111111111101;
        weights1[24420] <= 16'b1111111111111010;
        weights1[24421] <= 16'b1111111111110110;
        weights1[24422] <= 16'b0000000000001111;
        weights1[24423] <= 16'b1111111111101111;
        weights1[24424] <= 16'b0000000000001010;
        weights1[24425] <= 16'b1111111111111001;
        weights1[24426] <= 16'b1111111111111000;
        weights1[24427] <= 16'b1111111111111000;
        weights1[24428] <= 16'b0000000000000011;
        weights1[24429] <= 16'b1111111111110101;
        weights1[24430] <= 16'b0000000000000010;
        weights1[24431] <= 16'b0000000000000011;
        weights1[24432] <= 16'b1111111111111111;
        weights1[24433] <= 16'b0000000000010011;
        weights1[24434] <= 16'b1111111111111001;
        weights1[24435] <= 16'b1111111111101110;
        weights1[24436] <= 16'b1111111111111111;
        weights1[24437] <= 16'b0000000000001110;
        weights1[24438] <= 16'b1111111111110111;
        weights1[24439] <= 16'b0000000000000001;
        weights1[24440] <= 16'b0000000000010011;
        weights1[24441] <= 16'b0000000000010101;
        weights1[24442] <= 16'b1111111111111101;
        weights1[24443] <= 16'b0000000000000111;
        weights1[24444] <= 16'b1111111111111101;
        weights1[24445] <= 16'b0000000000000010;
        weights1[24446] <= 16'b0000000000000101;
        weights1[24447] <= 16'b1111111111110111;
        weights1[24448] <= 16'b1111111111111110;
        weights1[24449] <= 16'b1111111111111011;
        weights1[24450] <= 16'b1111111111110101;
        weights1[24451] <= 16'b0000000000001001;
        weights1[24452] <= 16'b1111111111111111;
        weights1[24453] <= 16'b0000000000001010;
        weights1[24454] <= 16'b0000000000000111;
        weights1[24455] <= 16'b0000000000000100;
        weights1[24456] <= 16'b0000000000001100;
        weights1[24457] <= 16'b1111111111111101;
        weights1[24458] <= 16'b0000000000000010;
        weights1[24459] <= 16'b1111111111111111;
        weights1[24460] <= 16'b0000000000000000;
        weights1[24461] <= 16'b0000000000000010;
        weights1[24462] <= 16'b1111111111110000;
        weights1[24463] <= 16'b1111111111111011;
        weights1[24464] <= 16'b0000000000000001;
        weights1[24465] <= 16'b0000000000000011;
        weights1[24466] <= 16'b0000000000000111;
        weights1[24467] <= 16'b0000000000000011;
        weights1[24468] <= 16'b0000000000001011;
        weights1[24469] <= 16'b1111111111110101;
        weights1[24470] <= 16'b1111111111111011;
        weights1[24471] <= 16'b1111111111111010;
        weights1[24472] <= 16'b0000000000000010;
        weights1[24473] <= 16'b0000000000000001;
        weights1[24474] <= 16'b1111111111111010;
        weights1[24475] <= 16'b1111111111111101;
        weights1[24476] <= 16'b0000000000001011;
        weights1[24477] <= 16'b0000000000000101;
        weights1[24478] <= 16'b1111111111111101;
        weights1[24479] <= 16'b1111111111011110;
        weights1[24480] <= 16'b1111111111111101;
        weights1[24481] <= 16'b1111111111110101;
        weights1[24482] <= 16'b1111111111111100;
        weights1[24483] <= 16'b1111111111100000;
        weights1[24484] <= 16'b0000000000000101;
        weights1[24485] <= 16'b0000000000000111;
        weights1[24486] <= 16'b0000000000000011;
        weights1[24487] <= 16'b0000000000001010;
        weights1[24488] <= 16'b1111111111111111;
        weights1[24489] <= 16'b1111111111110000;
        weights1[24490] <= 16'b1111111111111000;
        weights1[24491] <= 16'b1111111111110010;
        weights1[24492] <= 16'b1111111111110000;
        weights1[24493] <= 16'b0000000000000111;
        weights1[24494] <= 16'b1111111111101101;
        weights1[24495] <= 16'b1111111111111100;
        weights1[24496] <= 16'b0000000000001011;
        weights1[24497] <= 16'b0000000000001011;
        weights1[24498] <= 16'b0000000000000100;
        weights1[24499] <= 16'b1111111111111110;
        weights1[24500] <= 16'b0000000000000000;
        weights1[24501] <= 16'b0000000000000111;
        weights1[24502] <= 16'b0000000000000100;
        weights1[24503] <= 16'b0000000000000111;
        weights1[24504] <= 16'b1111111111111110;
        weights1[24505] <= 16'b0000000000000101;
        weights1[24506] <= 16'b0000000000001011;
        weights1[24507] <= 16'b0000000000000110;
        weights1[24508] <= 16'b1111111111110001;
        weights1[24509] <= 16'b0000000000000100;
        weights1[24510] <= 16'b1111111111110111;
        weights1[24511] <= 16'b0000000000001000;
        weights1[24512] <= 16'b1111111111110001;
        weights1[24513] <= 16'b1111111111110111;
        weights1[24514] <= 16'b1111111111110110;
        weights1[24515] <= 16'b1111111111110000;
        weights1[24516] <= 16'b1111111111110111;
        weights1[24517] <= 16'b1111111111111111;
        weights1[24518] <= 16'b1111111111111001;
        weights1[24519] <= 16'b0000000000000001;
        weights1[24520] <= 16'b1111111111110110;
        weights1[24521] <= 16'b0000000000001001;
        weights1[24522] <= 16'b1111111111111001;
        weights1[24523] <= 16'b0000000000010101;
        weights1[24524] <= 16'b0000000000000010;
        weights1[24525] <= 16'b1111111111111101;
        weights1[24526] <= 16'b1111111111111001;
        weights1[24527] <= 16'b1111111111111110;
        weights1[24528] <= 16'b0000000000001010;
        weights1[24529] <= 16'b0000000000000000;
        weights1[24530] <= 16'b0000000000001001;
        weights1[24531] <= 16'b0000000000001000;
        weights1[24532] <= 16'b0000000000001001;
        weights1[24533] <= 16'b0000000000000100;
        weights1[24534] <= 16'b0000000000001100;
        weights1[24535] <= 16'b0000000000000000;
        weights1[24536] <= 16'b0000000000010010;
        weights1[24537] <= 16'b1111111111111001;
        weights1[24538] <= 16'b0000000000000101;
        weights1[24539] <= 16'b1111111111111010;
        weights1[24540] <= 16'b0000000000001000;
        weights1[24541] <= 16'b1111111111111001;
        weights1[24542] <= 16'b0000000000001110;
        weights1[24543] <= 16'b1111111111111101;
        weights1[24544] <= 16'b1111111111111110;
        weights1[24545] <= 16'b0000000000010010;
        weights1[24546] <= 16'b1111111111110101;
        weights1[24547] <= 16'b1111111111111100;
        weights1[24548] <= 16'b1111111111111011;
        weights1[24549] <= 16'b0000000000001100;
        weights1[24550] <= 16'b1111111111110011;
        weights1[24551] <= 16'b1111111111110110;
        weights1[24552] <= 16'b0000000000000011;
        weights1[24553] <= 16'b0000000000001001;
        weights1[24554] <= 16'b1111111111110110;
        weights1[24555] <= 16'b1111111111110110;
        weights1[24556] <= 16'b0000000000000011;
        weights1[24557] <= 16'b0000000000000110;
        weights1[24558] <= 16'b0000000000001101;
        weights1[24559] <= 16'b1111111111111100;
        weights1[24560] <= 16'b0000000000001111;
        weights1[24561] <= 16'b0000000000001001;
        weights1[24562] <= 16'b1111111111111101;
        weights1[24563] <= 16'b0000000000001011;
        weights1[24564] <= 16'b1111111111111010;
        weights1[24565] <= 16'b0000000000000110;
        weights1[24566] <= 16'b0000000000001111;
        weights1[24567] <= 16'b1111111111111000;
        weights1[24568] <= 16'b1111111111110100;
        weights1[24569] <= 16'b1111111111110111;
        weights1[24570] <= 16'b0000000000000000;
        weights1[24571] <= 16'b0000000000000000;
        weights1[24572] <= 16'b1111111111111101;
        weights1[24573] <= 16'b1111111111111011;
        weights1[24574] <= 16'b0000000000000110;
        weights1[24575] <= 16'b0000000000000011;
        weights1[24576] <= 16'b1111111111111110;
        weights1[24577] <= 16'b0000000000010101;
        weights1[24578] <= 16'b0000000000001011;
        weights1[24579] <= 16'b0000000000000101;
        weights1[24580] <= 16'b1111111111110110;
        weights1[24581] <= 16'b0000000000000001;
        weights1[24582] <= 16'b1111111111101000;
        weights1[24583] <= 16'b1111111111110000;
        weights1[24584] <= 16'b0000000000000010;
        weights1[24585] <= 16'b1111111111110011;
        weights1[24586] <= 16'b1111111111111001;
        weights1[24587] <= 16'b1111111111110110;
        weights1[24588] <= 16'b1111111111101011;
        weights1[24589] <= 16'b1111111111111110;
        weights1[24590] <= 16'b1111111111110110;
        weights1[24591] <= 16'b1111111111111001;
        weights1[24592] <= 16'b1111111111111111;
        weights1[24593] <= 16'b1111111111111100;
        weights1[24594] <= 16'b1111111111110011;
        weights1[24595] <= 16'b1111111111111010;
        weights1[24596] <= 16'b0000000000001001;
        weights1[24597] <= 16'b0000000000010011;
        weights1[24598] <= 16'b1111111111110010;
        weights1[24599] <= 16'b0000000000000100;
        weights1[24600] <= 16'b1111111111111101;
        weights1[24601] <= 16'b0000000000000101;
        weights1[24602] <= 16'b0000000000000110;
        weights1[24603] <= 16'b0000000000000010;
        weights1[24604] <= 16'b1111111111110010;
        weights1[24605] <= 16'b0000000000000000;
        weights1[24606] <= 16'b1111111111110111;
        weights1[24607] <= 16'b0000000000000111;
        weights1[24608] <= 16'b1111111111111101;
        weights1[24609] <= 16'b1111111111111110;
        weights1[24610] <= 16'b1111111111101011;
        weights1[24611] <= 16'b1111111111110100;
        weights1[24612] <= 16'b0000000000001001;
        weights1[24613] <= 16'b0000000000000110;
        weights1[24614] <= 16'b0000000000000100;
        weights1[24615] <= 16'b0000000000000011;
        weights1[24616] <= 16'b0000000000001100;
        weights1[24617] <= 16'b0000000000001100;
        weights1[24618] <= 16'b0000000000000010;
        weights1[24619] <= 16'b0000000000000010;
        weights1[24620] <= 16'b1111111111101011;
        weights1[24621] <= 16'b0000000000001111;
        weights1[24622] <= 16'b0000000000010111;
        weights1[24623] <= 16'b1111111111101101;
        weights1[24624] <= 16'b1111111111111010;
        weights1[24625] <= 16'b0000000000000001;
        weights1[24626] <= 16'b1111111111111001;
        weights1[24627] <= 16'b1111111111110111;
        weights1[24628] <= 16'b1111111111110110;
        weights1[24629] <= 16'b1111111111111111;
        weights1[24630] <= 16'b1111111111111100;
        weights1[24631] <= 16'b1111111111111011;
        weights1[24632] <= 16'b1111111111110110;
        weights1[24633] <= 16'b0000000000001101;
        weights1[24634] <= 16'b1111111111111111;
        weights1[24635] <= 16'b1111111111111001;
        weights1[24636] <= 16'b0000000000000010;
        weights1[24637] <= 16'b1111111111111110;
        weights1[24638] <= 16'b0000000000000011;
        weights1[24639] <= 16'b0000000000000010;
        weights1[24640] <= 16'b0000000000001001;
        weights1[24641] <= 16'b0000000000001010;
        weights1[24642] <= 16'b0000000000010111;
        weights1[24643] <= 16'b0000000000001010;
        weights1[24644] <= 16'b0000000000000111;
        weights1[24645] <= 16'b0000000000010001;
        weights1[24646] <= 16'b0000000000010011;
        weights1[24647] <= 16'b0000000000010000;
        weights1[24648] <= 16'b0000000000010100;
        weights1[24649] <= 16'b0000000000000110;
        weights1[24650] <= 16'b1111111111111000;
        weights1[24651] <= 16'b0000000000001011;
        weights1[24652] <= 16'b0000000000001010;
        weights1[24653] <= 16'b1111111111111100;
        weights1[24654] <= 16'b1111111111110100;
        weights1[24655] <= 16'b0000000000001101;
        weights1[24656] <= 16'b0000000000001110;
        weights1[24657] <= 16'b1111111111111110;
        weights1[24658] <= 16'b1111111111110101;
        weights1[24659] <= 16'b0000000000010001;
        weights1[24660] <= 16'b0000000000000011;
        weights1[24661] <= 16'b0000000000001001;
        weights1[24662] <= 16'b0000000000010100;
        weights1[24663] <= 16'b1111111111111101;
        weights1[24664] <= 16'b0000000000001100;
        weights1[24665] <= 16'b0000000000000011;
        weights1[24666] <= 16'b1111111111111000;
        weights1[24667] <= 16'b0000000000000101;
        weights1[24668] <= 16'b0000000000000011;
        weights1[24669] <= 16'b0000000000000101;
        weights1[24670] <= 16'b0000000000011010;
        weights1[24671] <= 16'b0000000000001001;
        weights1[24672] <= 16'b0000000000000101;
        weights1[24673] <= 16'b0000000000100110;
        weights1[24674] <= 16'b1111111111111000;
        weights1[24675] <= 16'b0000000000010001;
        weights1[24676] <= 16'b0000000000001100;
        weights1[24677] <= 16'b0000000000001110;
        weights1[24678] <= 16'b0000000000001011;
        weights1[24679] <= 16'b1111111111110010;
        weights1[24680] <= 16'b0000000000000001;
        weights1[24681] <= 16'b1111111111110010;
        weights1[24682] <= 16'b1111111111111011;
        weights1[24683] <= 16'b0000000000000101;
        weights1[24684] <= 16'b1111111111111100;
        weights1[24685] <= 16'b0000000000010011;
        weights1[24686] <= 16'b0000000000010001;
        weights1[24687] <= 16'b1111111111110011;
        weights1[24688] <= 16'b0000000000000000;
        weights1[24689] <= 16'b0000000000000101;
        weights1[24690] <= 16'b1111111111111100;
        weights1[24691] <= 16'b1111111111110111;
        weights1[24692] <= 16'b0000000000000000;
        weights1[24693] <= 16'b0000000000000011;
        weights1[24694] <= 16'b1111111111111011;
        weights1[24695] <= 16'b0000000000000011;
        weights1[24696] <= 16'b1111111111111101;
        weights1[24697] <= 16'b0000000000010010;
        weights1[24698] <= 16'b0000000000001101;
        weights1[24699] <= 16'b0000000000001001;
        weights1[24700] <= 16'b0000000000001001;
        weights1[24701] <= 16'b0000000000000010;
        weights1[24702] <= 16'b0000000000001110;
        weights1[24703] <= 16'b0000000000000101;
        weights1[24704] <= 16'b0000000000000100;
        weights1[24705] <= 16'b1111111111111101;
        weights1[24706] <= 16'b0000000000000010;
        weights1[24707] <= 16'b0000000000001011;
        weights1[24708] <= 16'b0000000000000100;
        weights1[24709] <= 16'b1111111111111111;
        weights1[24710] <= 16'b1111111111111110;
        weights1[24711] <= 16'b1111111111110110;
        weights1[24712] <= 16'b0000000000000101;
        weights1[24713] <= 16'b0000000000001101;
        weights1[24714] <= 16'b0000000000000001;
        weights1[24715] <= 16'b0000000000000101;
        weights1[24716] <= 16'b1111111111111000;
        weights1[24717] <= 16'b1111111111111010;
        weights1[24718] <= 16'b1111111111110101;
        weights1[24719] <= 16'b0000000000000110;
        weights1[24720] <= 16'b0000000000001100;
        weights1[24721] <= 16'b0000000000000000;
        weights1[24722] <= 16'b1111111111110000;
        weights1[24723] <= 16'b0000000000000101;
        weights1[24724] <= 16'b0000000000001101;
        weights1[24725] <= 16'b0000000000001011;
        weights1[24726] <= 16'b0000000000001001;
        weights1[24727] <= 16'b0000000000001011;
        weights1[24728] <= 16'b1111111111111010;
        weights1[24729] <= 16'b1111111111101100;
        weights1[24730] <= 16'b0000000000000000;
        weights1[24731] <= 16'b1111111111101101;
        weights1[24732] <= 16'b0000000000000111;
        weights1[24733] <= 16'b1111111111101101;
        weights1[24734] <= 16'b1111111111111101;
        weights1[24735] <= 16'b0000000000000001;
        weights1[24736] <= 16'b1111111111101101;
        weights1[24737] <= 16'b1111111111110010;
        weights1[24738] <= 16'b1111111111100101;
        weights1[24739] <= 16'b1111111111101101;
        weights1[24740] <= 16'b0000000000001011;
        weights1[24741] <= 16'b1111111111111100;
        weights1[24742] <= 16'b0000000000001100;
        weights1[24743] <= 16'b0000000000001000;
        weights1[24744] <= 16'b1111111111111101;
        weights1[24745] <= 16'b0000000000001100;
        weights1[24746] <= 16'b0000000000000110;
        weights1[24747] <= 16'b0000000000001000;
        weights1[24748] <= 16'b0000000000001011;
        weights1[24749] <= 16'b1111111111111001;
        weights1[24750] <= 16'b0000000000000111;
        weights1[24751] <= 16'b1111111111111110;
        weights1[24752] <= 16'b0000000000001111;
        weights1[24753] <= 16'b0000000000001011;
        weights1[24754] <= 16'b0000000000001110;
        weights1[24755] <= 16'b0000000000000111;
        weights1[24756] <= 16'b0000000000001101;
        weights1[24757] <= 16'b1111111111110101;
        weights1[24758] <= 16'b1111111111110111;
        weights1[24759] <= 16'b1111111111101110;
        weights1[24760] <= 16'b0000000000000110;
        weights1[24761] <= 16'b0000000000000010;
        weights1[24762] <= 16'b0000000000000001;
        weights1[24763] <= 16'b0000000000010010;
        weights1[24764] <= 16'b0000000000000010;
        weights1[24765] <= 16'b1111111111101101;
        weights1[24766] <= 16'b1111111111011110;
        weights1[24767] <= 16'b1111111111100111;
        weights1[24768] <= 16'b0000000000000001;
        weights1[24769] <= 16'b0000000000001110;
        weights1[24770] <= 16'b0000000000001101;
        weights1[24771] <= 16'b0000000000001011;
        weights1[24772] <= 16'b1111111111111100;
        weights1[24773] <= 16'b0000000000000011;
        weights1[24774] <= 16'b1111111111110111;
        weights1[24775] <= 16'b0000000000001001;
        weights1[24776] <= 16'b0000000000010000;
        weights1[24777] <= 16'b0000000000010101;
        weights1[24778] <= 16'b0000000000000110;
        weights1[24779] <= 16'b0000000000000011;
        weights1[24780] <= 16'b0000000000000010;
        weights1[24781] <= 16'b1111111111111001;
        weights1[24782] <= 16'b0000000000000110;
        weights1[24783] <= 16'b1111111111100111;
        weights1[24784] <= 16'b0000000000000100;
        weights1[24785] <= 16'b1111111111101101;
        weights1[24786] <= 16'b1111111111100011;
        weights1[24787] <= 16'b1111111111110000;
        weights1[24788] <= 16'b1111111111101100;
        weights1[24789] <= 16'b0000000000000010;
        weights1[24790] <= 16'b0000000000100001;
        weights1[24791] <= 16'b0000000000001100;
        weights1[24792] <= 16'b1111111111110000;
        weights1[24793] <= 16'b1111111111101010;
        weights1[24794] <= 16'b1111111111101000;
        weights1[24795] <= 16'b1111111111101100;
        weights1[24796] <= 16'b0000000000010000;
        weights1[24797] <= 16'b0000000000011101;
        weights1[24798] <= 16'b0000000000000101;
        weights1[24799] <= 16'b0000000000001000;
        weights1[24800] <= 16'b1111111111110101;
        weights1[24801] <= 16'b0000000000000001;
        weights1[24802] <= 16'b1111111111111110;
        weights1[24803] <= 16'b0000000000000000;
        weights1[24804] <= 16'b0000000000011011;
        weights1[24805] <= 16'b0000000000000111;
        weights1[24806] <= 16'b0000000000001010;
        weights1[24807] <= 16'b0000000000000011;
        weights1[24808] <= 16'b1111111111111010;
        weights1[24809] <= 16'b1111111111101110;
        weights1[24810] <= 16'b1111111111110100;
        weights1[24811] <= 16'b1111111111101011;
        weights1[24812] <= 16'b1111111111110001;
        weights1[24813] <= 16'b1111111111100100;
        weights1[24814] <= 16'b1111111111010011;
        weights1[24815] <= 16'b1111111111101100;
        weights1[24816] <= 16'b0000000000100000;
        weights1[24817] <= 16'b0000000000100100;
        weights1[24818] <= 16'b0000000000101000;
        weights1[24819] <= 16'b0000000000010110;
        weights1[24820] <= 16'b1111111111110110;
        weights1[24821] <= 16'b1111111111100011;
        weights1[24822] <= 16'b1111111111000000;
        weights1[24823] <= 16'b1111111111011011;
        weights1[24824] <= 16'b0000000000101000;
        weights1[24825] <= 16'b0000000000101010;
        weights1[24826] <= 16'b0000000000010101;
        weights1[24827] <= 16'b1111111111111101;
        weights1[24828] <= 16'b1111111111111011;
        weights1[24829] <= 16'b1111111111100111;
        weights1[24830] <= 16'b0000000000000100;
        weights1[24831] <= 16'b0000000000010100;
        weights1[24832] <= 16'b0000000000010110;
        weights1[24833] <= 16'b0000000000001100;
        weights1[24834] <= 16'b0000000000001010;
        weights1[24835] <= 16'b0000000000001000;
        weights1[24836] <= 16'b1111111111110010;
        weights1[24837] <= 16'b1111111111101001;
        weights1[24838] <= 16'b1111111111100100;
        weights1[24839] <= 16'b1111111111010000;
        weights1[24840] <= 16'b1111111111000101;
        weights1[24841] <= 16'b1111111111100100;
        weights1[24842] <= 16'b1111111111110011;
        weights1[24843] <= 16'b1111111111111100;
        weights1[24844] <= 16'b0000000000110100;
        weights1[24845] <= 16'b0000000000011011;
        weights1[24846] <= 16'b0000000000010001;
        weights1[24847] <= 16'b0000000000000000;
        weights1[24848] <= 16'b1111111111101101;
        weights1[24849] <= 16'b1111111111010001;
        weights1[24850] <= 16'b1111111110100010;
        weights1[24851] <= 16'b1111111111101100;
        weights1[24852] <= 16'b0000000000101101;
        weights1[24853] <= 16'b0000000000010111;
        weights1[24854] <= 16'b0000000000010011;
        weights1[24855] <= 16'b0000000000001000;
        weights1[24856] <= 16'b1111111111100000;
        weights1[24857] <= 16'b1111111111010110;
        weights1[24858] <= 16'b1111111111111000;
        weights1[24859] <= 16'b1111111111111010;
        weights1[24860] <= 16'b0000000000001101;
        weights1[24861] <= 16'b0000000000010111;
        weights1[24862] <= 16'b0000000000001101;
        weights1[24863] <= 16'b0000000000001111;
        weights1[24864] <= 16'b1111111111101101;
        weights1[24865] <= 16'b1111111111100101;
        weights1[24866] <= 16'b1111111111011111;
        weights1[24867] <= 16'b1111111111001000;
        weights1[24868] <= 16'b1111111111001000;
        weights1[24869] <= 16'b1111111111011101;
        weights1[24870] <= 16'b1111111111110111;
        weights1[24871] <= 16'b0000000000101000;
        weights1[24872] <= 16'b0000000000110101;
        weights1[24873] <= 16'b0000000000010001;
        weights1[24874] <= 16'b0000000000010011;
        weights1[24875] <= 16'b1111111111100001;
        weights1[24876] <= 16'b1111111111011010;
        weights1[24877] <= 16'b1111111110011011;
        weights1[24878] <= 16'b1111111110110111;
        weights1[24879] <= 16'b0000000000001010;
        weights1[24880] <= 16'b0000000000111010;
        weights1[24881] <= 16'b0000000000100000;
        weights1[24882] <= 16'b0000000000000101;
        weights1[24883] <= 16'b0000000000010011;
        weights1[24884] <= 16'b1111111111101101;
        weights1[24885] <= 16'b1111111111001100;
        weights1[24886] <= 16'b1111111111001000;
        weights1[24887] <= 16'b1111111111101001;
        weights1[24888] <= 16'b0000000000000010;
        weights1[24889] <= 16'b0000000000010000;
        weights1[24890] <= 16'b0000000000010001;
        weights1[24891] <= 16'b0000000000000110;
        weights1[24892] <= 16'b1111111111101001;
        weights1[24893] <= 16'b1111111111011100;
        weights1[24894] <= 16'b1111111111001100;
        weights1[24895] <= 16'b1111111111011011;
        weights1[24896] <= 16'b1111111111101000;
        weights1[24897] <= 16'b0000000000000111;
        weights1[24898] <= 16'b0000000000001110;
        weights1[24899] <= 16'b0000000000101101;
        weights1[24900] <= 16'b0000000001010101;
        weights1[24901] <= 16'b0000000000010111;
        weights1[24902] <= 16'b0000000000011000;
        weights1[24903] <= 16'b1111111111001101;
        weights1[24904] <= 16'b1111111110110100;
        weights1[24905] <= 16'b1111111101111100;
        weights1[24906] <= 16'b1111111111000101;
        weights1[24907] <= 16'b0000000000100111;
        weights1[24908] <= 16'b0000000000111110;
        weights1[24909] <= 16'b0000000000100001;
        weights1[24910] <= 16'b0000000000001001;
        weights1[24911] <= 16'b1111111111111110;
        weights1[24912] <= 16'b1111111111111001;
        weights1[24913] <= 16'b1111111111010001;
        weights1[24914] <= 16'b1111111110111001;
        weights1[24915] <= 16'b1111111111100111;
        weights1[24916] <= 16'b1111111111110100;
        weights1[24917] <= 16'b0000000000000110;
        weights1[24918] <= 16'b0000000000010000;
        weights1[24919] <= 16'b0000000000001000;
        weights1[24920] <= 16'b1111111111101100;
        weights1[24921] <= 16'b1111111111100011;
        weights1[24922] <= 16'b1111111111110010;
        weights1[24923] <= 16'b1111111111110111;
        weights1[24924] <= 16'b1111111111111111;
        weights1[24925] <= 16'b0000000000101000;
        weights1[24926] <= 16'b0000000001000000;
        weights1[24927] <= 16'b0000000001001001;
        weights1[24928] <= 16'b0000000000100111;
        weights1[24929] <= 16'b0000000000000000;
        weights1[24930] <= 16'b1111111111000000;
        weights1[24931] <= 16'b1111111110011110;
        weights1[24932] <= 16'b1111111110001101;
        weights1[24933] <= 16'b1111111101110101;
        weights1[24934] <= 16'b1111111111100011;
        weights1[24935] <= 16'b0000000000110000;
        weights1[24936] <= 16'b0000000000101101;
        weights1[24937] <= 16'b0000000000101001;
        weights1[24938] <= 16'b0000000000101111;
        weights1[24939] <= 16'b0000000000010000;
        weights1[24940] <= 16'b0000000000000010;
        weights1[24941] <= 16'b1111111111000000;
        weights1[24942] <= 16'b1111111110011011;
        weights1[24943] <= 16'b1111111110111101;
        weights1[24944] <= 16'b1111111111011111;
        weights1[24945] <= 16'b1111111111111110;
        weights1[24946] <= 16'b0000000000000100;
        weights1[24947] <= 16'b0000000000000011;
        weights1[24948] <= 16'b1111111111101101;
        weights1[24949] <= 16'b1111111111110110;
        weights1[24950] <= 16'b0000000000010110;
        weights1[24951] <= 16'b0000000000011001;
        weights1[24952] <= 16'b0000000000101001;
        weights1[24953] <= 16'b0000000000111001;
        weights1[24954] <= 16'b0000000000101011;
        weights1[24955] <= 16'b0000000000100110;
        weights1[24956] <= 16'b1111111111110110;
        weights1[24957] <= 16'b1111111111001001;
        weights1[24958] <= 16'b1111111110011111;
        weights1[24959] <= 16'b1111111110001100;
        weights1[24960] <= 16'b1111111110001010;
        weights1[24961] <= 16'b1111111110001000;
        weights1[24962] <= 16'b1111111111010101;
        weights1[24963] <= 16'b0000000000111110;
        weights1[24964] <= 16'b0000000000111101;
        weights1[24965] <= 16'b0000000000110111;
        weights1[24966] <= 16'b0000000000101101;
        weights1[24967] <= 16'b0000000000011101;
        weights1[24968] <= 16'b1111111111110010;
        weights1[24969] <= 16'b1111111110110011;
        weights1[24970] <= 16'b1111111110101101;
        weights1[24971] <= 16'b1111111110111011;
        weights1[24972] <= 16'b1111111111001110;
        weights1[24973] <= 16'b1111111111100111;
        weights1[24974] <= 16'b1111111111110110;
        weights1[24975] <= 16'b1111111111111011;
        weights1[24976] <= 16'b0000000000001000;
        weights1[24977] <= 16'b0000000000001110;
        weights1[24978] <= 16'b0000000000011110;
        weights1[24979] <= 16'b0000000000100100;
        weights1[24980] <= 16'b0000000000101011;
        weights1[24981] <= 16'b0000000000110110;
        weights1[24982] <= 16'b0000000000110001;
        weights1[24983] <= 16'b0000000000000111;
        weights1[24984] <= 16'b1111111111000100;
        weights1[24985] <= 16'b1111111110001011;
        weights1[24986] <= 16'b1111111101111001;
        weights1[24987] <= 16'b1111111101100000;
        weights1[24988] <= 16'b1111111110011000;
        weights1[24989] <= 16'b1111111111010101;
        weights1[24990] <= 16'b0000000000001110;
        weights1[24991] <= 16'b0000000000111010;
        weights1[24992] <= 16'b0000000001000011;
        weights1[24993] <= 16'b0000000000101100;
        weights1[24994] <= 16'b0000000000100110;
        weights1[24995] <= 16'b0000000000100000;
        weights1[24996] <= 16'b1111111111111100;
        weights1[24997] <= 16'b1111111110111100;
        weights1[24998] <= 16'b1111111110111001;
        weights1[24999] <= 16'b1111111110111100;
        weights1[25000] <= 16'b1111111111001110;
        weights1[25001] <= 16'b1111111111100000;
        weights1[25002] <= 16'b1111111111110100;
        weights1[25003] <= 16'b1111111111110111;
        weights1[25004] <= 16'b0000000000001000;
        weights1[25005] <= 16'b0000000000001101;
        weights1[25006] <= 16'b0000000000100000;
        weights1[25007] <= 16'b0000000000100011;
        weights1[25008] <= 16'b0000000000101110;
        weights1[25009] <= 16'b0000000000100000;
        weights1[25010] <= 16'b1111111111111110;
        weights1[25011] <= 16'b1111111111011000;
        weights1[25012] <= 16'b1111111110100001;
        weights1[25013] <= 16'b1111111110001000;
        weights1[25014] <= 16'b1111111101111000;
        weights1[25015] <= 16'b1111111101111010;
        weights1[25016] <= 16'b1111111110100000;
        weights1[25017] <= 16'b1111111110110110;
        weights1[25018] <= 16'b1111111111111111;
        weights1[25019] <= 16'b0000000000101010;
        weights1[25020] <= 16'b0000000000001111;
        weights1[25021] <= 16'b0000000000101011;
        weights1[25022] <= 16'b0000000000101010;
        weights1[25023] <= 16'b0000000000100000;
        weights1[25024] <= 16'b1111111111111000;
        weights1[25025] <= 16'b1111111111011010;
        weights1[25026] <= 16'b1111111110111011;
        weights1[25027] <= 16'b1111111110111101;
        weights1[25028] <= 16'b1111111111010011;
        weights1[25029] <= 16'b1111111111101001;
        weights1[25030] <= 16'b1111111111110001;
        weights1[25031] <= 16'b1111111111111000;
        weights1[25032] <= 16'b0000000000000111;
        weights1[25033] <= 16'b0000000000000001;
        weights1[25034] <= 16'b0000000000000110;
        weights1[25035] <= 16'b0000000000001001;
        weights1[25036] <= 16'b1111111111111111;
        weights1[25037] <= 16'b1111111111111011;
        weights1[25038] <= 16'b1111111111010101;
        weights1[25039] <= 16'b1111111110100111;
        weights1[25040] <= 16'b1111111110001110;
        weights1[25041] <= 16'b1111111101111110;
        weights1[25042] <= 16'b1111111101111011;
        weights1[25043] <= 16'b1111111110111011;
        weights1[25044] <= 16'b1111111111111100;
        weights1[25045] <= 16'b1111111111111110;
        weights1[25046] <= 16'b0000000000100111;
        weights1[25047] <= 16'b0000000000000001;
        weights1[25048] <= 16'b0000000000010001;
        weights1[25049] <= 16'b0000000000100001;
        weights1[25050] <= 16'b0000000000100101;
        weights1[25051] <= 16'b0000000000100100;
        weights1[25052] <= 16'b0000000000001001;
        weights1[25053] <= 16'b1111111111001111;
        weights1[25054] <= 16'b1111111111000110;
        weights1[25055] <= 16'b1111111111010101;
        weights1[25056] <= 16'b1111111111100011;
        weights1[25057] <= 16'b1111111111101111;
        weights1[25058] <= 16'b1111111111110101;
        weights1[25059] <= 16'b1111111111111110;
        weights1[25060] <= 16'b0000000000000100;
        weights1[25061] <= 16'b0000000000000010;
        weights1[25062] <= 16'b0000000000000001;
        weights1[25063] <= 16'b0000000000000000;
        weights1[25064] <= 16'b1111111111110111;
        weights1[25065] <= 16'b1111111111010111;
        weights1[25066] <= 16'b1111111110111111;
        weights1[25067] <= 16'b1111111110010101;
        weights1[25068] <= 16'b1111111110000111;
        weights1[25069] <= 16'b1111111101111000;
        weights1[25070] <= 16'b1111111110010010;
        weights1[25071] <= 16'b1111111110110010;
        weights1[25072] <= 16'b1111111111101100;
        weights1[25073] <= 16'b1111111111110100;
        weights1[25074] <= 16'b0000000000000000;
        weights1[25075] <= 16'b0000000000011110;
        weights1[25076] <= 16'b0000000001000111;
        weights1[25077] <= 16'b0000000001010100;
        weights1[25078] <= 16'b0000000001000100;
        weights1[25079] <= 16'b0000000000110011;
        weights1[25080] <= 16'b0000000000010100;
        weights1[25081] <= 16'b1111111111101000;
        weights1[25082] <= 16'b1111111111011111;
        weights1[25083] <= 16'b1111111111100100;
        weights1[25084] <= 16'b1111111111110001;
        weights1[25085] <= 16'b1111111111111000;
        weights1[25086] <= 16'b1111111111111010;
        weights1[25087] <= 16'b0000000000000001;
        weights1[25088] <= 16'b0000000000000000;
        weights1[25089] <= 16'b1111111111111111;
        weights1[25090] <= 16'b1111111111111110;
        weights1[25091] <= 16'b1111111111111100;
        weights1[25092] <= 16'b1111111111111101;
        weights1[25093] <= 16'b1111111111111010;
        weights1[25094] <= 16'b1111111111111000;
        weights1[25095] <= 16'b1111111111111001;
        weights1[25096] <= 16'b1111111111110100;
        weights1[25097] <= 16'b1111111111110110;
        weights1[25098] <= 16'b1111111111111011;
        weights1[25099] <= 16'b1111111111111110;
        weights1[25100] <= 16'b0000000000001001;
        weights1[25101] <= 16'b0000000000001001;
        weights1[25102] <= 16'b1111111111111110;
        weights1[25103] <= 16'b1111111111111111;
        weights1[25104] <= 16'b1111111111111001;
        weights1[25105] <= 16'b1111111111110100;
        weights1[25106] <= 16'b1111111111100011;
        weights1[25107] <= 16'b1111111111010001;
        weights1[25108] <= 16'b1111111111011100;
        weights1[25109] <= 16'b1111111111011001;
        weights1[25110] <= 16'b1111111111011011;
        weights1[25111] <= 16'b1111111111011111;
        weights1[25112] <= 16'b1111111111101000;
        weights1[25113] <= 16'b1111111111110000;
        weights1[25114] <= 16'b1111111111110111;
        weights1[25115] <= 16'b1111111111111010;
        weights1[25116] <= 16'b1111111111111111;
        weights1[25117] <= 16'b1111111111111100;
        weights1[25118] <= 16'b1111111111110110;
        weights1[25119] <= 16'b1111111111111010;
        weights1[25120] <= 16'b1111111111111011;
        weights1[25121] <= 16'b1111111111111000;
        weights1[25122] <= 16'b1111111111110001;
        weights1[25123] <= 16'b1111111111110111;
        weights1[25124] <= 16'b1111111111111011;
        weights1[25125] <= 16'b1111111111110000;
        weights1[25126] <= 16'b1111111111111011;
        weights1[25127] <= 16'b0000000000000100;
        weights1[25128] <= 16'b0000000000001001;
        weights1[25129] <= 16'b0000000000000100;
        weights1[25130] <= 16'b0000000000000010;
        weights1[25131] <= 16'b1111111111111000;
        weights1[25132] <= 16'b0000000000000000;
        weights1[25133] <= 16'b0000000000001010;
        weights1[25134] <= 16'b1111111111111011;
        weights1[25135] <= 16'b1111111111101100;
        weights1[25136] <= 16'b1111111111010011;
        weights1[25137] <= 16'b1111111111010101;
        weights1[25138] <= 16'b1111111111001010;
        weights1[25139] <= 16'b1111111111010100;
        weights1[25140] <= 16'b1111111111011101;
        weights1[25141] <= 16'b1111111111100101;
        weights1[25142] <= 16'b1111111111110100;
        weights1[25143] <= 16'b1111111111110111;
        weights1[25144] <= 16'b1111111111111111;
        weights1[25145] <= 16'b1111111111111001;
        weights1[25146] <= 16'b1111111111111001;
        weights1[25147] <= 16'b1111111111110111;
        weights1[25148] <= 16'b1111111111110101;
        weights1[25149] <= 16'b1111111111110011;
        weights1[25150] <= 16'b1111111111101011;
        weights1[25151] <= 16'b1111111111111010;
        weights1[25152] <= 16'b0000000000000100;
        weights1[25153] <= 16'b0000000000000110;
        weights1[25154] <= 16'b1111111111111100;
        weights1[25155] <= 16'b1111111111101101;
        weights1[25156] <= 16'b1111111111111101;
        weights1[25157] <= 16'b0000000000000011;
        weights1[25158] <= 16'b0000000000010110;
        weights1[25159] <= 16'b0000000000001001;
        weights1[25160] <= 16'b0000000000000110;
        weights1[25161] <= 16'b0000000000001100;
        weights1[25162] <= 16'b0000000000001111;
        weights1[25163] <= 16'b0000000000001001;
        weights1[25164] <= 16'b1111111111110000;
        weights1[25165] <= 16'b1111111111100111;
        weights1[25166] <= 16'b1111111111001001;
        weights1[25167] <= 16'b1111111111001110;
        weights1[25168] <= 16'b1111111111010110;
        weights1[25169] <= 16'b1111111111011001;
        weights1[25170] <= 16'b1111111111101100;
        weights1[25171] <= 16'b1111111111101111;
        weights1[25172] <= 16'b1111111111111101;
        weights1[25173] <= 16'b1111111111111100;
        weights1[25174] <= 16'b1111111111111011;
        weights1[25175] <= 16'b1111111111110001;
        weights1[25176] <= 16'b1111111111110010;
        weights1[25177] <= 16'b1111111111110100;
        weights1[25178] <= 16'b1111111111110100;
        weights1[25179] <= 16'b1111111111111001;
        weights1[25180] <= 16'b1111111111111110;
        weights1[25181] <= 16'b1111111111111001;
        weights1[25182] <= 16'b1111111111101111;
        weights1[25183] <= 16'b1111111111110010;
        weights1[25184] <= 16'b0000000000001000;
        weights1[25185] <= 16'b0000000000001011;
        weights1[25186] <= 16'b0000000000011000;
        weights1[25187] <= 16'b1111111111111101;
        weights1[25188] <= 16'b0000000000011011;
        weights1[25189] <= 16'b0000000000100101;
        weights1[25190] <= 16'b0000000000001111;
        weights1[25191] <= 16'b0000000000010010;
        weights1[25192] <= 16'b0000000000010011;
        weights1[25193] <= 16'b1111111111110101;
        weights1[25194] <= 16'b1111111111011010;
        weights1[25195] <= 16'b1111111111001010;
        weights1[25196] <= 16'b1111111111001000;
        weights1[25197] <= 16'b1111111111001111;
        weights1[25198] <= 16'b1111111111011101;
        weights1[25199] <= 16'b1111111111100110;
        weights1[25200] <= 16'b1111111111111111;
        weights1[25201] <= 16'b1111111111111001;
        weights1[25202] <= 16'b1111111111110011;
        weights1[25203] <= 16'b1111111111101110;
        weights1[25204] <= 16'b1111111111101101;
        weights1[25205] <= 16'b1111111111110000;
        weights1[25206] <= 16'b1111111111111001;
        weights1[25207] <= 16'b1111111111101111;
        weights1[25208] <= 16'b1111111111111011;
        weights1[25209] <= 16'b1111111111111001;
        weights1[25210] <= 16'b1111111111110111;
        weights1[25211] <= 16'b0000000000000001;
        weights1[25212] <= 16'b0000000000001010;
        weights1[25213] <= 16'b1111111111110101;
        weights1[25214] <= 16'b0000000000010001;
        weights1[25215] <= 16'b0000000000011100;
        weights1[25216] <= 16'b0000000000100000;
        weights1[25217] <= 16'b0000000000110110;
        weights1[25218] <= 16'b0000000000101100;
        weights1[25219] <= 16'b0000000000010101;
        weights1[25220] <= 16'b0000000000101001;
        weights1[25221] <= 16'b0000000000001011;
        weights1[25222] <= 16'b1111111111110101;
        weights1[25223] <= 16'b1111111111011100;
        weights1[25224] <= 16'b1111111111001110;
        weights1[25225] <= 16'b1111111111000110;
        weights1[25226] <= 16'b1111111111010100;
        weights1[25227] <= 16'b1111111111101010;
        weights1[25228] <= 16'b0000000000000000;
        weights1[25229] <= 16'b1111111111110110;
        weights1[25230] <= 16'b1111111111101100;
        weights1[25231] <= 16'b1111111111101101;
        weights1[25232] <= 16'b1111111111100100;
        weights1[25233] <= 16'b1111111111100010;
        weights1[25234] <= 16'b1111111111101011;
        weights1[25235] <= 16'b1111111111110101;
        weights1[25236] <= 16'b1111111111011110;
        weights1[25237] <= 16'b1111111111101011;
        weights1[25238] <= 16'b1111111111110011;
        weights1[25239] <= 16'b1111111111101100;
        weights1[25240] <= 16'b0000000000000101;
        weights1[25241] <= 16'b0000000000000010;
        weights1[25242] <= 16'b0000000000000000;
        weights1[25243] <= 16'b0000000000011011;
        weights1[25244] <= 16'b0000000000010111;
        weights1[25245] <= 16'b0000000000101000;
        weights1[25246] <= 16'b0000000000011011;
        weights1[25247] <= 16'b0000000000101011;
        weights1[25248] <= 16'b0000000000110111;
        weights1[25249] <= 16'b0000000000010110;
        weights1[25250] <= 16'b0000000000000110;
        weights1[25251] <= 16'b1111111111101000;
        weights1[25252] <= 16'b1111111111011011;
        weights1[25253] <= 16'b1111111111010110;
        weights1[25254] <= 16'b1111111111011001;
        weights1[25255] <= 16'b1111111111011111;
        weights1[25256] <= 16'b1111111111111100;
        weights1[25257] <= 16'b1111111111110100;
        weights1[25258] <= 16'b1111111111101110;
        weights1[25259] <= 16'b1111111111110111;
        weights1[25260] <= 16'b1111111111101101;
        weights1[25261] <= 16'b1111111111101100;
        weights1[25262] <= 16'b1111111111111010;
        weights1[25263] <= 16'b1111111111101111;
        weights1[25264] <= 16'b1111111111101011;
        weights1[25265] <= 16'b1111111111101101;
        weights1[25266] <= 16'b1111111111100010;
        weights1[25267] <= 16'b1111111111110001;
        weights1[25268] <= 16'b1111111111110010;
        weights1[25269] <= 16'b1111111111111111;
        weights1[25270] <= 16'b1111111111101110;
        weights1[25271] <= 16'b0000000000000000;
        weights1[25272] <= 16'b0000000000001000;
        weights1[25273] <= 16'b0000000000100100;
        weights1[25274] <= 16'b0000000000101001;
        weights1[25275] <= 16'b0000000000101011;
        weights1[25276] <= 16'b0000000000110101;
        weights1[25277] <= 16'b0000000000101010;
        weights1[25278] <= 16'b0000000000011000;
        weights1[25279] <= 16'b0000000000000101;
        weights1[25280] <= 16'b1111111111011111;
        weights1[25281] <= 16'b1111111111010110;
        weights1[25282] <= 16'b1111111111010101;
        weights1[25283] <= 16'b1111111111011001;
        weights1[25284] <= 16'b1111111111111100;
        weights1[25285] <= 16'b1111111111110111;
        weights1[25286] <= 16'b1111111111110011;
        weights1[25287] <= 16'b1111111111110111;
        weights1[25288] <= 16'b1111111111110110;
        weights1[25289] <= 16'b1111111111101000;
        weights1[25290] <= 16'b1111111111110010;
        weights1[25291] <= 16'b1111111111111001;
        weights1[25292] <= 16'b1111111111110000;
        weights1[25293] <= 16'b1111111111110110;
        weights1[25294] <= 16'b1111111111110110;
        weights1[25295] <= 16'b1111111111111010;
        weights1[25296] <= 16'b1111111111110011;
        weights1[25297] <= 16'b1111111111101111;
        weights1[25298] <= 16'b1111111111101111;
        weights1[25299] <= 16'b1111111111110110;
        weights1[25300] <= 16'b0000000000001010;
        weights1[25301] <= 16'b0000000000101011;
        weights1[25302] <= 16'b0000000001000000;
        weights1[25303] <= 16'b0000000000110010;
        weights1[25304] <= 16'b0000000000110001;
        weights1[25305] <= 16'b0000000000101000;
        weights1[25306] <= 16'b0000000000011111;
        weights1[25307] <= 16'b0000000000010100;
        weights1[25308] <= 16'b1111111111110100;
        weights1[25309] <= 16'b1111111111100111;
        weights1[25310] <= 16'b1111111111011001;
        weights1[25311] <= 16'b1111111111100000;
        weights1[25312] <= 16'b1111111111111010;
        weights1[25313] <= 16'b1111111111111001;
        weights1[25314] <= 16'b1111111111110001;
        weights1[25315] <= 16'b1111111111110000;
        weights1[25316] <= 16'b1111111111111011;
        weights1[25317] <= 16'b1111111111101111;
        weights1[25318] <= 16'b1111111111011101;
        weights1[25319] <= 16'b0000000000000111;
        weights1[25320] <= 16'b1111111111111110;
        weights1[25321] <= 16'b1111111111100010;
        weights1[25322] <= 16'b1111111111110101;
        weights1[25323] <= 16'b1111111111101110;
        weights1[25324] <= 16'b1111111111110000;
        weights1[25325] <= 16'b1111111111100101;
        weights1[25326] <= 16'b1111111111011111;
        weights1[25327] <= 16'b1111111111110001;
        weights1[25328] <= 16'b1111111111110011;
        weights1[25329] <= 16'b0000000000011001;
        weights1[25330] <= 16'b0000000001000001;
        weights1[25331] <= 16'b0000000000110110;
        weights1[25332] <= 16'b0000000000100110;
        weights1[25333] <= 16'b0000000000111011;
        weights1[25334] <= 16'b0000000000100010;
        weights1[25335] <= 16'b0000000000011001;
        weights1[25336] <= 16'b1111111111110101;
        weights1[25337] <= 16'b1111111111011111;
        weights1[25338] <= 16'b1111111111100000;
        weights1[25339] <= 16'b1111111111011101;
        weights1[25340] <= 16'b0000000000000010;
        weights1[25341] <= 16'b1111111111111001;
        weights1[25342] <= 16'b1111111111110011;
        weights1[25343] <= 16'b1111111111110110;
        weights1[25344] <= 16'b0000000000000101;
        weights1[25345] <= 16'b1111111111111011;
        weights1[25346] <= 16'b0000000000001100;
        weights1[25347] <= 16'b1111111111111101;
        weights1[25348] <= 16'b1111111111111011;
        weights1[25349] <= 16'b1111111111111010;
        weights1[25350] <= 16'b0000000000000001;
        weights1[25351] <= 16'b0000000000000101;
        weights1[25352] <= 16'b1111111111110100;
        weights1[25353] <= 16'b1111111111101001;
        weights1[25354] <= 16'b1111111111100010;
        weights1[25355] <= 16'b1111111111010010;
        weights1[25356] <= 16'b1111111111010011;
        weights1[25357] <= 16'b1111111111111100;
        weights1[25358] <= 16'b0000000000111001;
        weights1[25359] <= 16'b0000000001000010;
        weights1[25360] <= 16'b0000000000101011;
        weights1[25361] <= 16'b0000000000101000;
        weights1[25362] <= 16'b0000000000011100;
        weights1[25363] <= 16'b0000000000010001;
        weights1[25364] <= 16'b0000000000000101;
        weights1[25365] <= 16'b1111111111101010;
        weights1[25366] <= 16'b1111111111100110;
        weights1[25367] <= 16'b1111111111100011;
        weights1[25368] <= 16'b0000000000000010;
        weights1[25369] <= 16'b0000000000000011;
        weights1[25370] <= 16'b1111111111111101;
        weights1[25371] <= 16'b0000000000001011;
        weights1[25372] <= 16'b0000000000000010;
        weights1[25373] <= 16'b0000000000001001;
        weights1[25374] <= 16'b1111111111111010;
        weights1[25375] <= 16'b1111111111111010;
        weights1[25376] <= 16'b1111111111110101;
        weights1[25377] <= 16'b0000000000000000;
        weights1[25378] <= 16'b1111111111100100;
        weights1[25379] <= 16'b1111111111101010;
        weights1[25380] <= 16'b1111111111101010;
        weights1[25381] <= 16'b1111111111100000;
        weights1[25382] <= 16'b1111111111010101;
        weights1[25383] <= 16'b1111111111011110;
        weights1[25384] <= 16'b1111111111000001;
        weights1[25385] <= 16'b1111111111111100;
        weights1[25386] <= 16'b0000000000101111;
        weights1[25387] <= 16'b0000000000111111;
        weights1[25388] <= 16'b0000000000111111;
        weights1[25389] <= 16'b0000000000101000;
        weights1[25390] <= 16'b0000000000101110;
        weights1[25391] <= 16'b0000000000100110;
        weights1[25392] <= 16'b1111111111111100;
        weights1[25393] <= 16'b1111111111110000;
        weights1[25394] <= 16'b1111111111100000;
        weights1[25395] <= 16'b1111111111100011;
        weights1[25396] <= 16'b0000000000000011;
        weights1[25397] <= 16'b0000000000001010;
        weights1[25398] <= 16'b0000000000001111;
        weights1[25399] <= 16'b0000000000001011;
        weights1[25400] <= 16'b1111111111111011;
        weights1[25401] <= 16'b1111111111111011;
        weights1[25402] <= 16'b1111111111110100;
        weights1[25403] <= 16'b1111111111110111;
        weights1[25404] <= 16'b1111111111101110;
        weights1[25405] <= 16'b1111111111111011;
        weights1[25406] <= 16'b1111111111101101;
        weights1[25407] <= 16'b1111111111111000;
        weights1[25408] <= 16'b1111111111101001;
        weights1[25409] <= 16'b1111111111110010;
        weights1[25410] <= 16'b1111111111101100;
        weights1[25411] <= 16'b1111111111011001;
        weights1[25412] <= 16'b1111111111001110;
        weights1[25413] <= 16'b1111111111101101;
        weights1[25414] <= 16'b0000000000010011;
        weights1[25415] <= 16'b0000000000101000;
        weights1[25416] <= 16'b0000000000110011;
        weights1[25417] <= 16'b0000000000100110;
        weights1[25418] <= 16'b0000000000101110;
        weights1[25419] <= 16'b0000000000100110;
        weights1[25420] <= 16'b0000000000000100;
        weights1[25421] <= 16'b1111111111101110;
        weights1[25422] <= 16'b1111111111100010;
        weights1[25423] <= 16'b1111111111111000;
        weights1[25424] <= 16'b0000000000000111;
        weights1[25425] <= 16'b0000000000001100;
        weights1[25426] <= 16'b0000000000001000;
        weights1[25427] <= 16'b1111111111111010;
        weights1[25428] <= 16'b1111111111110100;
        weights1[25429] <= 16'b0000000000000100;
        weights1[25430] <= 16'b1111111111110010;
        weights1[25431] <= 16'b1111111111100001;
        weights1[25432] <= 16'b0000000000000100;
        weights1[25433] <= 16'b1111111111101101;
        weights1[25434] <= 16'b1111111111101000;
        weights1[25435] <= 16'b1111111111111000;
        weights1[25436] <= 16'b1111111111110010;
        weights1[25437] <= 16'b1111111111110001;
        weights1[25438] <= 16'b1111111111101011;
        weights1[25439] <= 16'b1111111111010011;
        weights1[25440] <= 16'b1111111110111001;
        weights1[25441] <= 16'b1111111111001100;
        weights1[25442] <= 16'b0000000000000100;
        weights1[25443] <= 16'b0000000000011100;
        weights1[25444] <= 16'b0000000000100000;
        weights1[25445] <= 16'b0000000000010110;
        weights1[25446] <= 16'b0000000000011110;
        weights1[25447] <= 16'b0000000000001101;
        weights1[25448] <= 16'b0000000000000101;
        weights1[25449] <= 16'b1111111111111000;
        weights1[25450] <= 16'b1111111111100100;
        weights1[25451] <= 16'b1111111111101111;
        weights1[25452] <= 16'b0000000000000111;
        weights1[25453] <= 16'b0000000000010000;
        weights1[25454] <= 16'b0000000000000000;
        weights1[25455] <= 16'b1111111111101101;
        weights1[25456] <= 16'b1111111111111010;
        weights1[25457] <= 16'b1111111111111011;
        weights1[25458] <= 16'b1111111111110100;
        weights1[25459] <= 16'b1111111111101111;
        weights1[25460] <= 16'b0000000000000000;
        weights1[25461] <= 16'b1111111111101101;
        weights1[25462] <= 16'b1111111111110011;
        weights1[25463] <= 16'b1111111111111000;
        weights1[25464] <= 16'b1111111111111010;
        weights1[25465] <= 16'b1111111111110110;
        weights1[25466] <= 16'b1111111111011110;
        weights1[25467] <= 16'b1111111110111001;
        weights1[25468] <= 16'b1111111110111101;
        weights1[25469] <= 16'b1111111111011000;
        weights1[25470] <= 16'b0000000000000101;
        weights1[25471] <= 16'b0000000000011010;
        weights1[25472] <= 16'b0000000000000101;
        weights1[25473] <= 16'b0000000000010110;
        weights1[25474] <= 16'b0000000000001001;
        weights1[25475] <= 16'b0000000000011011;
        weights1[25476] <= 16'b1111111111111110;
        weights1[25477] <= 16'b1111111111110111;
        weights1[25478] <= 16'b1111111111100110;
        weights1[25479] <= 16'b1111111111101110;
        weights1[25480] <= 16'b0000000000001011;
        weights1[25481] <= 16'b0000000000001001;
        weights1[25482] <= 16'b1111111111111010;
        weights1[25483] <= 16'b1111111111111011;
        weights1[25484] <= 16'b1111111111100101;
        weights1[25485] <= 16'b0000000000000101;
        weights1[25486] <= 16'b1111111111101010;
        weights1[25487] <= 16'b1111111111111011;
        weights1[25488] <= 16'b1111111111110010;
        weights1[25489] <= 16'b1111111111111110;
        weights1[25490] <= 16'b0000000000000010;
        weights1[25491] <= 16'b0000000000000010;
        weights1[25492] <= 16'b1111111111110110;
        weights1[25493] <= 16'b1111111111111000;
        weights1[25494] <= 16'b1111111111011010;
        weights1[25495] <= 16'b1111111111010010;
        weights1[25496] <= 16'b1111111110111100;
        weights1[25497] <= 16'b1111111111101000;
        weights1[25498] <= 16'b0000000000001101;
        weights1[25499] <= 16'b0000000000000001;
        weights1[25500] <= 16'b0000000000010100;
        weights1[25501] <= 16'b0000000000001101;
        weights1[25502] <= 16'b0000000000010011;
        weights1[25503] <= 16'b0000000000011011;
        weights1[25504] <= 16'b1111111111111001;
        weights1[25505] <= 16'b1111111111110001;
        weights1[25506] <= 16'b1111111111101111;
        weights1[25507] <= 16'b1111111111111001;
        weights1[25508] <= 16'b0000000000001101;
        weights1[25509] <= 16'b0000000000000100;
        weights1[25510] <= 16'b0000000000000110;
        weights1[25511] <= 16'b0000000000000011;
        weights1[25512] <= 16'b1111111111111010;
        weights1[25513] <= 16'b0000000000010001;
        weights1[25514] <= 16'b1111111111110010;
        weights1[25515] <= 16'b0000000000001100;
        weights1[25516] <= 16'b0000000000000110;
        weights1[25517] <= 16'b0000000000001111;
        weights1[25518] <= 16'b1111111111110101;
        weights1[25519] <= 16'b1111111111101111;
        weights1[25520] <= 16'b1111111111101100;
        weights1[25521] <= 16'b1111111111110001;
        weights1[25522] <= 16'b1111111111011011;
        weights1[25523] <= 16'b1111111111010010;
        weights1[25524] <= 16'b1111111111010110;
        weights1[25525] <= 16'b1111111111110100;
        weights1[25526] <= 16'b0000000000010011;
        weights1[25527] <= 16'b0000000000010111;
        weights1[25528] <= 16'b0000000000001000;
        weights1[25529] <= 16'b0000000000001000;
        weights1[25530] <= 16'b0000000000010010;
        weights1[25531] <= 16'b0000000000000001;
        weights1[25532] <= 16'b1111111111110001;
        weights1[25533] <= 16'b1111111111110010;
        weights1[25534] <= 16'b1111111111101110;
        weights1[25535] <= 16'b0000000000000110;
        weights1[25536] <= 16'b0000000000001001;
        weights1[25537] <= 16'b0000000000001010;
        weights1[25538] <= 16'b0000000000010000;
        weights1[25539] <= 16'b1111111111111110;
        weights1[25540] <= 16'b0000000000001010;
        weights1[25541] <= 16'b0000000000000101;
        weights1[25542] <= 16'b1111111111111101;
        weights1[25543] <= 16'b0000000000000000;
        weights1[25544] <= 16'b0000000000001011;
        weights1[25545] <= 16'b1111111111111001;
        weights1[25546] <= 16'b1111111111101101;
        weights1[25547] <= 16'b1111111111110100;
        weights1[25548] <= 16'b1111111111100011;
        weights1[25549] <= 16'b1111111111011110;
        weights1[25550] <= 16'b1111111111010100;
        weights1[25551] <= 16'b1111111111011111;
        weights1[25552] <= 16'b1111111111110001;
        weights1[25553] <= 16'b0000000000000111;
        weights1[25554] <= 16'b0000000000001100;
        weights1[25555] <= 16'b0000000000001010;
        weights1[25556] <= 16'b0000000000010111;
        weights1[25557] <= 16'b0000000000010110;
        weights1[25558] <= 16'b0000000000000101;
        weights1[25559] <= 16'b1111111111111000;
        weights1[25560] <= 16'b0000000000000000;
        weights1[25561] <= 16'b1111111111111100;
        weights1[25562] <= 16'b1111111111110110;
        weights1[25563] <= 16'b0000000000000010;
        weights1[25564] <= 16'b0000000000001001;
        weights1[25565] <= 16'b0000000000001001;
        weights1[25566] <= 16'b0000000000011000;
        weights1[25567] <= 16'b0000000000000010;
        weights1[25568] <= 16'b0000000000011010;
        weights1[25569] <= 16'b0000000000000001;
        weights1[25570] <= 16'b1111111111111111;
        weights1[25571] <= 16'b1111111111111100;
        weights1[25572] <= 16'b1111111111111111;
        weights1[25573] <= 16'b1111111111111111;
        weights1[25574] <= 16'b1111111111111011;
        weights1[25575] <= 16'b1111111111110011;
        weights1[25576] <= 16'b1111111111100000;
        weights1[25577] <= 16'b1111111111110100;
        weights1[25578] <= 16'b1111111111101001;
        weights1[25579] <= 16'b1111111111110010;
        weights1[25580] <= 16'b1111111111110110;
        weights1[25581] <= 16'b0000000000000000;
        weights1[25582] <= 16'b0000000000001111;
        weights1[25583] <= 16'b0000000000010110;
        weights1[25584] <= 16'b0000000000001100;
        weights1[25585] <= 16'b1111111111110010;
        weights1[25586] <= 16'b1111111111110111;
        weights1[25587] <= 16'b1111111111100100;
        weights1[25588] <= 16'b1111111111101111;
        weights1[25589] <= 16'b1111111111110111;
        weights1[25590] <= 16'b1111111111111100;
        weights1[25591] <= 16'b0000000000000010;
        weights1[25592] <= 16'b0000000000000100;
        weights1[25593] <= 16'b0000000000000000;
        weights1[25594] <= 16'b0000000000001010;
        weights1[25595] <= 16'b0000000000000110;
        weights1[25596] <= 16'b0000000000001011;
        weights1[25597] <= 16'b0000000000010000;
        weights1[25598] <= 16'b0000000000010000;
        weights1[25599] <= 16'b1111111111111110;
        weights1[25600] <= 16'b0000000000000101;
        weights1[25601] <= 16'b0000000000000001;
        weights1[25602] <= 16'b0000000000010011;
        weights1[25603] <= 16'b1111111111101001;
        weights1[25604] <= 16'b1111111111100011;
        weights1[25605] <= 16'b1111111111101100;
        weights1[25606] <= 16'b1111111111110110;
        weights1[25607] <= 16'b1111111111110010;
        weights1[25608] <= 16'b1111111111110101;
        weights1[25609] <= 16'b1111111111111111;
        weights1[25610] <= 16'b1111111111111000;
        weights1[25611] <= 16'b0000000000001011;
        weights1[25612] <= 16'b1111111111101110;
        weights1[25613] <= 16'b1111111111101101;
        weights1[25614] <= 16'b1111111111101010;
        weights1[25615] <= 16'b1111111111100000;
        weights1[25616] <= 16'b1111111111101110;
        weights1[25617] <= 16'b1111111111110001;
        weights1[25618] <= 16'b1111111111111000;
        weights1[25619] <= 16'b1111111111111011;
        weights1[25620] <= 16'b0000000000000000;
        weights1[25621] <= 16'b1111111111111111;
        weights1[25622] <= 16'b1111111111111010;
        weights1[25623] <= 16'b0000000000000001;
        weights1[25624] <= 16'b1111111111110101;
        weights1[25625] <= 16'b0000000000000001;
        weights1[25626] <= 16'b0000000000000010;
        weights1[25627] <= 16'b1111111111111001;
        weights1[25628] <= 16'b0000000000001100;
        weights1[25629] <= 16'b0000000000010010;
        weights1[25630] <= 16'b0000000000000110;
        weights1[25631] <= 16'b0000000000000000;
        weights1[25632] <= 16'b1111111111111000;
        weights1[25633] <= 16'b1111111111111101;
        weights1[25634] <= 16'b0000000000001001;
        weights1[25635] <= 16'b0000000000000000;
        weights1[25636] <= 16'b1111111111111111;
        weights1[25637] <= 16'b0000000000000011;
        weights1[25638] <= 16'b1111111111111100;
        weights1[25639] <= 16'b0000000000000100;
        weights1[25640] <= 16'b1111111111110100;
        weights1[25641] <= 16'b1111111111110100;
        weights1[25642] <= 16'b1111111111111011;
        weights1[25643] <= 16'b1111111111111010;
        weights1[25644] <= 16'b1111111111110100;
        weights1[25645] <= 16'b1111111111111000;
        weights1[25646] <= 16'b1111111111111010;
        weights1[25647] <= 16'b0000000000000100;
        weights1[25648] <= 16'b1111111111111100;
        weights1[25649] <= 16'b1111111111111001;
        weights1[25650] <= 16'b1111111111110110;
        weights1[25651] <= 16'b0000000000000101;
        weights1[25652] <= 16'b0000000000000111;
        weights1[25653] <= 16'b0000000000001101;
        weights1[25654] <= 16'b0000000000000011;
        weights1[25655] <= 16'b1111111111110101;
        weights1[25656] <= 16'b1111111111111001;
        weights1[25657] <= 16'b1111111111111111;
        weights1[25658] <= 16'b0000000000011010;
        weights1[25659] <= 16'b0000000000000011;
        weights1[25660] <= 16'b0000000000001011;
        weights1[25661] <= 16'b0000000000001000;
        weights1[25662] <= 16'b0000000000001000;
        weights1[25663] <= 16'b0000000000000001;
        weights1[25664] <= 16'b1111111111110011;
        weights1[25665] <= 16'b0000000000001001;
        weights1[25666] <= 16'b0000000000000110;
        weights1[25667] <= 16'b1111111111111111;
        weights1[25668] <= 16'b1111111111110110;
        weights1[25669] <= 16'b0000000000000101;
        weights1[25670] <= 16'b1111111111111010;
        weights1[25671] <= 16'b0000000000001010;
        weights1[25672] <= 16'b1111111111110101;
        weights1[25673] <= 16'b0000000000000000;
        weights1[25674] <= 16'b0000000000000000;
        weights1[25675] <= 16'b0000000000001101;
        weights1[25676] <= 16'b1111111111111011;
        weights1[25677] <= 16'b0000000000000001;
        weights1[25678] <= 16'b1111111111110010;
        weights1[25679] <= 16'b1111111111111001;
        weights1[25680] <= 16'b0000000000001000;
        weights1[25681] <= 16'b0000000000010110;
        weights1[25682] <= 16'b0000000000000001;
        weights1[25683] <= 16'b1111111111111111;
        weights1[25684] <= 16'b1111111111110100;
        weights1[25685] <= 16'b1111111111111010;
        weights1[25686] <= 16'b1111111111111110;
        weights1[25687] <= 16'b0000000000010110;
        weights1[25688] <= 16'b0000000000001011;
        weights1[25689] <= 16'b0000000000000111;
        weights1[25690] <= 16'b0000000000000001;
        weights1[25691] <= 16'b1111111111111000;
        weights1[25692] <= 16'b0000000000000001;
        weights1[25693] <= 16'b1111111111111101;
        weights1[25694] <= 16'b1111111111110001;
        weights1[25695] <= 16'b1111111111111111;
        weights1[25696] <= 16'b1111111111110010;
        weights1[25697] <= 16'b1111111111111111;
        weights1[25698] <= 16'b1111111111111100;
        weights1[25699] <= 16'b0000000000010000;
        weights1[25700] <= 16'b0000000000001110;
        weights1[25701] <= 16'b0000000000000001;
        weights1[25702] <= 16'b0000000000000000;
        weights1[25703] <= 16'b0000000000001111;
        weights1[25704] <= 16'b1111111111111110;
        weights1[25705] <= 16'b1111111111111101;
        weights1[25706] <= 16'b1111111111111111;
        weights1[25707] <= 16'b1111111111111110;
        weights1[25708] <= 16'b1111111111111011;
        weights1[25709] <= 16'b1111111111111000;
        weights1[25710] <= 16'b1111111111110011;
        weights1[25711] <= 16'b0000000000001001;
        weights1[25712] <= 16'b1111111111111010;
        weights1[25713] <= 16'b0000000000001011;
        weights1[25714] <= 16'b0000000000010111;
        weights1[25715] <= 16'b0000000000010011;
        weights1[25716] <= 16'b0000000000010011;
        weights1[25717] <= 16'b0000000000000001;
        weights1[25718] <= 16'b1111111111111111;
        weights1[25719] <= 16'b1111111111110010;
        weights1[25720] <= 16'b0000000000001101;
        weights1[25721] <= 16'b1111111111111101;
        weights1[25722] <= 16'b1111111111111101;
        weights1[25723] <= 16'b1111111111111110;
        weights1[25724] <= 16'b1111111111111110;
        weights1[25725] <= 16'b0000000000000010;
        weights1[25726] <= 16'b1111111111111001;
        weights1[25727] <= 16'b0000000000011011;
        weights1[25728] <= 16'b0000000000000000;
        weights1[25729] <= 16'b1111111111111001;
        weights1[25730] <= 16'b0000000000001001;
        weights1[25731] <= 16'b0000000000001001;
        weights1[25732] <= 16'b1111111111111110;
        weights1[25733] <= 16'b0000000000000000;
        weights1[25734] <= 16'b1111111111111111;
        weights1[25735] <= 16'b1111111111111010;
        weights1[25736] <= 16'b1111111111111101;
        weights1[25737] <= 16'b1111111111110101;
        weights1[25738] <= 16'b0000000000001111;
        weights1[25739] <= 16'b0000000000001101;
        weights1[25740] <= 16'b0000000000000010;
        weights1[25741] <= 16'b1111111111111011;
        weights1[25742] <= 16'b0000000000011100;
        weights1[25743] <= 16'b0000000000010111;
        weights1[25744] <= 16'b0000000000001100;
        weights1[25745] <= 16'b0000000000000101;
        weights1[25746] <= 16'b0000000000001010;
        weights1[25747] <= 16'b1111111111111100;
        weights1[25748] <= 16'b0000000000010001;
        weights1[25749] <= 16'b0000000000000101;
        weights1[25750] <= 16'b1111111111110101;
        weights1[25751] <= 16'b1111111111111111;
        weights1[25752] <= 16'b1111111111111101;
        weights1[25753] <= 16'b0000000000001110;
        weights1[25754] <= 16'b0000000000000101;
        weights1[25755] <= 16'b0000000000001011;
        weights1[25756] <= 16'b0000000000000001;
        weights1[25757] <= 16'b1111111111111110;
        weights1[25758] <= 16'b1111111111111111;
        weights1[25759] <= 16'b0000000000000101;
        weights1[25760] <= 16'b0000000000000000;
        weights1[25761] <= 16'b1111111111111101;
        weights1[25762] <= 16'b1111111111111011;
        weights1[25763] <= 16'b1111111111111001;
        weights1[25764] <= 16'b0000000000000110;
        weights1[25765] <= 16'b0000000000011000;
        weights1[25766] <= 16'b0000000000010011;
        weights1[25767] <= 16'b0000000000000000;
        weights1[25768] <= 16'b1111111111111001;
        weights1[25769] <= 16'b0000000000010000;
        weights1[25770] <= 16'b0000000000011110;
        weights1[25771] <= 16'b0000000000001010;
        weights1[25772] <= 16'b0000000000000111;
        weights1[25773] <= 16'b1111111111110111;
        weights1[25774] <= 16'b1111111111101101;
        weights1[25775] <= 16'b1111111111101011;
        weights1[25776] <= 16'b0000000000001000;
        weights1[25777] <= 16'b1111111111111011;
        weights1[25778] <= 16'b1111111111111000;
        weights1[25779] <= 16'b0000000000000000;
        weights1[25780] <= 16'b0000000000000010;
        weights1[25781] <= 16'b0000000000001000;
        weights1[25782] <= 16'b1111111111111010;
        weights1[25783] <= 16'b1111111111111111;
        weights1[25784] <= 16'b0000000000000000;
        weights1[25785] <= 16'b0000000000000101;
        weights1[25786] <= 16'b1111111111111011;
        weights1[25787] <= 16'b1111111111111110;
        weights1[25788] <= 16'b1111111111111111;
        weights1[25789] <= 16'b1111111111111110;
        weights1[25790] <= 16'b1111111111111001;
        weights1[25791] <= 16'b1111111111111000;
        weights1[25792] <= 16'b1111111111111111;
        weights1[25793] <= 16'b0000000000000011;
        weights1[25794] <= 16'b0000000000000100;
        weights1[25795] <= 16'b0000000000001010;
        weights1[25796] <= 16'b0000000000010101;
        weights1[25797] <= 16'b0000000000011101;
        weights1[25798] <= 16'b0000000000011101;
        weights1[25799] <= 16'b0000000000000000;
        weights1[25800] <= 16'b1111111111111011;
        weights1[25801] <= 16'b1111111111111101;
        weights1[25802] <= 16'b1111111111110101;
        weights1[25803] <= 16'b1111111111110010;
        weights1[25804] <= 16'b1111111111110011;
        weights1[25805] <= 16'b1111111111111010;
        weights1[25806] <= 16'b1111111111111010;
        weights1[25807] <= 16'b1111111111110101;
        weights1[25808] <= 16'b1111111111110110;
        weights1[25809] <= 16'b0000000000001001;
        weights1[25810] <= 16'b1111111111111000;
        weights1[25811] <= 16'b1111111111111100;
        weights1[25812] <= 16'b1111111111111100;
        weights1[25813] <= 16'b1111111111111011;
        weights1[25814] <= 16'b1111111111111000;
        weights1[25815] <= 16'b1111111111111110;
        weights1[25816] <= 16'b1111111111111110;
        weights1[25817] <= 16'b0000000000000001;
        weights1[25818] <= 16'b1111111111111000;
        weights1[25819] <= 16'b1111111111111011;
        weights1[25820] <= 16'b1111111111111111;
        weights1[25821] <= 16'b1111111111110010;
        weights1[25822] <= 16'b1111111111110010;
        weights1[25823] <= 16'b1111111111111110;
        weights1[25824] <= 16'b0000000000001101;
        weights1[25825] <= 16'b0000000000001110;
        weights1[25826] <= 16'b0000000000000101;
        weights1[25827] <= 16'b1111111111110001;
        weights1[25828] <= 16'b1111111111101000;
        weights1[25829] <= 16'b1111111111111000;
        weights1[25830] <= 16'b1111111111111001;
        weights1[25831] <= 16'b0000000000000000;
        weights1[25832] <= 16'b1111111111111000;
        weights1[25833] <= 16'b0000000000000000;
        weights1[25834] <= 16'b1111111111110001;
        weights1[25835] <= 16'b1111111111110101;
        weights1[25836] <= 16'b0000000000001010;
        weights1[25837] <= 16'b0000000000000010;
        weights1[25838] <= 16'b1111111111111111;
        weights1[25839] <= 16'b1111111111111000;
        weights1[25840] <= 16'b1111111111110110;
        weights1[25841] <= 16'b1111111111110100;
        weights1[25842] <= 16'b1111111111111110;
        weights1[25843] <= 16'b1111111111111111;
        weights1[25844] <= 16'b1111111111111111;
        weights1[25845] <= 16'b1111111111111111;
        weights1[25846] <= 16'b1111111111111111;
        weights1[25847] <= 16'b0000000000000001;
        weights1[25848] <= 16'b1111111111111101;
        weights1[25849] <= 16'b0000000000000100;
        weights1[25850] <= 16'b0000000000000110;
        weights1[25851] <= 16'b0000000000000000;
        weights1[25852] <= 16'b1111111111110111;
        weights1[25853] <= 16'b1111111111100100;
        weights1[25854] <= 16'b1111111111101001;
        weights1[25855] <= 16'b1111111111110011;
        weights1[25856] <= 16'b1111111111110000;
        weights1[25857] <= 16'b1111111111101110;
        weights1[25858] <= 16'b1111111111101110;
        weights1[25859] <= 16'b1111111111110000;
        weights1[25860] <= 16'b1111111111101101;
        weights1[25861] <= 16'b1111111111110111;
        weights1[25862] <= 16'b1111111111110101;
        weights1[25863] <= 16'b1111111111110110;
        weights1[25864] <= 16'b1111111111111011;
        weights1[25865] <= 16'b1111111111110110;
        weights1[25866] <= 16'b1111111111111000;
        weights1[25867] <= 16'b1111111111111000;
        weights1[25868] <= 16'b1111111111111010;
        weights1[25869] <= 16'b1111111111111101;
        weights1[25870] <= 16'b1111111111111111;
        weights1[25871] <= 16'b0000000000000001;
        weights1[25872] <= 16'b0000000000000000;
        weights1[25873] <= 16'b0000000000000001;
        weights1[25874] <= 16'b0000000000000011;
        weights1[25875] <= 16'b0000000000001011;
        weights1[25876] <= 16'b0000000000001001;
        weights1[25877] <= 16'b0000000000001010;
        weights1[25878] <= 16'b0000000000001101;
        weights1[25879] <= 16'b0000000000010100;
        weights1[25880] <= 16'b0000000000000110;
        weights1[25881] <= 16'b0000000000001101;
        weights1[25882] <= 16'b0000000000001110;
        weights1[25883] <= 16'b0000000000011100;
        weights1[25884] <= 16'b0000000000001100;
        weights1[25885] <= 16'b0000000000011111;
        weights1[25886] <= 16'b0000000000010110;
        weights1[25887] <= 16'b0000000000001110;
        weights1[25888] <= 16'b0000000000001111;
        weights1[25889] <= 16'b0000000000001111;
        weights1[25890] <= 16'b0000000000010010;
        weights1[25891] <= 16'b0000000000000100;
        weights1[25892] <= 16'b0000000000000000;
        weights1[25893] <= 16'b0000000000011001;
        weights1[25894] <= 16'b1111111111111001;
        weights1[25895] <= 16'b1111111111111010;
        weights1[25896] <= 16'b1111111111111101;
        weights1[25897] <= 16'b1111111111101110;
        weights1[25898] <= 16'b1111111111111010;
        weights1[25899] <= 16'b1111111111111100;
        weights1[25900] <= 16'b0000000000000001;
        weights1[25901] <= 16'b0000000000000001;
        weights1[25902] <= 16'b0000000000000001;
        weights1[25903] <= 16'b0000000000000010;
        weights1[25904] <= 16'b0000000000001100;
        weights1[25905] <= 16'b0000000000001101;
        weights1[25906] <= 16'b0000000000000000;
        weights1[25907] <= 16'b0000000000010100;
        weights1[25908] <= 16'b1111111111111101;
        weights1[25909] <= 16'b0000000000001000;
        weights1[25910] <= 16'b0000000000001000;
        weights1[25911] <= 16'b0000000000000000;
        weights1[25912] <= 16'b0000000000000110;
        weights1[25913] <= 16'b0000000000001001;
        weights1[25914] <= 16'b1111111111111011;
        weights1[25915] <= 16'b1111111111110011;
        weights1[25916] <= 16'b1111111111111111;
        weights1[25917] <= 16'b0000000000000001;
        weights1[25918] <= 16'b0000000000000000;
        weights1[25919] <= 16'b1111111111111100;
        weights1[25920] <= 16'b0000000000000101;
        weights1[25921] <= 16'b0000000000000000;
        weights1[25922] <= 16'b0000000000000111;
        weights1[25923] <= 16'b0000000000000000;
        weights1[25924] <= 16'b0000000000000000;
        weights1[25925] <= 16'b1111111111111011;
        weights1[25926] <= 16'b1111111111110000;
        weights1[25927] <= 16'b1111111111111010;
        weights1[25928] <= 16'b0000000000000001;
        weights1[25929] <= 16'b0000000000000010;
        weights1[25930] <= 16'b1111111111111101;
        weights1[25931] <= 16'b1111111111111110;
        weights1[25932] <= 16'b0000000000001011;
        weights1[25933] <= 16'b0000000000001001;
        weights1[25934] <= 16'b0000000000001000;
        weights1[25935] <= 16'b0000000000000011;
        weights1[25936] <= 16'b1111111111110010;
        weights1[25937] <= 16'b1111111111111000;
        weights1[25938] <= 16'b0000000000000001;
        weights1[25939] <= 16'b1111111111110011;
        weights1[25940] <= 16'b1111111111111110;
        weights1[25941] <= 16'b1111111111110001;
        weights1[25942] <= 16'b0000000000001110;
        weights1[25943] <= 16'b1111111111110011;
        weights1[25944] <= 16'b0000000000000010;
        weights1[25945] <= 16'b0000000000001000;
        weights1[25946] <= 16'b1111111111110010;
        weights1[25947] <= 16'b1111111111111000;
        weights1[25948] <= 16'b1111111111101111;
        weights1[25949] <= 16'b1111111111111010;
        weights1[25950] <= 16'b0000000000001100;
        weights1[25951] <= 16'b1111111111110100;
        weights1[25952] <= 16'b1111111111111101;
        weights1[25953] <= 16'b1111111111111001;
        weights1[25954] <= 16'b1111111111111001;
        weights1[25955] <= 16'b1111111111110010;
        weights1[25956] <= 16'b1111111111111111;
        weights1[25957] <= 16'b0000000000000001;
        weights1[25958] <= 16'b0000000000000000;
        weights1[25959] <= 16'b0000000000000100;
        weights1[25960] <= 16'b0000000000010011;
        weights1[25961] <= 16'b0000000000000001;
        weights1[25962] <= 16'b0000000000000111;
        weights1[25963] <= 16'b1111111111111000;
        weights1[25964] <= 16'b1111111111110000;
        weights1[25965] <= 16'b0000000000000000;
        weights1[25966] <= 16'b0000000000000010;
        weights1[25967] <= 16'b0000000000000101;
        weights1[25968] <= 16'b0000000000000100;
        weights1[25969] <= 16'b0000000000001110;
        weights1[25970] <= 16'b1111111111111110;
        weights1[25971] <= 16'b0000000000001000;
        weights1[25972] <= 16'b0000000000000001;
        weights1[25973] <= 16'b1111111111111100;
        weights1[25974] <= 16'b1111111111111100;
        weights1[25975] <= 16'b0000000000001110;
        weights1[25976] <= 16'b1111111111111101;
        weights1[25977] <= 16'b1111111111111100;
        weights1[25978] <= 16'b1111111111111001;
        weights1[25979] <= 16'b0000000000001100;
        weights1[25980] <= 16'b1111111111111100;
        weights1[25981] <= 16'b1111111111111001;
        weights1[25982] <= 16'b1111111111101100;
        weights1[25983] <= 16'b1111111111110010;
        weights1[25984] <= 16'b1111111111111101;
        weights1[25985] <= 16'b1111111111111100;
        weights1[25986] <= 16'b1111111111111100;
        weights1[25987] <= 16'b1111111111110100;
        weights1[25988] <= 16'b0000000000001100;
        weights1[25989] <= 16'b0000000000000111;
        weights1[25990] <= 16'b1111111111111000;
        weights1[25991] <= 16'b1111111111110001;
        weights1[25992] <= 16'b1111111111110011;
        weights1[25993] <= 16'b1111111111101101;
        weights1[25994] <= 16'b1111111111111110;
        weights1[25995] <= 16'b1111111111101100;
        weights1[25996] <= 16'b1111111111101011;
        weights1[25997] <= 16'b1111111111111110;
        weights1[25998] <= 16'b1111111111110001;
        weights1[25999] <= 16'b1111111111111101;
        weights1[26000] <= 16'b1111111111110000;
        weights1[26001] <= 16'b1111111111110110;
        weights1[26002] <= 16'b1111111111111110;
        weights1[26003] <= 16'b1111111111101111;
        weights1[26004] <= 16'b1111111111101010;
        weights1[26005] <= 16'b1111111111110101;
        weights1[26006] <= 16'b1111111111111110;
        weights1[26007] <= 16'b1111111111110001;
        weights1[26008] <= 16'b1111111111101000;
        weights1[26009] <= 16'b1111111111110100;
        weights1[26010] <= 16'b1111111111101100;
        weights1[26011] <= 16'b1111111111101001;
        weights1[26012] <= 16'b1111111111111000;
        weights1[26013] <= 16'b1111111111110010;
        weights1[26014] <= 16'b1111111111110101;
        weights1[26015] <= 16'b1111111111110111;
        weights1[26016] <= 16'b1111111111110010;
        weights1[26017] <= 16'b1111111111110110;
        weights1[26018] <= 16'b1111111111111111;
        weights1[26019] <= 16'b1111111111011011;
        weights1[26020] <= 16'b1111111111100101;
        weights1[26021] <= 16'b1111111111101110;
        weights1[26022] <= 16'b1111111111101111;
        weights1[26023] <= 16'b1111111111011010;
        weights1[26024] <= 16'b1111111111111011;
        weights1[26025] <= 16'b1111111111101111;
        weights1[26026] <= 16'b0000000000000001;
        weights1[26027] <= 16'b1111111111110111;
        weights1[26028] <= 16'b0000000000000111;
        weights1[26029] <= 16'b0000000000000001;
        weights1[26030] <= 16'b0000000000000111;
        weights1[26031] <= 16'b1111111111110011;
        weights1[26032] <= 16'b1111111111111101;
        weights1[26033] <= 16'b0000000000000010;
        weights1[26034] <= 16'b1111111111111000;
        weights1[26035] <= 16'b1111111111101100;
        weights1[26036] <= 16'b1111111111110011;
        weights1[26037] <= 16'b1111111111110100;
        weights1[26038] <= 16'b1111111111101110;
        weights1[26039] <= 16'b1111111111100101;
        weights1[26040] <= 16'b1111111111111000;
        weights1[26041] <= 16'b1111111111110011;
        weights1[26042] <= 16'b1111111111101001;
        weights1[26043] <= 16'b1111111111011111;
        weights1[26044] <= 16'b1111111111110011;
        weights1[26045] <= 16'b0000000000001110;
        weights1[26046] <= 16'b1111111111111010;
        weights1[26047] <= 16'b1111111111101100;
        weights1[26048] <= 16'b1111111111101011;
        weights1[26049] <= 16'b1111111111110101;
        weights1[26050] <= 16'b1111111111100111;
        weights1[26051] <= 16'b1111111111111000;
        weights1[26052] <= 16'b1111111111100001;
        weights1[26053] <= 16'b1111111111110011;
        weights1[26054] <= 16'b1111111111010001;
        weights1[26055] <= 16'b1111111111101001;
        weights1[26056] <= 16'b1111111111101110;
        weights1[26057] <= 16'b1111111111101000;
        weights1[26058] <= 16'b1111111111110010;
        weights1[26059] <= 16'b1111111111011100;
        weights1[26060] <= 16'b1111111111110111;
        weights1[26061] <= 16'b1111111111100001;
        weights1[26062] <= 16'b1111111111101101;
        weights1[26063] <= 16'b1111111111110001;
        weights1[26064] <= 16'b1111111111111000;
        weights1[26065] <= 16'b1111111111110100;
        weights1[26066] <= 16'b1111111111100100;
        weights1[26067] <= 16'b1111111111010001;
        weights1[26068] <= 16'b1111111111110011;
        weights1[26069] <= 16'b1111111111100101;
        weights1[26070] <= 16'b1111111111101001;
        weights1[26071] <= 16'b1111111111100101;
        weights1[26072] <= 16'b1111111111100111;
        weights1[26073] <= 16'b0000000000010001;
        weights1[26074] <= 16'b1111111111100110;
        weights1[26075] <= 16'b1111111111101110;
        weights1[26076] <= 16'b1111111111101000;
        weights1[26077] <= 16'b0000000000001010;
        weights1[26078] <= 16'b1111111111100011;
        weights1[26079] <= 16'b1111111111101101;
        weights1[26080] <= 16'b1111111111110001;
        weights1[26081] <= 16'b1111111111010011;
        weights1[26082] <= 16'b1111111111101110;
        weights1[26083] <= 16'b1111111111111100;
        weights1[26084] <= 16'b1111111111101011;
        weights1[26085] <= 16'b1111111111110110;
        weights1[26086] <= 16'b1111111111011001;
        weights1[26087] <= 16'b1111111111100101;
        weights1[26088] <= 16'b1111111111010010;
        weights1[26089] <= 16'b1111111111010010;
        weights1[26090] <= 16'b1111111111101111;
        weights1[26091] <= 16'b1111111111100000;
        weights1[26092] <= 16'b1111111111101011;
        weights1[26093] <= 16'b1111111111010111;
        weights1[26094] <= 16'b1111111111100001;
        weights1[26095] <= 16'b1111111111010100;
        weights1[26096] <= 16'b1111111111111000;
        weights1[26097] <= 16'b1111111111100110;
        weights1[26098] <= 16'b1111111111011010;
        weights1[26099] <= 16'b1111111111011110;
        weights1[26100] <= 16'b1111111111010110;
        weights1[26101] <= 16'b1111111111011000;
        weights1[26102] <= 16'b1111111111011110;
        weights1[26103] <= 16'b1111111111100100;
        weights1[26104] <= 16'b1111111111010110;
        weights1[26105] <= 16'b1111111111110001;
        weights1[26106] <= 16'b1111111111110010;
        weights1[26107] <= 16'b1111111111101011;
        weights1[26108] <= 16'b1111111111100100;
        weights1[26109] <= 16'b1111111111110000;
        weights1[26110] <= 16'b1111111111100010;
        weights1[26111] <= 16'b1111111111101100;
        weights1[26112] <= 16'b1111111111101011;
        weights1[26113] <= 16'b1111111111110000;
        weights1[26114] <= 16'b1111111111101111;
        weights1[26115] <= 16'b1111111111100010;
        weights1[26116] <= 16'b1111111111011110;
        weights1[26117] <= 16'b1111111111010101;
        weights1[26118] <= 16'b1111111111010011;
        weights1[26119] <= 16'b1111111111100110;
        weights1[26120] <= 16'b1111111111100111;
        weights1[26121] <= 16'b1111111111010110;
        weights1[26122] <= 16'b1111111111101000;
        weights1[26123] <= 16'b1111111111011011;
        weights1[26124] <= 16'b1111111111111010;
        weights1[26125] <= 16'b1111111111101111;
        weights1[26126] <= 16'b1111111111011000;
        weights1[26127] <= 16'b1111111111011010;
        weights1[26128] <= 16'b1111111111100101;
        weights1[26129] <= 16'b1111111111001101;
        weights1[26130] <= 16'b1111111111000001;
        weights1[26131] <= 16'b1111111111100001;
        weights1[26132] <= 16'b1111111111011010;
        weights1[26133] <= 16'b1111111111011010;
        weights1[26134] <= 16'b1111111111011111;
        weights1[26135] <= 16'b1111111111100101;
        weights1[26136] <= 16'b1111111111010101;
        weights1[26137] <= 16'b1111111111101000;
        weights1[26138] <= 16'b1111111111100010;
        weights1[26139] <= 16'b1111111111110100;
        weights1[26140] <= 16'b1111111111100011;
        weights1[26141] <= 16'b1111111111100110;
        weights1[26142] <= 16'b1111111111011111;
        weights1[26143] <= 16'b1111111111010111;
        weights1[26144] <= 16'b1111111111110000;
        weights1[26145] <= 16'b1111111111110110;
        weights1[26146] <= 16'b1111111111101011;
        weights1[26147] <= 16'b1111111111011010;
        weights1[26148] <= 16'b1111111111100100;
        weights1[26149] <= 16'b1111111111001010;
        weights1[26150] <= 16'b1111111111011101;
        weights1[26151] <= 16'b1111111111011011;
        weights1[26152] <= 16'b1111111111110100;
        weights1[26153] <= 16'b1111111111110001;
        weights1[26154] <= 16'b1111111111011101;
        weights1[26155] <= 16'b1111111111010101;
        weights1[26156] <= 16'b1111111111001011;
        weights1[26157] <= 16'b1111111111101111;
        weights1[26158] <= 16'b1111111111110011;
        weights1[26159] <= 16'b1111111111111011;
        weights1[26160] <= 16'b1111111111110001;
        weights1[26161] <= 16'b0000000000000000;
        weights1[26162] <= 16'b1111111111110000;
        weights1[26163] <= 16'b1111111111101111;
        weights1[26164] <= 16'b1111111111110011;
        weights1[26165] <= 16'b1111111111110010;
        weights1[26166] <= 16'b1111111111100111;
        weights1[26167] <= 16'b1111111111100110;
        weights1[26168] <= 16'b1111111111110011;
        weights1[26169] <= 16'b1111111111111011;
        weights1[26170] <= 16'b1111111111110111;
        weights1[26171] <= 16'b1111111111111010;
        weights1[26172] <= 16'b1111111111111000;
        weights1[26173] <= 16'b1111111111110111;
        weights1[26174] <= 16'b1111111111111110;
        weights1[26175] <= 16'b1111111111010111;
        weights1[26176] <= 16'b1111111111010111;
        weights1[26177] <= 16'b1111111111010000;
        weights1[26178] <= 16'b1111111111010110;
        weights1[26179] <= 16'b1111111111011000;
        weights1[26180] <= 16'b1111111111111100;
        weights1[26181] <= 16'b0000000000000100;
        weights1[26182] <= 16'b1111111111110001;
        weights1[26183] <= 16'b1111111111110000;
        weights1[26184] <= 16'b0000000000011110;
        weights1[26185] <= 16'b0000000000101100;
        weights1[26186] <= 16'b0000000000001101;
        weights1[26187] <= 16'b1111111111111101;
        weights1[26188] <= 16'b0000000000010000;
        weights1[26189] <= 16'b0000000000001100;
        weights1[26190] <= 16'b0000000000000101;
        weights1[26191] <= 16'b0000000000001010;
        weights1[26192] <= 16'b0000000000001000;
        weights1[26193] <= 16'b0000000000000001;
        weights1[26194] <= 16'b0000000000000010;
        weights1[26195] <= 16'b1111111111110111;
        weights1[26196] <= 16'b0000000000010000;
        weights1[26197] <= 16'b1111111111110000;
        weights1[26198] <= 16'b1111111111101101;
        weights1[26199] <= 16'b1111111111110110;
        weights1[26200] <= 16'b1111111111111001;
        weights1[26201] <= 16'b0000000000000011;
        weights1[26202] <= 16'b1111111111011100;
        weights1[26203] <= 16'b1111111111100100;
        weights1[26204] <= 16'b1111111111101110;
        weights1[26205] <= 16'b1111111111110110;
        weights1[26206] <= 16'b1111111111010011;
        weights1[26207] <= 16'b1111111111111010;
        weights1[26208] <= 16'b0000000000000110;
        weights1[26209] <= 16'b0000000000010001;
        weights1[26210] <= 16'b0000000000011001;
        weights1[26211] <= 16'b0000000000010000;
        weights1[26212] <= 16'b0000000000010111;
        weights1[26213] <= 16'b0000000000000111;
        weights1[26214] <= 16'b0000000000011101;
        weights1[26215] <= 16'b0000000000010111;
        weights1[26216] <= 16'b0000000001000000;
        weights1[26217] <= 16'b0000000000010101;
        weights1[26218] <= 16'b0000000000100101;
        weights1[26219] <= 16'b0000000000100010;
        weights1[26220] <= 16'b0000000000011001;
        weights1[26221] <= 16'b0000000000001000;
        weights1[26222] <= 16'b0000000000001000;
        weights1[26223] <= 16'b0000000000001011;
        weights1[26224] <= 16'b0000000000011100;
        weights1[26225] <= 16'b0000000000010000;
        weights1[26226] <= 16'b1111111111111111;
        weights1[26227] <= 16'b0000000000001000;
        weights1[26228] <= 16'b1111111111110000;
        weights1[26229] <= 16'b1111111111111011;
        weights1[26230] <= 16'b0000000000010100;
        weights1[26231] <= 16'b0000000000000110;
        weights1[26232] <= 16'b1111111111101000;
        weights1[26233] <= 16'b1111111111110101;
        weights1[26234] <= 16'b1111111111111011;
        weights1[26235] <= 16'b0000000000010111;
        weights1[26236] <= 16'b0000000000010101;
        weights1[26237] <= 16'b0000000000100100;
        weights1[26238] <= 16'b0000000000011111;
        weights1[26239] <= 16'b0000000000011111;
        weights1[26240] <= 16'b0000000000001011;
        weights1[26241] <= 16'b0000000000010011;
        weights1[26242] <= 16'b0000000000100001;
        weights1[26243] <= 16'b0000000000001011;
        weights1[26244] <= 16'b0000000000000000;
        weights1[26245] <= 16'b0000000000010101;
        weights1[26246] <= 16'b0000000000101010;
        weights1[26247] <= 16'b0000000000011001;
        weights1[26248] <= 16'b0000000000001100;
        weights1[26249] <= 16'b0000000000101010;
        weights1[26250] <= 16'b0000000000010110;
        weights1[26251] <= 16'b0000000000010100;
        weights1[26252] <= 16'b0000000000101100;
        weights1[26253] <= 16'b0000000000010111;
        weights1[26254] <= 16'b0000000000010011;
        weights1[26255] <= 16'b0000000000101000;
        weights1[26256] <= 16'b0000000000001011;
        weights1[26257] <= 16'b0000000000001110;
        weights1[26258] <= 16'b0000000000000100;
        weights1[26259] <= 16'b0000000000101001;
        weights1[26260] <= 16'b0000000000110111;
        weights1[26261] <= 16'b0000000000010001;
        weights1[26262] <= 16'b0000000000010000;
        weights1[26263] <= 16'b0000000000010011;
        weights1[26264] <= 16'b0000000000010000;
        weights1[26265] <= 16'b0000000000010100;
        weights1[26266] <= 16'b0000000000100001;
        weights1[26267] <= 16'b0000000000010001;
        weights1[26268] <= 16'b0000000000011001;
        weights1[26269] <= 16'b0000000000111001;
        weights1[26270] <= 16'b0000000000010000;
        weights1[26271] <= 16'b0000000000100011;
        weights1[26272] <= 16'b0000000000011001;
        weights1[26273] <= 16'b0000000000011111;
        weights1[26274] <= 16'b0000000000010011;
        weights1[26275] <= 16'b0000000000100100;
        weights1[26276] <= 16'b0000000000101000;
        weights1[26277] <= 16'b0000000000011001;
        weights1[26278] <= 16'b0000000000100000;
        weights1[26279] <= 16'b0000000000100001;
        weights1[26280] <= 16'b0000000000101101;
        weights1[26281] <= 16'b0000000000100001;
        weights1[26282] <= 16'b0000000000010011;
        weights1[26283] <= 16'b0000000000100111;
        weights1[26284] <= 16'b0000000000100001;
        weights1[26285] <= 16'b0000000000010111;
        weights1[26286] <= 16'b0000000000110000;
        weights1[26287] <= 16'b0000000000100111;
        weights1[26288] <= 16'b0000000000011010;
        weights1[26289] <= 16'b0000000000101111;
        weights1[26290] <= 16'b0000000000011111;
        weights1[26291] <= 16'b0000000000010000;
        weights1[26292] <= 16'b0000000000001111;
        weights1[26293] <= 16'b0000000000011101;
        weights1[26294] <= 16'b0000000000010011;
        weights1[26295] <= 16'b0000000000100011;
        weights1[26296] <= 16'b0000000000001010;
        weights1[26297] <= 16'b1111111111111100;
        weights1[26298] <= 16'b0000000000010111;
        weights1[26299] <= 16'b0000000000011001;
        weights1[26300] <= 16'b0000000000011010;
        weights1[26301] <= 16'b0000000000010110;
        weights1[26302] <= 16'b0000000000011001;
        weights1[26303] <= 16'b0000000000100001;
        weights1[26304] <= 16'b0000000000011010;
        weights1[26305] <= 16'b0000000000001001;
        weights1[26306] <= 16'b0000000000001011;
        weights1[26307] <= 16'b0000000000101001;
        weights1[26308] <= 16'b0000000000011010;
        weights1[26309] <= 16'b0000000000101001;
        weights1[26310] <= 16'b0000000000000110;
        weights1[26311] <= 16'b0000000000101101;
        weights1[26312] <= 16'b0000000000010000;
        weights1[26313] <= 16'b0000000000010011;
        weights1[26314] <= 16'b0000000000011110;
        weights1[26315] <= 16'b0000000000100100;
        weights1[26316] <= 16'b0000000000011001;
        weights1[26317] <= 16'b0000000000101101;
        weights1[26318] <= 16'b0000000001001011;
        weights1[26319] <= 16'b0000000000101000;
        weights1[26320] <= 16'b0000000000001101;
        weights1[26321] <= 16'b0000000000001101;
        weights1[26322] <= 16'b0000000000010001;
        weights1[26323] <= 16'b0000000000010011;
        weights1[26324] <= 16'b0000000000000110;
        weights1[26325] <= 16'b0000000000001111;
        weights1[26326] <= 16'b0000000000100000;
        weights1[26327] <= 16'b0000000000010001;
        weights1[26328] <= 16'b0000000000001100;
        weights1[26329] <= 16'b0000000000001000;
        weights1[26330] <= 16'b0000000000010000;
        weights1[26331] <= 16'b0000000000001110;
        weights1[26332] <= 16'b0000000000011101;
        weights1[26333] <= 16'b0000000000101001;
        weights1[26334] <= 16'b0000000000010111;
        weights1[26335] <= 16'b0000000000101101;
        weights1[26336] <= 16'b0000000000011110;
        weights1[26337] <= 16'b0000000000110111;
        weights1[26338] <= 16'b0000000000110011;
        weights1[26339] <= 16'b0000000000100000;
        weights1[26340] <= 16'b0000000000110000;
        weights1[26341] <= 16'b0000000000101001;
        weights1[26342] <= 16'b0000000000100111;
        weights1[26343] <= 16'b0000000000100110;
        weights1[26344] <= 16'b0000000000111011;
        weights1[26345] <= 16'b0000000000101101;
        weights1[26346] <= 16'b0000000000100100;
        weights1[26347] <= 16'b0000000000101101;
        weights1[26348] <= 16'b1111111111111100;
        weights1[26349] <= 16'b0000000000000000;
        weights1[26350] <= 16'b1111111111110111;
        weights1[26351] <= 16'b0000000000010100;
        weights1[26352] <= 16'b0000000000001011;
        weights1[26353] <= 16'b1111111111110100;
        weights1[26354] <= 16'b0000000000010101;
        weights1[26355] <= 16'b1111111111111100;
        weights1[26356] <= 16'b0000000000001101;
        weights1[26357] <= 16'b0000000000001010;
        weights1[26358] <= 16'b0000000000000011;
        weights1[26359] <= 16'b0000000000011101;
        weights1[26360] <= 16'b1111111111111001;
        weights1[26361] <= 16'b0000000000001110;
        weights1[26362] <= 16'b0000000000011010;
        weights1[26363] <= 16'b0000000000010011;
        weights1[26364] <= 16'b0000000000001011;
        weights1[26365] <= 16'b1111111111111101;
        weights1[26366] <= 16'b0000000000100011;
        weights1[26367] <= 16'b0000000000010000;
        weights1[26368] <= 16'b0000000000101001;
        weights1[26369] <= 16'b0000000000101100;
        weights1[26370] <= 16'b0000000000001110;
        weights1[26371] <= 16'b0000000000101100;
        weights1[26372] <= 16'b0000000000110110;
        weights1[26373] <= 16'b0000000000111010;
        weights1[26374] <= 16'b0000000000100011;
        weights1[26375] <= 16'b0000000000011010;
        weights1[26376] <= 16'b0000000000000001;
        weights1[26377] <= 16'b1111111111111100;
        weights1[26378] <= 16'b1111111111011011;
        weights1[26379] <= 16'b0000000000000100;
        weights1[26380] <= 16'b0000000000000000;
        weights1[26381] <= 16'b1111111111100111;
        weights1[26382] <= 16'b1111111111110111;
        weights1[26383] <= 16'b1111111111101111;
        weights1[26384] <= 16'b0000000000000100;
        weights1[26385] <= 16'b0000000000010000;
        weights1[26386] <= 16'b0000000000001100;
        weights1[26387] <= 16'b1111111111110011;
        weights1[26388] <= 16'b0000000000000011;
        weights1[26389] <= 16'b1111111111110111;
        weights1[26390] <= 16'b1111111111111110;
        weights1[26391] <= 16'b1111111111101111;
        weights1[26392] <= 16'b1111111111111101;
        weights1[26393] <= 16'b0000000000001000;
        weights1[26394] <= 16'b0000000000001100;
        weights1[26395] <= 16'b1111111111110011;
        weights1[26396] <= 16'b0000000000100110;
        weights1[26397] <= 16'b0000000000010010;
        weights1[26398] <= 16'b0000000000100010;
        weights1[26399] <= 16'b0000000000011110;
        weights1[26400] <= 16'b0000000000011000;
        weights1[26401] <= 16'b0000000000011010;
        weights1[26402] <= 16'b0000000000000110;
        weights1[26403] <= 16'b0000000000000111;
        weights1[26404] <= 16'b1111111111111001;
        weights1[26405] <= 16'b1111111111101110;
        weights1[26406] <= 16'b1111111111100110;
        weights1[26407] <= 16'b1111111111100100;
        weights1[26408] <= 16'b0000000000000110;
        weights1[26409] <= 16'b1111111111011111;
        weights1[26410] <= 16'b0000000000000100;
        weights1[26411] <= 16'b0000000000001111;
        weights1[26412] <= 16'b1111111111101111;
        weights1[26413] <= 16'b1111111111100000;
        weights1[26414] <= 16'b1111111111111100;
        weights1[26415] <= 16'b0000000000000001;
        weights1[26416] <= 16'b1111111111111110;
        weights1[26417] <= 16'b1111111111101111;
        weights1[26418] <= 16'b1111111111101001;
        weights1[26419] <= 16'b1111111111111000;
        weights1[26420] <= 16'b1111111111110110;
        weights1[26421] <= 16'b1111111111110100;
        weights1[26422] <= 16'b1111111111100110;
        weights1[26423] <= 16'b1111111111100101;
        weights1[26424] <= 16'b1111111111111110;
        weights1[26425] <= 16'b0000000000000101;
        weights1[26426] <= 16'b0000000000000000;
        weights1[26427] <= 16'b0000000000010100;
        weights1[26428] <= 16'b0000000000010010;
        weights1[26429] <= 16'b1111111111100001;
        weights1[26430] <= 16'b1111111111111101;
        weights1[26431] <= 16'b1111111111111111;
        weights1[26432] <= 16'b1111111111110111;
        weights1[26433] <= 16'b1111111111011101;
        weights1[26434] <= 16'b1111111111011010;
        weights1[26435] <= 16'b1111111111001011;
        weights1[26436] <= 16'b1111111111101010;
        weights1[26437] <= 16'b1111111111100011;
        weights1[26438] <= 16'b1111111111111010;
        weights1[26439] <= 16'b0000000000000100;
        weights1[26440] <= 16'b0000000000000011;
        weights1[26441] <= 16'b1111111111111000;
        weights1[26442] <= 16'b1111111111110011;
        weights1[26443] <= 16'b1111111111111111;
        weights1[26444] <= 16'b0000000000000011;
        weights1[26445] <= 16'b0000000000000110;
        weights1[26446] <= 16'b1111111111111010;
        weights1[26447] <= 16'b0000000000001100;
        weights1[26448] <= 16'b1111111111110100;
        weights1[26449] <= 16'b1111111111111001;
        weights1[26450] <= 16'b1111111111111001;
        weights1[26451] <= 16'b1111111111100011;
        weights1[26452] <= 16'b1111111111011001;
        weights1[26453] <= 16'b1111111111100010;
        weights1[26454] <= 16'b1111111111100110;
        weights1[26455] <= 16'b1111111111100001;
        weights1[26456] <= 16'b1111111111010010;
        weights1[26457] <= 16'b1111111111000000;
        weights1[26458] <= 16'b1111111111010010;
        weights1[26459] <= 16'b1111111111011110;
        weights1[26460] <= 16'b1111111111111100;
        weights1[26461] <= 16'b1111111111110101;
        weights1[26462] <= 16'b1111111111100110;
        weights1[26463] <= 16'b1111111111001001;
        weights1[26464] <= 16'b1111111111000101;
        weights1[26465] <= 16'b1111111111000101;
        weights1[26466] <= 16'b1111111111011100;
        weights1[26467] <= 16'b1111111111110011;
        weights1[26468] <= 16'b1111111111111010;
        weights1[26469] <= 16'b1111111111100110;
        weights1[26470] <= 16'b1111111111111000;
        weights1[26471] <= 16'b1111111111110111;
        weights1[26472] <= 16'b0000000000100111;
        weights1[26473] <= 16'b0000000000010101;
        weights1[26474] <= 16'b0000000000000100;
        weights1[26475] <= 16'b1111111111111011;
        weights1[26476] <= 16'b1111111111011110;
        weights1[26477] <= 16'b1111111111111011;
        weights1[26478] <= 16'b1111111111110000;
        weights1[26479] <= 16'b1111111111100101;
        weights1[26480] <= 16'b1111111111010111;
        weights1[26481] <= 16'b1111111111010011;
        weights1[26482] <= 16'b1111111110111101;
        weights1[26483] <= 16'b1111111110111110;
        weights1[26484] <= 16'b1111111110100111;
        weights1[26485] <= 16'b1111111110110111;
        weights1[26486] <= 16'b1111111111000100;
        weights1[26487] <= 16'b1111111111011001;
        weights1[26488] <= 16'b1111111111111001;
        weights1[26489] <= 16'b1111111111111000;
        weights1[26490] <= 16'b1111111111101100;
        weights1[26491] <= 16'b1111111111011001;
        weights1[26492] <= 16'b1111111111010000;
        weights1[26493] <= 16'b1111111111000010;
        weights1[26494] <= 16'b1111111111001110;
        weights1[26495] <= 16'b1111111110111101;
        weights1[26496] <= 16'b1111111111011001;
        weights1[26497] <= 16'b1111111111001010;
        weights1[26498] <= 16'b0000000000000000;
        weights1[26499] <= 16'b1111111111100001;
        weights1[26500] <= 16'b1111111111100011;
        weights1[26501] <= 16'b1111111111101001;
        weights1[26502] <= 16'b1111111111100001;
        weights1[26503] <= 16'b1111111111101000;
        weights1[26504] <= 16'b1111111111110011;
        weights1[26505] <= 16'b1111111111100001;
        weights1[26506] <= 16'b1111111111110100;
        weights1[26507] <= 16'b1111111111011000;
        weights1[26508] <= 16'b1111111111010111;
        weights1[26509] <= 16'b1111111111000111;
        weights1[26510] <= 16'b1111111110110000;
        weights1[26511] <= 16'b1111111110100101;
        weights1[26512] <= 16'b1111111110101000;
        weights1[26513] <= 16'b1111111110111111;
        weights1[26514] <= 16'b1111111111010100;
        weights1[26515] <= 16'b1111111111011010;
        weights1[26516] <= 16'b1111111111111011;
        weights1[26517] <= 16'b1111111111110011;
        weights1[26518] <= 16'b1111111111101100;
        weights1[26519] <= 16'b1111111111010111;
        weights1[26520] <= 16'b1111111111000100;
        weights1[26521] <= 16'b1111111110111011;
        weights1[26522] <= 16'b1111111110111001;
        weights1[26523] <= 16'b1111111110100011;
        weights1[26524] <= 16'b1111111110110100;
        weights1[26525] <= 16'b1111111110001110;
        weights1[26526] <= 16'b1111111110101101;
        weights1[26527] <= 16'b1111111110100101;
        weights1[26528] <= 16'b1111111110111001;
        weights1[26529] <= 16'b1111111111010011;
        weights1[26530] <= 16'b1111111111001001;
        weights1[26531] <= 16'b1111111111101000;
        weights1[26532] <= 16'b1111111111011000;
        weights1[26533] <= 16'b1111111111001110;
        weights1[26534] <= 16'b1111111111011001;
        weights1[26535] <= 16'b1111111111011101;
        weights1[26536] <= 16'b1111111111011001;
        weights1[26537] <= 16'b1111111110110110;
        weights1[26538] <= 16'b1111111111000010;
        weights1[26539] <= 16'b1111111110110111;
        weights1[26540] <= 16'b1111111110110111;
        weights1[26541] <= 16'b1111111111010000;
        weights1[26542] <= 16'b1111111111100010;
        weights1[26543] <= 16'b1111111111100110;
        weights1[26544] <= 16'b1111111111111101;
        weights1[26545] <= 16'b1111111111110110;
        weights1[26546] <= 16'b1111111111100101;
        weights1[26547] <= 16'b1111111111011000;
        weights1[26548] <= 16'b1111111111010101;
        weights1[26549] <= 16'b1111111111001101;
        weights1[26550] <= 16'b1111111111000001;
        weights1[26551] <= 16'b1111111110110111;
        weights1[26552] <= 16'b1111111110110100;
        weights1[26553] <= 16'b1111111111000101;
        weights1[26554] <= 16'b1111111110101000;
        weights1[26555] <= 16'b1111111111010101;
        weights1[26556] <= 16'b1111111111000111;
        weights1[26557] <= 16'b1111111110110110;
        weights1[26558] <= 16'b1111111111011110;
        weights1[26559] <= 16'b1111111111011001;
        weights1[26560] <= 16'b1111111111010101;
        weights1[26561] <= 16'b1111111111010000;
        weights1[26562] <= 16'b1111111111011100;
        weights1[26563] <= 16'b1111111111000111;
        weights1[26564] <= 16'b1111111110100111;
        weights1[26565] <= 16'b1111111110111110;
        weights1[26566] <= 16'b1111111110111111;
        weights1[26567] <= 16'b1111111111010011;
        weights1[26568] <= 16'b1111111111010101;
        weights1[26569] <= 16'b1111111111011101;
        weights1[26570] <= 16'b1111111111100001;
        weights1[26571] <= 16'b1111111111100111;
        weights1[26572] <= 16'b0000000000000000;
        weights1[26573] <= 16'b1111111111110101;
        weights1[26574] <= 16'b1111111111100111;
        weights1[26575] <= 16'b1111111111100011;
        weights1[26576] <= 16'b1111111111100000;
        weights1[26577] <= 16'b1111111111010000;
        weights1[26578] <= 16'b1111111111000100;
        weights1[26579] <= 16'b1111111111000011;
        weights1[26580] <= 16'b1111111110111111;
        weights1[26581] <= 16'b1111111110011100;
        weights1[26582] <= 16'b1111111110011101;
        weights1[26583] <= 16'b1111111110100110;
        weights1[26584] <= 16'b1111111110001001;
        weights1[26585] <= 16'b1111111110010000;
        weights1[26586] <= 16'b1111111110101101;
        weights1[26587] <= 16'b1111111110010101;
        weights1[26588] <= 16'b1111111110010100;
        weights1[26589] <= 16'b1111111110011001;
        weights1[26590] <= 16'b1111111110000100;
        weights1[26591] <= 16'b1111111110010100;
        weights1[26592] <= 16'b1111111110010111;
        weights1[26593] <= 16'b1111111110110011;
        weights1[26594] <= 16'b1111111110111101;
        weights1[26595] <= 16'b1111111111010100;
        weights1[26596] <= 16'b1111111111011000;
        weights1[26597] <= 16'b1111111111100101;
        weights1[26598] <= 16'b1111111111101000;
        weights1[26599] <= 16'b1111111111110001;
        weights1[26600] <= 16'b1111111111111110;
        weights1[26601] <= 16'b1111111111111001;
        weights1[26602] <= 16'b1111111111110011;
        weights1[26603] <= 16'b1111111111110000;
        weights1[26604] <= 16'b1111111111101000;
        weights1[26605] <= 16'b1111111111011000;
        weights1[26606] <= 16'b1111111111001010;
        weights1[26607] <= 16'b1111111111000001;
        weights1[26608] <= 16'b1111111110111111;
        weights1[26609] <= 16'b1111111110111010;
        weights1[26610] <= 16'b1111111110110000;
        weights1[26611] <= 16'b1111111110011110;
        weights1[26612] <= 16'b1111111110011001;
        weights1[26613] <= 16'b1111111110001010;
        weights1[26614] <= 16'b1111111110001001;
        weights1[26615] <= 16'b1111111110010000;
        weights1[26616] <= 16'b1111111110011100;
        weights1[26617] <= 16'b1111111110010010;
        weights1[26618] <= 16'b1111111110101000;
        weights1[26619] <= 16'b1111111110101110;
        weights1[26620] <= 16'b1111111110110001;
        weights1[26621] <= 16'b1111111111000110;
        weights1[26622] <= 16'b1111111111010001;
        weights1[26623] <= 16'b1111111111100010;
        weights1[26624] <= 16'b1111111111100101;
        weights1[26625] <= 16'b1111111111101001;
        weights1[26626] <= 16'b1111111111110000;
        weights1[26627] <= 16'b1111111111110111;
        weights1[26628] <= 16'b1111111111111011;
        weights1[26629] <= 16'b1111111111111010;
        weights1[26630] <= 16'b1111111111111010;
        weights1[26631] <= 16'b1111111111111001;
        weights1[26632] <= 16'b1111111111110000;
        weights1[26633] <= 16'b1111111111101000;
        weights1[26634] <= 16'b1111111111100001;
        weights1[26635] <= 16'b1111111111001101;
        weights1[26636] <= 16'b1111111111001000;
        weights1[26637] <= 16'b1111111111001101;
        weights1[26638] <= 16'b1111111111000101;
        weights1[26639] <= 16'b1111111110110010;
        weights1[26640] <= 16'b1111111110110011;
        weights1[26641] <= 16'b1111111110110000;
        weights1[26642] <= 16'b1111111110100110;
        weights1[26643] <= 16'b1111111110111000;
        weights1[26644] <= 16'b1111111110111101;
        weights1[26645] <= 16'b1111111110111101;
        weights1[26646] <= 16'b1111111111000101;
        weights1[26647] <= 16'b1111111111001101;
        weights1[26648] <= 16'b1111111111010001;
        weights1[26649] <= 16'b1111111111010110;
        weights1[26650] <= 16'b1111111111100100;
        weights1[26651] <= 16'b1111111111101101;
        weights1[26652] <= 16'b1111111111101101;
        weights1[26653] <= 16'b1111111111110100;
        weights1[26654] <= 16'b1111111111111001;
        weights1[26655] <= 16'b1111111111111100;
        weights1[26656] <= 16'b0000000000000001;
        weights1[26657] <= 16'b1111111111111111;
        weights1[26658] <= 16'b1111111111111110;
        weights1[26659] <= 16'b0000000000000001;
        weights1[26660] <= 16'b0000000000000011;
        weights1[26661] <= 16'b0000000000001000;
        weights1[26662] <= 16'b0000000000000001;
        weights1[26663] <= 16'b0000000000001101;
        weights1[26664] <= 16'b0000000000010110;
        weights1[26665] <= 16'b0000000000001110;
        weights1[26666] <= 16'b0000000000000111;
        weights1[26667] <= 16'b0000000000000101;
        weights1[26668] <= 16'b1111111111110011;
        weights1[26669] <= 16'b1111111111011000;
        weights1[26670] <= 16'b1111111111000001;
        weights1[26671] <= 16'b1111111111000011;
        weights1[26672] <= 16'b1111111111010110;
        weights1[26673] <= 16'b1111111111011101;
        weights1[26674] <= 16'b1111111111110100;
        weights1[26675] <= 16'b1111111111111110;
        weights1[26676] <= 16'b0000000000010000;
        weights1[26677] <= 16'b0000000000011000;
        weights1[26678] <= 16'b0000000000010000;
        weights1[26679] <= 16'b0000000000010010;
        weights1[26680] <= 16'b0000000000001010;
        weights1[26681] <= 16'b0000000000000010;
        weights1[26682] <= 16'b0000000000000110;
        weights1[26683] <= 16'b0000000000000001;
        weights1[26684] <= 16'b1111111111111110;
        weights1[26685] <= 16'b1111111111111110;
        weights1[26686] <= 16'b0000000000000001;
        weights1[26687] <= 16'b0000000000000010;
        weights1[26688] <= 16'b0000000000000101;
        weights1[26689] <= 16'b0000000000000010;
        weights1[26690] <= 16'b1111111111111110;
        weights1[26691] <= 16'b0000000000010101;
        weights1[26692] <= 16'b0000000000100001;
        weights1[26693] <= 16'b0000000000001001;
        weights1[26694] <= 16'b0000000000010011;
        weights1[26695] <= 16'b0000000000001101;
        weights1[26696] <= 16'b0000000000010001;
        weights1[26697] <= 16'b1111111111100110;
        weights1[26698] <= 16'b1111111111001101;
        weights1[26699] <= 16'b1111111111000010;
        weights1[26700] <= 16'b1111111111001001;
        weights1[26701] <= 16'b1111111111011011;
        weights1[26702] <= 16'b1111111111011111;
        weights1[26703] <= 16'b0000000000010001;
        weights1[26704] <= 16'b0000000000011111;
        weights1[26705] <= 16'b0000000000011011;
        weights1[26706] <= 16'b0000000000010101;
        weights1[26707] <= 16'b0000000000010100;
        weights1[26708] <= 16'b0000000000001100;
        weights1[26709] <= 16'b0000000000010001;
        weights1[26710] <= 16'b0000000000001111;
        weights1[26711] <= 16'b0000000000001001;
        weights1[26712] <= 16'b0000000000000010;
        weights1[26713] <= 16'b0000000000000010;
        weights1[26714] <= 16'b0000000000000010;
        weights1[26715] <= 16'b0000000000000010;
        weights1[26716] <= 16'b0000000000000100;
        weights1[26717] <= 16'b1111111111111101;
        weights1[26718] <= 16'b1111111111110010;
        weights1[26719] <= 16'b0000000000000000;
        weights1[26720] <= 16'b0000000000011001;
        weights1[26721] <= 16'b0000000000001100;
        weights1[26722] <= 16'b1111111111110011;
        weights1[26723] <= 16'b0000000000000011;
        weights1[26724] <= 16'b0000000000000110;
        weights1[26725] <= 16'b1111111111010101;
        weights1[26726] <= 16'b1111111111000001;
        weights1[26727] <= 16'b1111111110101111;
        weights1[26728] <= 16'b1111111110101101;
        weights1[26729] <= 16'b1111111110111001;
        weights1[26730] <= 16'b1111111111010000;
        weights1[26731] <= 16'b0000000000000101;
        weights1[26732] <= 16'b0000000000101100;
        weights1[26733] <= 16'b0000000000100100;
        weights1[26734] <= 16'b0000000000011100;
        weights1[26735] <= 16'b0000000000100000;
        weights1[26736] <= 16'b0000000000010010;
        weights1[26737] <= 16'b0000000000010000;
        weights1[26738] <= 16'b0000000000010000;
        weights1[26739] <= 16'b0000000000001010;
        weights1[26740] <= 16'b0000000000000110;
        weights1[26741] <= 16'b0000000000001001;
        weights1[26742] <= 16'b0000000000000010;
        weights1[26743] <= 16'b0000000000000101;
        weights1[26744] <= 16'b0000000000000100;
        weights1[26745] <= 16'b1111111111101111;
        weights1[26746] <= 16'b1111111111111001;
        weights1[26747] <= 16'b0000000000001011;
        weights1[26748] <= 16'b0000000000010010;
        weights1[26749] <= 16'b0000000000000111;
        weights1[26750] <= 16'b1111111111111001;
        weights1[26751] <= 16'b1111111111110101;
        weights1[26752] <= 16'b1111111111110101;
        weights1[26753] <= 16'b1111111111001110;
        weights1[26754] <= 16'b1111111111010000;
        weights1[26755] <= 16'b1111111110101011;
        weights1[26756] <= 16'b1111111110000001;
        weights1[26757] <= 16'b1111111110100110;
        weights1[26758] <= 16'b1111111111001101;
        weights1[26759] <= 16'b1111111111111100;
        weights1[26760] <= 16'b0000000000010110;
        weights1[26761] <= 16'b0000000000000101;
        weights1[26762] <= 16'b0000000000010010;
        weights1[26763] <= 16'b0000000000011000;
        weights1[26764] <= 16'b0000000000011101;
        weights1[26765] <= 16'b0000000000010000;
        weights1[26766] <= 16'b0000000000001111;
        weights1[26767] <= 16'b0000000000001001;
        weights1[26768] <= 16'b0000000000000100;
        weights1[26769] <= 16'b0000000000000011;
        weights1[26770] <= 16'b1111111111111011;
        weights1[26771] <= 16'b1111111111111100;
        weights1[26772] <= 16'b1111111111111010;
        weights1[26773] <= 16'b1111111111110111;
        weights1[26774] <= 16'b1111111111111001;
        weights1[26775] <= 16'b1111111111111100;
        weights1[26776] <= 16'b0000000000001000;
        weights1[26777] <= 16'b0000000000011001;
        weights1[26778] <= 16'b1111111111110001;
        weights1[26779] <= 16'b0000000000000100;
        weights1[26780] <= 16'b1111111111111111;
        weights1[26781] <= 16'b1111111111010010;
        weights1[26782] <= 16'b1111111111011111;
        weights1[26783] <= 16'b1111111110100011;
        weights1[26784] <= 16'b1111111101101101;
        weights1[26785] <= 16'b1111111110000001;
        weights1[26786] <= 16'b1111111110111100;
        weights1[26787] <= 16'b1111111111100101;
        weights1[26788] <= 16'b0000000000010110;
        weights1[26789] <= 16'b0000000000010101;
        weights1[26790] <= 16'b0000000000011011;
        weights1[26791] <= 16'b0000000000100001;
        weights1[26792] <= 16'b0000000000101001;
        weights1[26793] <= 16'b0000000000001001;
        weights1[26794] <= 16'b0000000000000110;
        weights1[26795] <= 16'b0000000000001100;
        weights1[26796] <= 16'b0000000000000101;
        weights1[26797] <= 16'b1111111111111101;
        weights1[26798] <= 16'b1111111111111100;
        weights1[26799] <= 16'b1111111111111000;
        weights1[26800] <= 16'b1111111111101000;
        weights1[26801] <= 16'b1111111111111010;
        weights1[26802] <= 16'b1111111111101111;
        weights1[26803] <= 16'b0000000000000000;
        weights1[26804] <= 16'b0000000000001110;
        weights1[26805] <= 16'b1111111111111000;
        weights1[26806] <= 16'b0000000000000001;
        weights1[26807] <= 16'b1111111111111011;
        weights1[26808] <= 16'b0000000000001101;
        weights1[26809] <= 16'b1111111111110101;
        weights1[26810] <= 16'b1111111111010101;
        weights1[26811] <= 16'b1111111110111001;
        weights1[26812] <= 16'b1111111101011101;
        weights1[26813] <= 16'b1111111101010011;
        weights1[26814] <= 16'b1111111111100110;
        weights1[26815] <= 16'b0000000000010000;
        weights1[26816] <= 16'b0000000000011001;
        weights1[26817] <= 16'b0000000000101001;
        weights1[26818] <= 16'b0000000000011111;
        weights1[26819] <= 16'b0000000000101101;
        weights1[26820] <= 16'b0000000000001111;
        weights1[26821] <= 16'b0000000000001001;
        weights1[26822] <= 16'b0000000000000001;
        weights1[26823] <= 16'b1111111111111111;
        weights1[26824] <= 16'b0000000000000011;
        weights1[26825] <= 16'b0000000000000010;
        weights1[26826] <= 16'b1111111111110111;
        weights1[26827] <= 16'b1111111111111001;
        weights1[26828] <= 16'b1111111111111101;
        weights1[26829] <= 16'b0000000000000000;
        weights1[26830] <= 16'b0000000000000010;
        weights1[26831] <= 16'b0000000000000010;
        weights1[26832] <= 16'b0000000000001001;
        weights1[26833] <= 16'b0000000000010010;
        weights1[26834] <= 16'b0000000000000111;
        weights1[26835] <= 16'b1111111111111001;
        weights1[26836] <= 16'b1111111111111001;
        weights1[26837] <= 16'b1111111111101010;
        weights1[26838] <= 16'b1111111111111110;
        weights1[26839] <= 16'b1111111111000111;
        weights1[26840] <= 16'b1111111100110001;
        weights1[26841] <= 16'b1111111101000100;
        weights1[26842] <= 16'b1111111111011111;
        weights1[26843] <= 16'b0000000000111001;
        weights1[26844] <= 16'b0000000000010011;
        weights1[26845] <= 16'b0000000000010000;
        weights1[26846] <= 16'b0000000000011001;
        weights1[26847] <= 16'b0000000000100010;
        weights1[26848] <= 16'b0000000000010001;
        weights1[26849] <= 16'b1111111111111101;
        weights1[26850] <= 16'b1111111111111001;
        weights1[26851] <= 16'b1111111111111101;
        weights1[26852] <= 16'b0000000000001000;
        weights1[26853] <= 16'b0000000000000110;
        weights1[26854] <= 16'b1111111111111100;
        weights1[26855] <= 16'b1111111111110110;
        weights1[26856] <= 16'b1111111111111101;
        weights1[26857] <= 16'b1111111111100101;
        weights1[26858] <= 16'b1111111111101110;
        weights1[26859] <= 16'b1111111111111110;
        weights1[26860] <= 16'b0000000000010111;
        weights1[26861] <= 16'b0000000000001100;
        weights1[26862] <= 16'b0000000000010011;
        weights1[26863] <= 16'b0000000000000000;
        weights1[26864] <= 16'b0000000000001101;
        weights1[26865] <= 16'b1111111111111111;
        weights1[26866] <= 16'b1111111111110100;
        weights1[26867] <= 16'b1111111111100001;
        weights1[26868] <= 16'b1111111100001100;
        weights1[26869] <= 16'b1111111100110111;
        weights1[26870] <= 16'b0000000000100111;
        weights1[26871] <= 16'b0000000001000110;
        weights1[26872] <= 16'b0000000000100110;
        weights1[26873] <= 16'b0000000000010001;
        weights1[26874] <= 16'b0000000000011101;
        weights1[26875] <= 16'b0000000000101110;
        weights1[26876] <= 16'b0000000000001010;
        weights1[26877] <= 16'b1111111111101100;
        weights1[26878] <= 16'b1111111111101001;
        weights1[26879] <= 16'b1111111111101101;
        weights1[26880] <= 16'b0000000000000011;
        weights1[26881] <= 16'b1111111111111111;
        weights1[26882] <= 16'b0000000000000011;
        weights1[26883] <= 16'b1111111111111101;
        weights1[26884] <= 16'b1111111111110100;
        weights1[26885] <= 16'b1111111111100110;
        weights1[26886] <= 16'b1111111111100000;
        weights1[26887] <= 16'b1111111111110111;
        weights1[26888] <= 16'b1111111111100101;
        weights1[26889] <= 16'b0000000000000111;
        weights1[26890] <= 16'b0000000000100010;
        weights1[26891] <= 16'b0000000000001110;
        weights1[26892] <= 16'b0000000000101000;
        weights1[26893] <= 16'b0000000000001000;
        weights1[26894] <= 16'b1111111111101110;
        weights1[26895] <= 16'b1111111110101011;
        weights1[26896] <= 16'b1111111011111011;
        weights1[26897] <= 16'b1111111110100101;
        weights1[26898] <= 16'b0000000000111000;
        weights1[26899] <= 16'b0000000000100000;
        weights1[26900] <= 16'b0000000000011110;
        weights1[26901] <= 16'b1111111111100110;
        weights1[26902] <= 16'b0000000000100010;
        weights1[26903] <= 16'b0000000000100011;
        weights1[26904] <= 16'b1111111111101111;
        weights1[26905] <= 16'b1111111111111001;
        weights1[26906] <= 16'b1111111111001000;
        weights1[26907] <= 16'b1111111111011111;
        weights1[26908] <= 16'b0000000000000110;
        weights1[26909] <= 16'b1111111111111111;
        weights1[26910] <= 16'b0000000000010001;
        weights1[26911] <= 16'b0000000000000001;
        weights1[26912] <= 16'b1111111111110000;
        weights1[26913] <= 16'b1111111111111101;
        weights1[26914] <= 16'b1111111111101100;
        weights1[26915] <= 16'b1111111111110100;
        weights1[26916] <= 16'b0000000000000111;
        weights1[26917] <= 16'b1111111111111110;
        weights1[26918] <= 16'b0000000000000100;
        weights1[26919] <= 16'b0000000000010110;
        weights1[26920] <= 16'b0000000000011110;
        weights1[26921] <= 16'b0000000000100100;
        weights1[26922] <= 16'b1111111111101110;
        weights1[26923] <= 16'b1111111101101100;
        weights1[26924] <= 16'b1111111011110011;
        weights1[26925] <= 16'b1111111111111001;
        weights1[26926] <= 16'b0000000000101111;
        weights1[26927] <= 16'b0000000000000101;
        weights1[26928] <= 16'b0000000000100010;
        weights1[26929] <= 16'b0000000000001000;
        weights1[26930] <= 16'b0000000000010010;
        weights1[26931] <= 16'b0000000000000011;
        weights1[26932] <= 16'b1111111111110111;
        weights1[26933] <= 16'b1111111111011001;
        weights1[26934] <= 16'b1111111111010011;
        weights1[26935] <= 16'b1111111111100001;
        weights1[26936] <= 16'b0000000000000101;
        weights1[26937] <= 16'b0000000000000111;
        weights1[26938] <= 16'b0000000000000001;
        weights1[26939] <= 16'b1111111111111001;
        weights1[26940] <= 16'b1111111111110000;
        weights1[26941] <= 16'b1111111111110111;
        weights1[26942] <= 16'b1111111111101001;
        weights1[26943] <= 16'b0000000000000011;
        weights1[26944] <= 16'b0000000000001111;
        weights1[26945] <= 16'b0000000000010000;
        weights1[26946] <= 16'b0000000000001101;
        weights1[26947] <= 16'b0000000000011000;
        weights1[26948] <= 16'b0000000000100011;
        weights1[26949] <= 16'b0000000000100110;
        weights1[26950] <= 16'b1111111111111110;
        weights1[26951] <= 16'b1111111101010100;
        weights1[26952] <= 16'b1111111101011111;
        weights1[26953] <= 16'b0000000000001111;
        weights1[26954] <= 16'b0000000000010000;
        weights1[26955] <= 16'b0000000000010011;
        weights1[26956] <= 16'b0000000000010011;
        weights1[26957] <= 16'b0000000000001111;
        weights1[26958] <= 16'b0000000000000111;
        weights1[26959] <= 16'b0000000000000000;
        weights1[26960] <= 16'b1111111111110011;
        weights1[26961] <= 16'b1111111111011011;
        weights1[26962] <= 16'b1111111111010101;
        weights1[26963] <= 16'b1111111111100100;
        weights1[26964] <= 16'b0000000000000010;
        weights1[26965] <= 16'b0000000000001010;
        weights1[26966] <= 16'b1111111111111001;
        weights1[26967] <= 16'b1111111111110100;
        weights1[26968] <= 16'b1111111111011010;
        weights1[26969] <= 16'b1111111111110011;
        weights1[26970] <= 16'b1111111111110101;
        weights1[26971] <= 16'b0000000000000000;
        weights1[26972] <= 16'b1111111111110010;
        weights1[26973] <= 16'b0000000000000000;
        weights1[26974] <= 16'b0000000000010111;
        weights1[26975] <= 16'b0000000000001110;
        weights1[26976] <= 16'b0000000000110100;
        weights1[26977] <= 16'b0000000000010100;
        weights1[26978] <= 16'b1111111111010100;
        weights1[26979] <= 16'b1111111101111101;
        weights1[26980] <= 16'b1111111110100000;
        weights1[26981] <= 16'b1111111111110110;
        weights1[26982] <= 16'b0000000000101011;
        weights1[26983] <= 16'b0000000000001101;
        weights1[26984] <= 16'b0000000000000000;
        weights1[26985] <= 16'b0000000000010111;
        weights1[26986] <= 16'b0000000000001110;
        weights1[26987] <= 16'b0000000000001001;
        weights1[26988] <= 16'b1111111111100101;
        weights1[26989] <= 16'b1111111111011010;
        weights1[26990] <= 16'b1111111111011111;
        weights1[26991] <= 16'b1111111111100101;
        weights1[26992] <= 16'b0000000000000001;
        weights1[26993] <= 16'b0000000000010100;
        weights1[26994] <= 16'b0000000000001101;
        weights1[26995] <= 16'b0000000000000010;
        weights1[26996] <= 16'b1111111111101100;
        weights1[26997] <= 16'b1111111111101011;
        weights1[26998] <= 16'b1111111111110011;
        weights1[26999] <= 16'b1111111111100100;
        weights1[27000] <= 16'b0000000000000000;
        weights1[27001] <= 16'b0000000000000101;
        weights1[27002] <= 16'b0000000000001101;
        weights1[27003] <= 16'b0000000000010101;
        weights1[27004] <= 16'b0000000000011000;
        weights1[27005] <= 16'b0000000000101110;
        weights1[27006] <= 16'b1111111111110010;
        weights1[27007] <= 16'b1111111110101100;
        weights1[27008] <= 16'b1111111111001111;
        weights1[27009] <= 16'b1111111111111101;
        weights1[27010] <= 16'b0000000000010010;
        weights1[27011] <= 16'b0000000000100101;
        weights1[27012] <= 16'b0000000000010000;
        weights1[27013] <= 16'b0000000000010011;
        weights1[27014] <= 16'b0000000000001110;
        weights1[27015] <= 16'b1111111111111000;
        weights1[27016] <= 16'b1111111111100111;
        weights1[27017] <= 16'b1111111111100000;
        weights1[27018] <= 16'b1111111111101000;
        weights1[27019] <= 16'b1111111111110000;
        weights1[27020] <= 16'b1111111111111110;
        weights1[27021] <= 16'b0000000000010000;
        weights1[27022] <= 16'b0000000000000101;
        weights1[27023] <= 16'b0000000000001011;
        weights1[27024] <= 16'b0000000000000101;
        weights1[27025] <= 16'b1111111111101011;
        weights1[27026] <= 16'b0000000000010100;
        weights1[27027] <= 16'b1111111111110011;
        weights1[27028] <= 16'b0000000000000001;
        weights1[27029] <= 16'b1111111111110110;
        weights1[27030] <= 16'b0000000000001101;
        weights1[27031] <= 16'b0000000000001000;
        weights1[27032] <= 16'b0000000000011001;
        weights1[27033] <= 16'b1111111111111011;
        weights1[27034] <= 16'b1111111111100011;
        weights1[27035] <= 16'b1111111111011110;
        weights1[27036] <= 16'b1111111111011010;
        weights1[27037] <= 16'b0000000000001101;
        weights1[27038] <= 16'b0000000000010000;
        weights1[27039] <= 16'b0000000000100000;
        weights1[27040] <= 16'b0000000000011001;
        weights1[27041] <= 16'b0000000000001001;
        weights1[27042] <= 16'b0000000000000010;
        weights1[27043] <= 16'b1111111111100010;
        weights1[27044] <= 16'b1111111111110110;
        weights1[27045] <= 16'b1111111111011100;
        weights1[27046] <= 16'b1111111111101011;
        weights1[27047] <= 16'b1111111111110000;
        weights1[27048] <= 16'b1111111111111011;
        weights1[27049] <= 16'b0000000000000011;
        weights1[27050] <= 16'b0000000000001010;
        weights1[27051] <= 16'b0000000000001100;
        weights1[27052] <= 16'b0000000000001101;
        weights1[27053] <= 16'b1111111111110000;
        weights1[27054] <= 16'b0000000000001001;
        weights1[27055] <= 16'b1111111111110001;
        weights1[27056] <= 16'b0000000000000011;
        weights1[27057] <= 16'b0000000000010100;
        weights1[27058] <= 16'b1111111111111101;
        weights1[27059] <= 16'b0000000000010000;
        weights1[27060] <= 16'b0000000000001101;
        weights1[27061] <= 16'b0000000000000001;
        weights1[27062] <= 16'b1111111111101110;
        weights1[27063] <= 16'b1111111111011011;
        weights1[27064] <= 16'b1111111111111100;
        weights1[27065] <= 16'b0000000000010001;
        weights1[27066] <= 16'b0000000000001101;
        weights1[27067] <= 16'b0000000000010010;
        weights1[27068] <= 16'b0000000000000001;
        weights1[27069] <= 16'b0000000000010101;
        weights1[27070] <= 16'b1111111111111110;
        weights1[27071] <= 16'b1111111111110110;
        weights1[27072] <= 16'b1111111111110111;
        weights1[27073] <= 16'b1111111111110101;
        weights1[27074] <= 16'b1111111111100111;
        weights1[27075] <= 16'b1111111111110000;
        weights1[27076] <= 16'b0000000000001011;
        weights1[27077] <= 16'b0000000000001101;
        weights1[27078] <= 16'b0000000000011000;
        weights1[27079] <= 16'b0000000000001101;
        weights1[27080] <= 16'b1111111111111001;
        weights1[27081] <= 16'b0000000000000101;
        weights1[27082] <= 16'b1111111111110010;
        weights1[27083] <= 16'b0000000000000101;
        weights1[27084] <= 16'b0000000000000001;
        weights1[27085] <= 16'b1111111111111101;
        weights1[27086] <= 16'b0000000000001100;
        weights1[27087] <= 16'b0000000000000101;
        weights1[27088] <= 16'b1111111111111100;
        weights1[27089] <= 16'b1111111111111011;
        weights1[27090] <= 16'b1111111111101111;
        weights1[27091] <= 16'b1111111111101001;
        weights1[27092] <= 16'b0000000000000011;
        weights1[27093] <= 16'b0000000000010010;
        weights1[27094] <= 16'b0000000000001101;
        weights1[27095] <= 16'b0000000000011001;
        weights1[27096] <= 16'b0000000000001010;
        weights1[27097] <= 16'b1111111111111111;
        weights1[27098] <= 16'b1111111111111111;
        weights1[27099] <= 16'b1111111111111000;
        weights1[27100] <= 16'b1111111111100010;
        weights1[27101] <= 16'b1111111111111110;
        weights1[27102] <= 16'b1111111111111010;
        weights1[27103] <= 16'b1111111111110010;
        weights1[27104] <= 16'b0000000000000110;
        weights1[27105] <= 16'b0000000000001011;
        weights1[27106] <= 16'b0000000000001111;
        weights1[27107] <= 16'b0000000000000110;
        weights1[27108] <= 16'b1111111111111010;
        weights1[27109] <= 16'b1111111111111010;
        weights1[27110] <= 16'b0000000000000110;
        weights1[27111] <= 16'b1111111111111111;
        weights1[27112] <= 16'b1111111111100110;
        weights1[27113] <= 16'b1111111111111011;
        weights1[27114] <= 16'b1111111111111101;
        weights1[27115] <= 16'b0000000000000100;
        weights1[27116] <= 16'b1111111111110011;
        weights1[27117] <= 16'b1111111111111010;
        weights1[27118] <= 16'b0000000000000010;
        weights1[27119] <= 16'b0000000000000111;
        weights1[27120] <= 16'b0000000000000100;
        weights1[27121] <= 16'b0000000000001000;
        weights1[27122] <= 16'b1111111111111011;
        weights1[27123] <= 16'b1111111111110101;
        weights1[27124] <= 16'b1111111111111101;
        weights1[27125] <= 16'b0000000000000001;
        weights1[27126] <= 16'b0000000000000111;
        weights1[27127] <= 16'b1111111111100011;
        weights1[27128] <= 16'b1111111111110101;
        weights1[27129] <= 16'b1111111111111110;
        weights1[27130] <= 16'b1111111111111101;
        weights1[27131] <= 16'b1111111111111000;
        weights1[27132] <= 16'b0000000000000110;
        weights1[27133] <= 16'b0000000000000001;
        weights1[27134] <= 16'b0000000000010011;
        weights1[27135] <= 16'b0000000000000110;
        weights1[27136] <= 16'b1111111111110111;
        weights1[27137] <= 16'b0000000000000010;
        weights1[27138] <= 16'b0000000000001000;
        weights1[27139] <= 16'b1111111111111000;
        weights1[27140] <= 16'b1111111111100011;
        weights1[27141] <= 16'b1111111111110101;
        weights1[27142] <= 16'b1111111111111111;
        weights1[27143] <= 16'b1111111111100111;
        weights1[27144] <= 16'b1111111111111110;
        weights1[27145] <= 16'b1111111111110001;
        weights1[27146] <= 16'b1111111111101111;
        weights1[27147] <= 16'b1111111111111011;
        weights1[27148] <= 16'b1111111111111000;
        weights1[27149] <= 16'b0000000000010001;
        weights1[27150] <= 16'b0000000000000101;
        weights1[27151] <= 16'b1111111111111100;
        weights1[27152] <= 16'b1111111111111101;
        weights1[27153] <= 16'b0000000000001101;
        weights1[27154] <= 16'b0000000000000000;
        weights1[27155] <= 16'b1111111111111100;
        weights1[27156] <= 16'b0000000000001001;
        weights1[27157] <= 16'b0000000000001111;
        weights1[27158] <= 16'b1111111111111100;
        weights1[27159] <= 16'b0000000000000001;
        weights1[27160] <= 16'b1111111111110110;
        weights1[27161] <= 16'b1111111111111011;
        weights1[27162] <= 16'b1111111111111101;
        weights1[27163] <= 16'b0000000000000100;
        weights1[27164] <= 16'b0000000000001110;
        weights1[27165] <= 16'b0000000000000000;
        weights1[27166] <= 16'b1111111111110110;
        weights1[27167] <= 16'b0000000000001000;
        weights1[27168] <= 16'b1111111111110101;
        weights1[27169] <= 16'b0000000000001101;
        weights1[27170] <= 16'b1111111111111111;
        weights1[27171] <= 16'b0000000000000010;
        weights1[27172] <= 16'b1111111111111111;
        weights1[27173] <= 16'b0000000000000110;
        weights1[27174] <= 16'b1111111111110111;
        weights1[27175] <= 16'b0000000000001101;
        weights1[27176] <= 16'b0000000000010000;
        weights1[27177] <= 16'b1111111111110110;
        weights1[27178] <= 16'b1111111111111110;
        weights1[27179] <= 16'b1111111111110111;
        weights1[27180] <= 16'b1111111111101100;
        weights1[27181] <= 16'b0000000000000101;
        weights1[27182] <= 16'b1111111111111010;
        weights1[27183] <= 16'b0000000000001000;
        weights1[27184] <= 16'b1111111111111101;
        weights1[27185] <= 16'b0000000000010010;
        weights1[27186] <= 16'b1111111111111110;
        weights1[27187] <= 16'b0000000000000110;
        weights1[27188] <= 16'b1111111111111110;
        weights1[27189] <= 16'b1111111111111100;
        weights1[27190] <= 16'b1111111111110110;
        weights1[27191] <= 16'b1111111111101111;
        weights1[27192] <= 16'b0000000000000001;
        weights1[27193] <= 16'b0000000000010111;
        weights1[27194] <= 16'b1111111111111010;
        weights1[27195] <= 16'b1111111111101011;
        weights1[27196] <= 16'b1111111111111011;
        weights1[27197] <= 16'b1111111111110111;
        weights1[27198] <= 16'b1111111111101101;
        weights1[27199] <= 16'b1111111111110111;
        weights1[27200] <= 16'b1111111111101000;
        weights1[27201] <= 16'b1111111111110001;
        weights1[27202] <= 16'b0000000000000001;
        weights1[27203] <= 16'b0000000000000001;
        weights1[27204] <= 16'b1111111111101110;
        weights1[27205] <= 16'b1111111111110110;
        weights1[27206] <= 16'b1111111111111111;
        weights1[27207] <= 16'b1111111111111011;
        weights1[27208] <= 16'b0000000000000001;
        weights1[27209] <= 16'b1111111111110010;
        weights1[27210] <= 16'b0000000000010100;
        weights1[27211] <= 16'b1111111111111101;
        weights1[27212] <= 16'b1111111111111101;
        weights1[27213] <= 16'b0000000000000011;
        weights1[27214] <= 16'b0000000000001010;
        weights1[27215] <= 16'b0000000000000110;
        weights1[27216] <= 16'b1111111111111011;
        weights1[27217] <= 16'b1111111111111001;
        weights1[27218] <= 16'b1111111111101011;
        weights1[27219] <= 16'b1111111111110101;
        weights1[27220] <= 16'b1111111111111101;
        weights1[27221] <= 16'b1111111111110100;
        weights1[27222] <= 16'b1111111111111010;
        weights1[27223] <= 16'b1111111111111110;
        weights1[27224] <= 16'b1111111111110100;
        weights1[27225] <= 16'b1111111111110110;
        weights1[27226] <= 16'b0000000000010011;
        weights1[27227] <= 16'b0000000000000110;
        weights1[27228] <= 16'b1111111111111111;
        weights1[27229] <= 16'b0000000000000000;
        weights1[27230] <= 16'b0000000000000001;
        weights1[27231] <= 16'b0000000000000111;
        weights1[27232] <= 16'b0000000000010001;
        weights1[27233] <= 16'b0000000000001011;
        weights1[27234] <= 16'b1111111111111000;
        weights1[27235] <= 16'b1111111111111000;
        weights1[27236] <= 16'b1111111111110001;
        weights1[27237] <= 16'b0000000000001001;
        weights1[27238] <= 16'b0000000000001100;
        weights1[27239] <= 16'b0000000000001100;
        weights1[27240] <= 16'b0000000000001100;
        weights1[27241] <= 16'b0000000000000100;
        weights1[27242] <= 16'b0000000000000011;
        weights1[27243] <= 16'b0000000000000101;
        weights1[27244] <= 16'b1111111111111010;
        weights1[27245] <= 16'b1111111111111010;
        weights1[27246] <= 16'b1111111111101110;
        weights1[27247] <= 16'b1111111111100110;
        weights1[27248] <= 16'b1111111111111111;
        weights1[27249] <= 16'b1111111111111001;
        weights1[27250] <= 16'b1111111111100101;
        weights1[27251] <= 16'b0000000000000001;
        weights1[27252] <= 16'b1111111111101101;
        weights1[27253] <= 16'b0000000000010000;
        weights1[27254] <= 16'b0000000000000010;
        weights1[27255] <= 16'b1111111111111100;
        weights1[27256] <= 16'b1111111111111010;
        weights1[27257] <= 16'b0000000000000000;
        weights1[27258] <= 16'b1111111111101101;
        weights1[27259] <= 16'b1111111111111111;
        weights1[27260] <= 16'b1111111111110101;
        weights1[27261] <= 16'b0000000000000100;
        weights1[27262] <= 16'b0000000000000010;
        weights1[27263] <= 16'b0000000000010100;
        weights1[27264] <= 16'b0000000000000000;
        weights1[27265] <= 16'b0000000000000000;
        weights1[27266] <= 16'b1111111111111011;
        weights1[27267] <= 16'b1111111111111110;
        weights1[27268] <= 16'b1111111111111100;
        weights1[27269] <= 16'b1111111111111100;
        weights1[27270] <= 16'b0000000000000011;
        weights1[27271] <= 16'b0000000000000100;
        weights1[27272] <= 16'b0000000000000010;
        weights1[27273] <= 16'b1111111111111000;
        weights1[27274] <= 16'b1111111111111110;
        weights1[27275] <= 16'b1111111111110000;
        weights1[27276] <= 16'b0000000000000000;
        weights1[27277] <= 16'b1111111111110010;
        weights1[27278] <= 16'b0000000000000000;
        weights1[27279] <= 16'b0000000000000101;
        weights1[27280] <= 16'b1111111111111100;
        weights1[27281] <= 16'b0000000000001111;
        weights1[27282] <= 16'b1111111111111110;
        weights1[27283] <= 16'b0000000000000100;
        weights1[27284] <= 16'b0000000000000000;
        weights1[27285] <= 16'b0000000000000111;
        weights1[27286] <= 16'b1111111111110100;
        weights1[27287] <= 16'b1111111111111110;
        weights1[27288] <= 16'b1111111111110100;
        weights1[27289] <= 16'b1111111111110110;
        weights1[27290] <= 16'b0000000000000011;
        weights1[27291] <= 16'b1111111111100001;
        weights1[27292] <= 16'b0000000000100100;
        weights1[27293] <= 16'b0000000000001010;
        weights1[27294] <= 16'b0000000000001011;
        weights1[27295] <= 16'b0000000000000011;
        weights1[27296] <= 16'b1111111111110000;
        weights1[27297] <= 16'b1111111111110111;
        weights1[27298] <= 16'b0000000000000110;
        weights1[27299] <= 16'b0000000000000000;
        weights1[27300] <= 16'b1111111111111011;
        weights1[27301] <= 16'b1111111111111011;
        weights1[27302] <= 16'b0000000000001110;
        weights1[27303] <= 16'b1111111111111001;
        weights1[27304] <= 16'b0000000000000010;
        weights1[27305] <= 16'b0000000000000100;
        weights1[27306] <= 16'b0000000000001000;
        weights1[27307] <= 16'b0000000000001111;
        weights1[27308] <= 16'b1111111111110100;
        weights1[27309] <= 16'b0000000000010001;
        weights1[27310] <= 16'b1111111111111101;
        weights1[27311] <= 16'b1111111111111100;
        weights1[27312] <= 16'b1111111111111000;
        weights1[27313] <= 16'b1111111111101001;
        weights1[27314] <= 16'b0000000000000010;
        weights1[27315] <= 16'b1111111111110000;
        weights1[27316] <= 16'b1111111111111101;
        weights1[27317] <= 16'b0000000000000100;
        weights1[27318] <= 16'b1111111111101010;
        weights1[27319] <= 16'b0000000000001001;
        weights1[27320] <= 16'b0000000000000101;
        weights1[27321] <= 16'b1111111111111111;
        weights1[27322] <= 16'b0000000000000000;
        weights1[27323] <= 16'b0000000000000100;
        weights1[27324] <= 16'b0000000000010001;
        weights1[27325] <= 16'b0000000000010000;
        weights1[27326] <= 16'b0000000000000100;
        weights1[27327] <= 16'b0000000000000001;
        weights1[27328] <= 16'b0000000000000101;
        weights1[27329] <= 16'b1111111111111101;
        weights1[27330] <= 16'b0000000000001000;
        weights1[27331] <= 16'b0000000000000110;
        weights1[27332] <= 16'b1111111111111101;
        weights1[27333] <= 16'b0000000000000101;
        weights1[27334] <= 16'b1111111111111100;
        weights1[27335] <= 16'b0000000000010010;
        weights1[27336] <= 16'b1111111111111000;
        weights1[27337] <= 16'b1111111111110001;
        weights1[27338] <= 16'b1111111111111011;
        weights1[27339] <= 16'b1111111111111010;
        weights1[27340] <= 16'b0000000000000010;
        weights1[27341] <= 16'b0000000000010000;
        weights1[27342] <= 16'b0000000000000110;
        weights1[27343] <= 16'b1111111111111010;
        weights1[27344] <= 16'b1111111111111111;
        weights1[27345] <= 16'b0000000000000000;
        weights1[27346] <= 16'b1111111111100111;
        weights1[27347] <= 16'b1111111111111001;
        weights1[27348] <= 16'b1111111111110111;
        weights1[27349] <= 16'b1111111111110110;
        weights1[27350] <= 16'b0000000000000011;
        weights1[27351] <= 16'b0000000000000000;
        weights1[27352] <= 16'b1111111111111110;
        weights1[27353] <= 16'b0000000000001101;
        weights1[27354] <= 16'b0000000000001101;
        weights1[27355] <= 16'b0000000000000110;
        weights1[27356] <= 16'b0000000000000110;
        weights1[27357] <= 16'b0000000000000000;
        weights1[27358] <= 16'b1111111111111100;
        weights1[27359] <= 16'b1111111111111011;
        weights1[27360] <= 16'b0000000000000100;
        weights1[27361] <= 16'b1111111111111100;
        weights1[27362] <= 16'b0000000000000111;
        weights1[27363] <= 16'b1111111111111111;
        weights1[27364] <= 16'b0000000000000100;
        weights1[27365] <= 16'b0000000000001100;
        weights1[27366] <= 16'b0000000000001000;
        weights1[27367] <= 16'b0000000000000101;
        weights1[27368] <= 16'b0000000000000011;
        weights1[27369] <= 16'b0000000000000010;
        weights1[27370] <= 16'b1111111111101110;
        weights1[27371] <= 16'b0000000000001011;
        weights1[27372] <= 16'b1111111111110101;
        weights1[27373] <= 16'b1111111111111000;
        weights1[27374] <= 16'b0000000000000100;
        weights1[27375] <= 16'b0000000000000001;
        weights1[27376] <= 16'b1111111111101011;
        weights1[27377] <= 16'b1111111111101111;
        weights1[27378] <= 16'b1111111111110101;
        weights1[27379] <= 16'b0000000000000010;
        weights1[27380] <= 16'b1111111111110011;
        weights1[27381] <= 16'b0000000000000011;
        weights1[27382] <= 16'b0000000000001000;
        weights1[27383] <= 16'b0000000000000110;
        weights1[27384] <= 16'b0000000000000100;
        weights1[27385] <= 16'b0000000000000010;
        weights1[27386] <= 16'b0000000000000001;
        weights1[27387] <= 16'b0000000000000100;
        weights1[27388] <= 16'b0000000000000000;
        weights1[27389] <= 16'b0000000000001000;
        weights1[27390] <= 16'b0000000000001001;
        weights1[27391] <= 16'b0000000000001100;
        weights1[27392] <= 16'b0000000000000010;
        weights1[27393] <= 16'b0000000000001011;
        weights1[27394] <= 16'b1111111111111110;
        weights1[27395] <= 16'b1111111111110111;
        weights1[27396] <= 16'b1111111111111011;
        weights1[27397] <= 16'b1111111111110101;
        weights1[27398] <= 16'b1111111111110100;
        weights1[27399] <= 16'b1111111111111001;
        weights1[27400] <= 16'b1111111111111011;
        weights1[27401] <= 16'b1111111111111000;
        weights1[27402] <= 16'b0000000000001001;
        weights1[27403] <= 16'b0000000000000110;
        weights1[27404] <= 16'b0000000000011011;
        weights1[27405] <= 16'b0000000000011011;
        weights1[27406] <= 16'b0000000000010100;
        weights1[27407] <= 16'b0000000000000010;
        weights1[27408] <= 16'b1111111111110100;
        weights1[27409] <= 16'b1111111111111101;
        weights1[27410] <= 16'b1111111111111100;
        weights1[27411] <= 16'b0000000000000001;
        weights1[27412] <= 16'b0000000000000001;
        weights1[27413] <= 16'b0000000000000011;
        weights1[27414] <= 16'b1111111111111011;
        weights1[27415] <= 16'b0000000000000000;
        weights1[27416] <= 16'b1111111111101010;
        weights1[27417] <= 16'b1111111111111001;
        weights1[27418] <= 16'b0000000000010010;
        weights1[27419] <= 16'b0000000000001011;
        weights1[27420] <= 16'b1111111111111111;
        weights1[27421] <= 16'b0000000000000100;
        weights1[27422] <= 16'b0000000000000110;
        weights1[27423] <= 16'b0000000000001001;
        weights1[27424] <= 16'b0000000000000011;
        weights1[27425] <= 16'b0000000000001000;
        weights1[27426] <= 16'b0000000000000101;
        weights1[27427] <= 16'b0000000000001010;
        weights1[27428] <= 16'b0000000000001010;
        weights1[27429] <= 16'b0000000000001100;
        weights1[27430] <= 16'b0000000000000110;
        weights1[27431] <= 16'b0000000000001101;
        weights1[27432] <= 16'b0000000000010001;
        weights1[27433] <= 16'b0000000000001110;
        weights1[27434] <= 16'b0000000000010001;
        weights1[27435] <= 16'b0000000000000101;
        weights1[27436] <= 16'b1111111111111011;
        weights1[27437] <= 16'b1111111111111101;
        weights1[27438] <= 16'b1111111111111101;
        weights1[27439] <= 16'b0000000000000010;
        weights1[27440] <= 16'b0000000000000001;
        weights1[27441] <= 16'b0000000000000001;
        weights1[27442] <= 16'b0000000000000011;
        weights1[27443] <= 16'b0000000000001110;
        weights1[27444] <= 16'b0000000000010111;
        weights1[27445] <= 16'b0000000000010011;
        weights1[27446] <= 16'b0000000000100001;
        weights1[27447] <= 16'b0000000000011000;
        weights1[27448] <= 16'b0000000000011010;
        weights1[27449] <= 16'b0000000000100011;
        weights1[27450] <= 16'b0000000000011101;
        weights1[27451] <= 16'b0000000000000011;
        weights1[27452] <= 16'b0000000000100111;
        weights1[27453] <= 16'b0000000000011000;
        weights1[27454] <= 16'b0000000000010100;
        weights1[27455] <= 16'b0000000000000110;
        weights1[27456] <= 16'b0000000000001111;
        weights1[27457] <= 16'b0000000000010010;
        weights1[27458] <= 16'b0000000000010111;
        weights1[27459] <= 16'b0000000000001111;
        weights1[27460] <= 16'b0000000000000011;
        weights1[27461] <= 16'b0000000000001001;
        weights1[27462] <= 16'b0000000000001111;
        weights1[27463] <= 16'b0000000000001010;
        weights1[27464] <= 16'b0000000000000001;
        weights1[27465] <= 16'b0000000000000011;
        weights1[27466] <= 16'b1111111111111101;
        weights1[27467] <= 16'b1111111111111111;
        weights1[27468] <= 16'b0000000000000000;
        weights1[27469] <= 16'b0000000000000011;
        weights1[27470] <= 16'b0000000000010001;
        weights1[27471] <= 16'b0000000000011000;
        weights1[27472] <= 16'b0000000000011011;
        weights1[27473] <= 16'b0000000000010000;
        weights1[27474] <= 16'b0000000000011010;
        weights1[27475] <= 16'b0000000000010000;
        weights1[27476] <= 16'b1111111111111001;
        weights1[27477] <= 16'b0000000000001011;
        weights1[27478] <= 16'b1111111111111111;
        weights1[27479] <= 16'b1111111111101110;
        weights1[27480] <= 16'b0000000000000110;
        weights1[27481] <= 16'b0000000000001011;
        weights1[27482] <= 16'b1111111111111010;
        weights1[27483] <= 16'b0000000000001000;
        weights1[27484] <= 16'b0000000000001101;
        weights1[27485] <= 16'b0000000000000000;
        weights1[27486] <= 16'b1111111111111111;
        weights1[27487] <= 16'b0000000000001100;
        weights1[27488] <= 16'b1111111111110111;
        weights1[27489] <= 16'b0000000000001111;
        weights1[27490] <= 16'b0000000000001011;
        weights1[27491] <= 16'b1111111111111111;
        weights1[27492] <= 16'b1111111111111000;
        weights1[27493] <= 16'b0000000000001001;
        weights1[27494] <= 16'b0000000000000111;
        weights1[27495] <= 16'b0000000000000100;
        weights1[27496] <= 16'b1111111111111101;
        weights1[27497] <= 16'b0000000000001001;
        weights1[27498] <= 16'b0000000000001111;
        weights1[27499] <= 16'b0000000000001010;
        weights1[27500] <= 16'b0000000000001000;
        weights1[27501] <= 16'b0000000000010011;
        weights1[27502] <= 16'b0000000000011010;
        weights1[27503] <= 16'b0000000000000101;
        weights1[27504] <= 16'b1111111111111100;
        weights1[27505] <= 16'b0000000000001110;
        weights1[27506] <= 16'b0000000000000100;
        weights1[27507] <= 16'b1111111111111011;
        weights1[27508] <= 16'b1111111111110011;
        weights1[27509] <= 16'b0000000000000111;
        weights1[27510] <= 16'b1111111111111010;
        weights1[27511] <= 16'b1111111111110110;
        weights1[27512] <= 16'b1111111111111001;
        weights1[27513] <= 16'b1111111111101110;
        weights1[27514] <= 16'b0000000000010001;
        weights1[27515] <= 16'b0000000000000001;
        weights1[27516] <= 16'b0000000000000100;
        weights1[27517] <= 16'b0000000000001110;
        weights1[27518] <= 16'b1111111111111101;
        weights1[27519] <= 16'b1111111111101101;
        weights1[27520] <= 16'b0000000000000011;
        weights1[27521] <= 16'b1111111111111000;
        weights1[27522] <= 16'b1111111111111001;
        weights1[27523] <= 16'b0000000000001000;
        weights1[27524] <= 16'b1111111111111011;
        weights1[27525] <= 16'b0000000000000111;
        weights1[27526] <= 16'b0000000000000011;
        weights1[27527] <= 16'b0000000000000011;
        weights1[27528] <= 16'b0000000000011101;
        weights1[27529] <= 16'b0000000000000111;
        weights1[27530] <= 16'b0000000000000110;
        weights1[27531] <= 16'b0000000000001110;
        weights1[27532] <= 16'b1111111111110101;
        weights1[27533] <= 16'b1111111111111011;
        weights1[27534] <= 16'b1111111111111001;
        weights1[27535] <= 16'b1111111111101010;
        weights1[27536] <= 16'b1111111111110100;
        weights1[27537] <= 16'b1111111111101110;
        weights1[27538] <= 16'b1111111111111000;
        weights1[27539] <= 16'b1111111111110011;
        weights1[27540] <= 16'b1111111111111111;
        weights1[27541] <= 16'b0000000000000001;
        weights1[27542] <= 16'b1111111111110100;
        weights1[27543] <= 16'b0000000000000100;
        weights1[27544] <= 16'b1111111111111010;
        weights1[27545] <= 16'b1111111111111000;
        weights1[27546] <= 16'b1111111111111111;
        weights1[27547] <= 16'b0000000000000110;
        weights1[27548] <= 16'b1111111111111010;
        weights1[27549] <= 16'b0000000000001000;
        weights1[27550] <= 16'b1111111111111110;
        weights1[27551] <= 16'b1111111111111110;
        weights1[27552] <= 16'b1111111111111011;
        weights1[27553] <= 16'b0000000000000000;
        weights1[27554] <= 16'b1111111111111010;
        weights1[27555] <= 16'b1111111111111011;
        weights1[27556] <= 16'b0000000000000100;
        weights1[27557] <= 16'b0000000000000110;
        weights1[27558] <= 16'b1111111111111101;
        weights1[27559] <= 16'b1111111111110001;
        weights1[27560] <= 16'b1111111111110111;
        weights1[27561] <= 16'b0000000000001000;
        weights1[27562] <= 16'b1111111111110011;
        weights1[27563] <= 16'b1111111111110111;
        weights1[27564] <= 16'b1111111111111111;
        weights1[27565] <= 16'b1111111111111001;
        weights1[27566] <= 16'b1111111111110110;
        weights1[27567] <= 16'b1111111111110110;
        weights1[27568] <= 16'b1111111111110100;
        weights1[27569] <= 16'b0000000000000001;
        weights1[27570] <= 16'b1111111111111110;
        weights1[27571] <= 16'b1111111111110010;
        weights1[27572] <= 16'b1111111111111001;
        weights1[27573] <= 16'b1111111111111111;
        weights1[27574] <= 16'b1111111111101111;
        weights1[27575] <= 16'b1111111111111010;
        weights1[27576] <= 16'b1111111111111000;
        weights1[27577] <= 16'b0000000000000100;
        weights1[27578] <= 16'b0000000000000110;
        weights1[27579] <= 16'b1111111111110100;
        weights1[27580] <= 16'b1111111111110111;
        weights1[27581] <= 16'b1111111111111100;
        weights1[27582] <= 16'b1111111111111011;
        weights1[27583] <= 16'b1111111111110110;
        weights1[27584] <= 16'b1111111111111110;
        weights1[27585] <= 16'b1111111111111111;
        weights1[27586] <= 16'b0000000000001100;
        weights1[27587] <= 16'b1111111111110011;
        weights1[27588] <= 16'b1111111111110110;
        weights1[27589] <= 16'b1111111111111101;
        weights1[27590] <= 16'b1111111111111111;
        weights1[27591] <= 16'b1111111111110111;
        weights1[27592] <= 16'b1111111111111100;
        weights1[27593] <= 16'b1111111111110111;
        weights1[27594] <= 16'b1111111111110001;
        weights1[27595] <= 16'b1111111111111000;
        weights1[27596] <= 16'b1111111111110010;
        weights1[27597] <= 16'b1111111111110001;
        weights1[27598] <= 16'b1111111111100100;
        weights1[27599] <= 16'b1111111111110111;
        weights1[27600] <= 16'b1111111111111100;
        weights1[27601] <= 16'b1111111111100100;
        weights1[27602] <= 16'b1111111111111001;
        weights1[27603] <= 16'b1111111111111111;
        weights1[27604] <= 16'b0000000000000101;
        weights1[27605] <= 16'b0000000000001010;
        weights1[27606] <= 16'b1111111111111010;
        weights1[27607] <= 16'b1111111111111000;
        weights1[27608] <= 16'b1111111111111000;
        weights1[27609] <= 16'b0000000000000100;
        weights1[27610] <= 16'b1111111111111001;
        weights1[27611] <= 16'b1111111111110001;
        weights1[27612] <= 16'b0000000000001001;
        weights1[27613] <= 16'b1111111111110111;
        weights1[27614] <= 16'b1111111111110110;
        weights1[27615] <= 16'b1111111111111110;
        weights1[27616] <= 16'b0000000000000001;
        weights1[27617] <= 16'b1111111111111011;
        weights1[27618] <= 16'b1111111111111111;
        weights1[27619] <= 16'b1111111111110000;
        weights1[27620] <= 16'b1111111111111111;
        weights1[27621] <= 16'b1111111111111110;
        weights1[27622] <= 16'b1111111111111111;
        weights1[27623] <= 16'b1111111111111100;
        weights1[27624] <= 16'b1111111111110011;
        weights1[27625] <= 16'b1111111111111011;
        weights1[27626] <= 16'b0000000000000101;
        weights1[27627] <= 16'b1111111111101101;
        weights1[27628] <= 16'b1111111111110110;
        weights1[27629] <= 16'b0000000000000110;
        weights1[27630] <= 16'b0000000000001000;
        weights1[27631] <= 16'b1111111111111111;
        weights1[27632] <= 16'b1111111111100101;
        weights1[27633] <= 16'b1111111111110010;
        weights1[27634] <= 16'b1111111111111101;
        weights1[27635] <= 16'b1111111111110111;
        weights1[27636] <= 16'b1111111111111101;
        weights1[27637] <= 16'b0000000000000101;
        weights1[27638] <= 16'b1111111111111100;
        weights1[27639] <= 16'b0000000000000000;
        weights1[27640] <= 16'b0000000000000011;
        weights1[27641] <= 16'b0000000000000101;
        weights1[27642] <= 16'b0000000000000100;
        weights1[27643] <= 16'b0000000000000011;
        weights1[27644] <= 16'b1111111111111011;
        weights1[27645] <= 16'b0000000000000010;
        weights1[27646] <= 16'b1111111111110110;
        weights1[27647] <= 16'b0000000000000010;
        weights1[27648] <= 16'b1111111111111010;
        weights1[27649] <= 16'b1111111111110110;
        weights1[27650] <= 16'b0000000000001010;
        weights1[27651] <= 16'b1111111111111111;
        weights1[27652] <= 16'b0000000000000010;
        weights1[27653] <= 16'b1111111111111111;
        weights1[27654] <= 16'b0000000000000011;
        weights1[27655] <= 16'b0000000000000101;
        weights1[27656] <= 16'b0000000000001110;
        weights1[27657] <= 16'b1111111111110101;
        weights1[27658] <= 16'b1111111111110000;
        weights1[27659] <= 16'b1111111111111010;
        weights1[27660] <= 16'b1111111111111010;
        weights1[27661] <= 16'b0000000000000001;
        weights1[27662] <= 16'b1111111111111011;
        weights1[27663] <= 16'b1111111111101100;
        weights1[27664] <= 16'b1111111111110010;
        weights1[27665] <= 16'b0000000000000000;
        weights1[27666] <= 16'b1111111111110101;
        weights1[27667] <= 16'b1111111111110101;
        weights1[27668] <= 16'b0000000000000100;
        weights1[27669] <= 16'b1111111111111000;
        weights1[27670] <= 16'b1111111111110101;
        weights1[27671] <= 16'b1111111111111001;
        weights1[27672] <= 16'b1111111111111001;
        weights1[27673] <= 16'b0000000000001101;
        weights1[27674] <= 16'b1111111111111000;
        weights1[27675] <= 16'b0000000000001010;
        weights1[27676] <= 16'b0000000000000001;
        weights1[27677] <= 16'b0000000000000011;
        weights1[27678] <= 16'b0000000000000000;
        weights1[27679] <= 16'b0000000000000111;
        weights1[27680] <= 16'b1111111111111110;
        weights1[27681] <= 16'b0000000000000010;
        weights1[27682] <= 16'b0000000000001001;
        weights1[27683] <= 16'b1111111111111101;
        weights1[27684] <= 16'b1111111111110010;
        weights1[27685] <= 16'b1111111111110001;
        weights1[27686] <= 16'b1111111111101101;
        weights1[27687] <= 16'b0000000000000100;
        weights1[27688] <= 16'b0000000000000001;
        weights1[27689] <= 16'b0000000000001111;
        weights1[27690] <= 16'b1111111111110011;
        weights1[27691] <= 16'b1111111111110111;
        weights1[27692] <= 16'b1111111111111001;
        weights1[27693] <= 16'b1111111111110100;
        weights1[27694] <= 16'b0000000000000000;
        weights1[27695] <= 16'b1111111111110110;
        weights1[27696] <= 16'b1111111111111111;
        weights1[27697] <= 16'b0000000000001000;
        weights1[27698] <= 16'b1111111111101100;
        weights1[27699] <= 16'b1111111111111101;
        weights1[27700] <= 16'b1111111111111111;
        weights1[27701] <= 16'b0000000000001001;
        weights1[27702] <= 16'b0000000000010000;
        weights1[27703] <= 16'b1111111111111010;
        weights1[27704] <= 16'b0000000000010000;
        weights1[27705] <= 16'b0000000000001001;
        weights1[27706] <= 16'b0000000000001111;
        weights1[27707] <= 16'b0000000000001000;
        weights1[27708] <= 16'b1111111111111111;
        weights1[27709] <= 16'b1111111111110001;
        weights1[27710] <= 16'b0000000000000101;
        weights1[27711] <= 16'b0000000000000011;
        weights1[27712] <= 16'b0000000000001100;
        weights1[27713] <= 16'b1111111111111101;
        weights1[27714] <= 16'b0000000000010010;
        weights1[27715] <= 16'b1111111111111011;
        weights1[27716] <= 16'b0000000000001001;
        weights1[27717] <= 16'b0000000000000000;
        weights1[27718] <= 16'b1111111111101011;
        weights1[27719] <= 16'b0000000000000001;
        weights1[27720] <= 16'b1111111111111011;
        weights1[27721] <= 16'b0000000000000000;
        weights1[27722] <= 16'b0000000000001000;
        weights1[27723] <= 16'b1111111111111001;
        weights1[27724] <= 16'b1111111111111101;
        weights1[27725] <= 16'b1111111111111110;
        weights1[27726] <= 16'b0000000000000011;
        weights1[27727] <= 16'b0000000000001100;
        weights1[27728] <= 16'b0000000000000010;
        weights1[27729] <= 16'b0000000000000011;
        weights1[27730] <= 16'b0000000000010011;
        weights1[27731] <= 16'b0000000000001011;
        weights1[27732] <= 16'b0000000000001010;
        weights1[27733] <= 16'b1111111111111100;
        weights1[27734] <= 16'b1111111111111100;
        weights1[27735] <= 16'b1111111111111110;
        weights1[27736] <= 16'b0000000000000110;
        weights1[27737] <= 16'b0000000000001000;
        weights1[27738] <= 16'b1111111111111110;
        weights1[27739] <= 16'b0000000000001010;
        weights1[27740] <= 16'b1111111111111101;
        weights1[27741] <= 16'b0000000000000001;
        weights1[27742] <= 16'b0000000000010000;
        weights1[27743] <= 16'b0000000000001001;
        weights1[27744] <= 16'b1111111111101111;
        weights1[27745] <= 16'b0000000000001101;
        weights1[27746] <= 16'b0000000000000010;
        weights1[27747] <= 16'b0000000000001101;
        weights1[27748] <= 16'b1111111111111101;
        weights1[27749] <= 16'b0000000000001001;
        weights1[27750] <= 16'b0000000000001111;
        weights1[27751] <= 16'b0000000000011110;
        weights1[27752] <= 16'b0000000000001001;
        weights1[27753] <= 16'b1111111111111000;
        weights1[27754] <= 16'b1111111111111101;
        weights1[27755] <= 16'b1111111111111110;
        weights1[27756] <= 16'b0000000000001011;
        weights1[27757] <= 16'b0000000000001011;
        weights1[27758] <= 16'b0000000000001001;
        weights1[27759] <= 16'b1111111111111011;
        weights1[27760] <= 16'b0000000000000001;
        weights1[27761] <= 16'b1111111111111001;
        weights1[27762] <= 16'b0000000000001100;
        weights1[27763] <= 16'b0000000000000010;
        weights1[27764] <= 16'b0000000000000001;
        weights1[27765] <= 16'b0000000000000101;
        weights1[27766] <= 16'b0000000000001011;
        weights1[27767] <= 16'b0000000000001000;
        weights1[27768] <= 16'b0000000000000111;
        weights1[27769] <= 16'b0000000000011010;
        weights1[27770] <= 16'b0000000000000000;
        weights1[27771] <= 16'b0000000000011000;
        weights1[27772] <= 16'b0000000000001100;
        weights1[27773] <= 16'b0000000000010010;
        weights1[27774] <= 16'b0000000000000010;
        weights1[27775] <= 16'b0000000000001001;
        weights1[27776] <= 16'b0000000000000111;
        weights1[27777] <= 16'b0000000000001111;
        weights1[27778] <= 16'b0000000000011111;
        weights1[27779] <= 16'b1111111111111110;
        weights1[27780] <= 16'b0000000000000100;
        weights1[27781] <= 16'b0000000000010100;
        weights1[27782] <= 16'b0000000000001011;
        weights1[27783] <= 16'b0000000000000010;
        weights1[27784] <= 16'b1111111111110000;
        weights1[27785] <= 16'b0000000000000100;
        weights1[27786] <= 16'b1111111111111011;
        weights1[27787] <= 16'b0000000000010101;
        weights1[27788] <= 16'b0000000000011000;
        weights1[27789] <= 16'b0000000000000110;
        weights1[27790] <= 16'b0000000000000010;
        weights1[27791] <= 16'b0000000000001011;
        weights1[27792] <= 16'b1111111111111110;
        weights1[27793] <= 16'b0000000000000101;
        weights1[27794] <= 16'b0000000000000010;
        weights1[27795] <= 16'b1111111111111111;
        weights1[27796] <= 16'b0000000000000111;
        weights1[27797] <= 16'b0000000000000010;
        weights1[27798] <= 16'b0000000000001000;
        weights1[27799] <= 16'b0000000000011010;
        weights1[27800] <= 16'b1111111111111111;
        weights1[27801] <= 16'b0000000000001001;
        weights1[27802] <= 16'b0000000000010000;
        weights1[27803] <= 16'b0000000000010101;
        weights1[27804] <= 16'b0000000000001101;
        weights1[27805] <= 16'b0000000000001110;
        weights1[27806] <= 16'b0000000000010000;
        weights1[27807] <= 16'b0000000000010010;
        weights1[27808] <= 16'b0000000000000111;
        weights1[27809] <= 16'b0000000000001100;
        weights1[27810] <= 16'b1111111111111001;
        weights1[27811] <= 16'b0000000000000001;
        weights1[27812] <= 16'b0000000000011010;
        weights1[27813] <= 16'b1111111111111100;
        weights1[27814] <= 16'b0000000000000101;
        weights1[27815] <= 16'b1111111111111101;
        weights1[27816] <= 16'b0000000000000010;
        weights1[27817] <= 16'b0000000000000111;
        weights1[27818] <= 16'b0000000000001000;
        weights1[27819] <= 16'b0000000000001000;
        weights1[27820] <= 16'b0000000000000101;
        weights1[27821] <= 16'b0000000000001101;
        weights1[27822] <= 16'b0000000000001100;
        weights1[27823] <= 16'b0000000000010111;
        weights1[27824] <= 16'b1111111111110110;
        weights1[27825] <= 16'b0000000000010010;
        weights1[27826] <= 16'b0000000000011000;
        weights1[27827] <= 16'b0000000000001011;
        weights1[27828] <= 16'b0000000000010000;
        weights1[27829] <= 16'b0000000000001011;
        weights1[27830] <= 16'b0000000000001010;
        weights1[27831] <= 16'b0000000000001011;
        weights1[27832] <= 16'b0000000000001010;
        weights1[27833] <= 16'b0000000000001000;
        weights1[27834] <= 16'b0000000000001100;
        weights1[27835] <= 16'b0000000000011111;
        weights1[27836] <= 16'b0000000000010000;
        weights1[27837] <= 16'b0000000000011011;
        weights1[27838] <= 16'b0000000000010011;
        weights1[27839] <= 16'b0000000000001110;
        weights1[27840] <= 16'b0000000000010000;
        weights1[27841] <= 16'b0000000000001010;
        weights1[27842] <= 16'b0000000000001010;
        weights1[27843] <= 16'b1111111111111010;
        weights1[27844] <= 16'b0000000000000111;
        weights1[27845] <= 16'b0000000000001100;
        weights1[27846] <= 16'b0000000000001110;
        weights1[27847] <= 16'b1111111111111011;
        weights1[27848] <= 16'b0000000000001110;
        weights1[27849] <= 16'b1111111111111111;
        weights1[27850] <= 16'b0000000000000110;
        weights1[27851] <= 16'b0000000000010010;
        weights1[27852] <= 16'b0000000000000110;
        weights1[27853] <= 16'b0000000000000011;
        weights1[27854] <= 16'b0000000000010011;
        weights1[27855] <= 16'b0000000000100001;
        weights1[27856] <= 16'b0000000000010000;
        weights1[27857] <= 16'b0000000000001010;
        weights1[27858] <= 16'b1111111111111100;
        weights1[27859] <= 16'b0000000000000011;
        weights1[27860] <= 16'b0000000000000000;
        weights1[27861] <= 16'b0000000000001110;
        weights1[27862] <= 16'b0000000000001101;
        weights1[27863] <= 16'b0000000000010010;
        weights1[27864] <= 16'b0000000000001011;
        weights1[27865] <= 16'b0000000000000111;
        weights1[27866] <= 16'b1111111111101011;
        weights1[27867] <= 16'b0000000000010101;
        weights1[27868] <= 16'b0000000000000100;
        weights1[27869] <= 16'b0000000000000111;
        weights1[27870] <= 16'b0000000000010000;
        weights1[27871] <= 16'b0000000000000000;
        weights1[27872] <= 16'b0000000000000111;
        weights1[27873] <= 16'b0000000000011100;
        weights1[27874] <= 16'b1111111111111110;
        weights1[27875] <= 16'b0000000000001011;
        weights1[27876] <= 16'b0000000000010100;
        weights1[27877] <= 16'b0000000000010000;
        weights1[27878] <= 16'b0000000000100000;
        weights1[27879] <= 16'b0000000000001110;
        weights1[27880] <= 16'b0000000000011101;
        weights1[27881] <= 16'b0000000000000111;
        weights1[27882] <= 16'b0000000000001110;
        weights1[27883] <= 16'b0000000000001101;
        weights1[27884] <= 16'b0000000000001101;
        weights1[27885] <= 16'b0000000000000110;
        weights1[27886] <= 16'b1111111111110001;
        weights1[27887] <= 16'b0000000000000010;
        weights1[27888] <= 16'b0000000000000011;
        weights1[27889] <= 16'b1111111111111101;
        weights1[27890] <= 16'b1111111111111001;
        weights1[27891] <= 16'b0000000000000110;
        weights1[27892] <= 16'b0000000000010111;
        weights1[27893] <= 16'b0000000000011001;
        weights1[27894] <= 16'b0000000000001111;
        weights1[27895] <= 16'b0000000000011000;
        weights1[27896] <= 16'b0000000000001110;
        weights1[27897] <= 16'b0000000000001100;
        weights1[27898] <= 16'b0000000000000111;
        weights1[27899] <= 16'b0000000000010000;
        weights1[27900] <= 16'b0000000000010110;
        weights1[27901] <= 16'b0000000000001101;
        weights1[27902] <= 16'b0000000000001110;
        weights1[27903] <= 16'b0000000000010101;
        weights1[27904] <= 16'b0000000000010111;
        weights1[27905] <= 16'b0000000000010101;
        weights1[27906] <= 16'b0000000000000000;
        weights1[27907] <= 16'b0000000000010111;
        weights1[27908] <= 16'b0000000000010011;
        weights1[27909] <= 16'b0000000000010110;
        weights1[27910] <= 16'b1111111111111110;
        weights1[27911] <= 16'b0000000000001000;
        weights1[27912] <= 16'b0000000000000101;
        weights1[27913] <= 16'b0000000000001001;
        weights1[27914] <= 16'b1111111111101101;
        weights1[27915] <= 16'b1111111111101101;
        weights1[27916] <= 16'b0000000000000001;
        weights1[27917] <= 16'b1111111111111100;
        weights1[27918] <= 16'b1111111111111001;
        weights1[27919] <= 16'b0000000000000001;
        weights1[27920] <= 16'b0000000000000100;
        weights1[27921] <= 16'b1111111111101010;
        weights1[27922] <= 16'b0000000000010101;
        weights1[27923] <= 16'b0000000000001110;
        weights1[27924] <= 16'b1111111111111101;
        weights1[27925] <= 16'b0000000000000110;
        weights1[27926] <= 16'b0000000000000000;
        weights1[27927] <= 16'b0000000000000000;
        weights1[27928] <= 16'b0000000000001100;
        weights1[27929] <= 16'b1111111111111111;
        weights1[27930] <= 16'b0000000000000110;
        weights1[27931] <= 16'b0000000000000001;
        weights1[27932] <= 16'b0000000000011010;
        weights1[27933] <= 16'b0000000000001010;
        weights1[27934] <= 16'b0000000000001011;
        weights1[27935] <= 16'b0000000000010110;
        weights1[27936] <= 16'b0000000000010110;
        weights1[27937] <= 16'b0000000000010111;
        weights1[27938] <= 16'b0000000000010001;
        weights1[27939] <= 16'b0000000000001000;
        weights1[27940] <= 16'b1111111111101100;
        weights1[27941] <= 16'b1111111111100111;
        weights1[27942] <= 16'b1111111111101000;
        weights1[27943] <= 16'b1111111111011000;
        weights1[27944] <= 16'b1111111111111101;
        weights1[27945] <= 16'b1111111111101111;
        weights1[27946] <= 16'b1111111111101010;
        weights1[27947] <= 16'b0000000000000001;
        weights1[27948] <= 16'b0000000000000011;
        weights1[27949] <= 16'b1111111111111001;
        weights1[27950] <= 16'b1111111111110011;
        weights1[27951] <= 16'b1111111111111010;
        weights1[27952] <= 16'b0000000000011010;
        weights1[27953] <= 16'b1111111111111111;
        weights1[27954] <= 16'b0000000000001011;
        weights1[27955] <= 16'b0000000000000101;
        weights1[27956] <= 16'b1111111111111000;
        weights1[27957] <= 16'b0000000000001011;
        weights1[27958] <= 16'b1111111111111001;
        weights1[27959] <= 16'b0000000000000100;
        weights1[27960] <= 16'b1111111111110111;
        weights1[27961] <= 16'b0000000000010000;
        weights1[27962] <= 16'b0000000000100001;
        weights1[27963] <= 16'b0000000000011010;
        weights1[27964] <= 16'b0000000000001111;
        weights1[27965] <= 16'b0000000000001101;
        weights1[27966] <= 16'b1111111111101001;
        weights1[27967] <= 16'b1111111111101100;
        weights1[27968] <= 16'b1111111111100010;
        weights1[27969] <= 16'b1111111111001100;
        weights1[27970] <= 16'b1111111110111110;
        weights1[27971] <= 16'b1111111111001011;
        weights1[27972] <= 16'b1111111111111000;
        weights1[27973] <= 16'b1111111111101010;
        weights1[27974] <= 16'b1111111111101011;
        weights1[27975] <= 16'b1111111111110111;
        weights1[27976] <= 16'b1111111111101001;
        weights1[27977] <= 16'b1111111111111011;
        weights1[27978] <= 16'b1111111111101010;
        weights1[27979] <= 16'b1111111111101100;
        weights1[27980] <= 16'b1111111111110100;
        weights1[27981] <= 16'b1111111111100001;
        weights1[27982] <= 16'b1111111111011011;
        weights1[27983] <= 16'b1111111111110001;
        weights1[27984] <= 16'b1111111111110101;
        weights1[27985] <= 16'b1111111111111100;
        weights1[27986] <= 16'b1111111111111101;
        weights1[27987] <= 16'b0000000000000101;
        weights1[27988] <= 16'b1111111111110001;
        weights1[27989] <= 16'b1111111111101001;
        weights1[27990] <= 16'b1111111111101101;
        weights1[27991] <= 16'b1111111111101101;
        weights1[27992] <= 16'b1111111111011100;
        weights1[27993] <= 16'b1111111111001010;
        weights1[27994] <= 16'b1111111110111111;
        weights1[27995] <= 16'b1111111110101110;
        weights1[27996] <= 16'b1111111110111010;
        weights1[27997] <= 16'b1111111110111101;
        weights1[27998] <= 16'b1111111110111101;
        weights1[27999] <= 16'b1111111111001110;
        weights1[28000] <= 16'b1111111111110010;
        weights1[28001] <= 16'b1111111111100110;
        weights1[28002] <= 16'b1111111111100101;
        weights1[28003] <= 16'b1111111111010101;
        weights1[28004] <= 16'b1111111111010011;
        weights1[28005] <= 16'b1111111111100000;
        weights1[28006] <= 16'b1111111111010011;
        weights1[28007] <= 16'b1111111111000110;
        weights1[28008] <= 16'b1111111111100001;
        weights1[28009] <= 16'b1111111111010010;
        weights1[28010] <= 16'b1111111111001111;
        weights1[28011] <= 16'b1111111111011100;
        weights1[28012] <= 16'b1111111111011111;
        weights1[28013] <= 16'b1111111111001001;
        weights1[28014] <= 16'b1111111111010011;
        weights1[28015] <= 16'b1111111111001010;
        weights1[28016] <= 16'b1111111110111000;
        weights1[28017] <= 16'b1111111110011100;
        weights1[28018] <= 16'b1111111101111011;
        weights1[28019] <= 16'b1111111101111111;
        weights1[28020] <= 16'b1111111101101010;
        weights1[28021] <= 16'b1111111101011100;
        weights1[28022] <= 16'b1111111110010000;
        weights1[28023] <= 16'b1111111110100010;
        weights1[28024] <= 16'b1111111110110000;
        weights1[28025] <= 16'b1111111110100110;
        weights1[28026] <= 16'b1111111111001101;
        weights1[28027] <= 16'b1111111111010001;
        weights1[28028] <= 16'b1111111111110111;
        weights1[28029] <= 16'b1111111111100100;
        weights1[28030] <= 16'b1111111111011100;
        weights1[28031] <= 16'b1111111111010100;
        weights1[28032] <= 16'b1111111111000010;
        weights1[28033] <= 16'b1111111110110011;
        weights1[28034] <= 16'b1111111110100011;
        weights1[28035] <= 16'b1111111110011111;
        weights1[28036] <= 16'b1111111110011100;
        weights1[28037] <= 16'b1111111101111011;
        weights1[28038] <= 16'b1111111110001001;
        weights1[28039] <= 16'b1111111101110011;
        weights1[28040] <= 16'b1111111101110001;
        weights1[28041] <= 16'b1111111101101111;
        weights1[28042] <= 16'b1111111101100111;
        weights1[28043] <= 16'b1111111101100001;
        weights1[28044] <= 16'b1111111101100011;
        weights1[28045] <= 16'b1111111101011111;
        weights1[28046] <= 16'b1111111110000000;
        weights1[28047] <= 16'b1111111101111100;
        weights1[28048] <= 16'b1111111110010100;
        weights1[28049] <= 16'b1111111110101000;
        weights1[28050] <= 16'b1111111110101100;
        weights1[28051] <= 16'b1111111111000000;
        weights1[28052] <= 16'b1111111111010110;
        weights1[28053] <= 16'b1111111111010011;
        weights1[28054] <= 16'b1111111111011011;
        weights1[28055] <= 16'b1111111111100110;
        weights1[28056] <= 16'b1111111111110110;
        weights1[28057] <= 16'b1111111111101111;
        weights1[28058] <= 16'b1111111111100101;
        weights1[28059] <= 16'b1111111111100000;
        weights1[28060] <= 16'b1111111111011011;
        weights1[28061] <= 16'b1111111111011100;
        weights1[28062] <= 16'b1111111111001010;
        weights1[28063] <= 16'b1111111111000011;
        weights1[28064] <= 16'b1111111111000000;
        weights1[28065] <= 16'b1111111110111000;
        weights1[28066] <= 16'b1111111111000000;
        weights1[28067] <= 16'b1111111110100111;
        weights1[28068] <= 16'b1111111110111011;
        weights1[28069] <= 16'b1111111110100011;
        weights1[28070] <= 16'b1111111110101000;
        weights1[28071] <= 16'b1111111110011100;
        weights1[28072] <= 16'b1111111110101010;
        weights1[28073] <= 16'b1111111110100101;
        weights1[28074] <= 16'b1111111110110001;
        weights1[28075] <= 16'b1111111110101010;
        weights1[28076] <= 16'b1111111111000010;
        weights1[28077] <= 16'b1111111111000010;
        weights1[28078] <= 16'b1111111111010011;
        weights1[28079] <= 16'b1111111111010000;
        weights1[28080] <= 16'b1111111111100100;
        weights1[28081] <= 16'b1111111111101100;
        weights1[28082] <= 16'b1111111111101111;
        weights1[28083] <= 16'b1111111111101010;
        weights1[28084] <= 16'b0000000000000000;
        weights1[28085] <= 16'b1111111111111001;
        weights1[28086] <= 16'b1111111111111001;
        weights1[28087] <= 16'b1111111111110101;
        weights1[28088] <= 16'b1111111111110001;
        weights1[28089] <= 16'b1111111111101111;
        weights1[28090] <= 16'b1111111111101010;
        weights1[28091] <= 16'b1111111111100101;
        weights1[28092] <= 16'b1111111111100110;
        weights1[28093] <= 16'b1111111111010101;
        weights1[28094] <= 16'b1111111111100101;
        weights1[28095] <= 16'b1111111111010000;
        weights1[28096] <= 16'b1111111111010101;
        weights1[28097] <= 16'b1111111111001101;
        weights1[28098] <= 16'b1111111111001001;
        weights1[28099] <= 16'b1111111110111010;
        weights1[28100] <= 16'b1111111111001010;
        weights1[28101] <= 16'b1111111111000111;
        weights1[28102] <= 16'b1111111111001011;
        weights1[28103] <= 16'b1111111110111011;
        weights1[28104] <= 16'b1111111111001111;
        weights1[28105] <= 16'b1111111111010111;
        weights1[28106] <= 16'b1111111111011010;
        weights1[28107] <= 16'b1111111111101110;
        weights1[28108] <= 16'b1111111111101100;
        weights1[28109] <= 16'b1111111111110010;
        weights1[28110] <= 16'b1111111111110111;
        weights1[28111] <= 16'b1111111111110100;
        weights1[28112] <= 16'b0000000000000011;
        weights1[28113] <= 16'b0000000000000000;
        weights1[28114] <= 16'b1111111111111010;
        weights1[28115] <= 16'b1111111111111011;
        weights1[28116] <= 16'b1111111111111110;
        weights1[28117] <= 16'b0000000000000100;
        weights1[28118] <= 16'b0000000000000001;
        weights1[28119] <= 16'b1111111111110100;
        weights1[28120] <= 16'b1111111111111111;
        weights1[28121] <= 16'b1111111111110110;
        weights1[28122] <= 16'b1111111111010001;
        weights1[28123] <= 16'b1111111111100001;
        weights1[28124] <= 16'b1111111111101000;
        weights1[28125] <= 16'b1111111111001111;
        weights1[28126] <= 16'b1111111111011100;
        weights1[28127] <= 16'b1111111111101010;
        weights1[28128] <= 16'b1111111111100000;
        weights1[28129] <= 16'b1111111111011101;
        weights1[28130] <= 16'b1111111111100010;
        weights1[28131] <= 16'b1111111111011000;
        weights1[28132] <= 16'b1111111111010110;
        weights1[28133] <= 16'b1111111111010110;
        weights1[28134] <= 16'b1111111111101111;
        weights1[28135] <= 16'b1111111111110000;
        weights1[28136] <= 16'b1111111111111001;
        weights1[28137] <= 16'b1111111111110101;
        weights1[28138] <= 16'b1111111111111001;
        weights1[28139] <= 16'b1111111111111011;
        weights1[28140] <= 16'b0000000000000011;
        weights1[28141] <= 16'b1111111111111110;
        weights1[28142] <= 16'b1111111111111011;
        weights1[28143] <= 16'b0000000000000001;
        weights1[28144] <= 16'b1111111111111110;
        weights1[28145] <= 16'b0000000000000011;
        weights1[28146] <= 16'b0000000000000010;
        weights1[28147] <= 16'b0000000000000000;
        weights1[28148] <= 16'b1111111111111011;
        weights1[28149] <= 16'b1111111111101110;
        weights1[28150] <= 16'b1111111111101011;
        weights1[28151] <= 16'b1111111111110100;
        weights1[28152] <= 16'b1111111111101101;
        weights1[28153] <= 16'b1111111111101000;
        weights1[28154] <= 16'b1111111111100111;
        weights1[28155] <= 16'b1111111111110111;
        weights1[28156] <= 16'b1111111111100111;
        weights1[28157] <= 16'b1111111111100110;
        weights1[28158] <= 16'b1111111111110110;
        weights1[28159] <= 16'b1111111111011101;
        weights1[28160] <= 16'b1111111111100101;
        weights1[28161] <= 16'b1111111111111000;
        weights1[28162] <= 16'b1111111111111001;
        weights1[28163] <= 16'b1111111111110010;
        weights1[28164] <= 16'b1111111111111000;
        weights1[28165] <= 16'b1111111111111010;
        weights1[28166] <= 16'b1111111111111111;
        weights1[28167] <= 16'b1111111111111101;
        weights1[28168] <= 16'b0000000000000001;
        weights1[28169] <= 16'b0000000000000001;
        weights1[28170] <= 16'b0000000000000001;
        weights1[28171] <= 16'b0000000000000010;
        weights1[28172] <= 16'b1111111111111111;
        weights1[28173] <= 16'b1111111111111010;
        weights1[28174] <= 16'b1111111111111100;
        weights1[28175] <= 16'b1111111111111111;
        weights1[28176] <= 16'b1111111111101111;
        weights1[28177] <= 16'b1111111111111000;
        weights1[28178] <= 16'b1111111111111010;
        weights1[28179] <= 16'b1111111111110100;
        weights1[28180] <= 16'b1111111111110111;
        weights1[28181] <= 16'b1111111111110011;
        weights1[28182] <= 16'b1111111111111010;
        weights1[28183] <= 16'b1111111111111110;
        weights1[28184] <= 16'b1111111111101110;
        weights1[28185] <= 16'b1111111111111000;
        weights1[28186] <= 16'b1111111111111010;
        weights1[28187] <= 16'b1111111111110000;
        weights1[28188] <= 16'b1111111111101000;
        weights1[28189] <= 16'b1111111111111100;
        weights1[28190] <= 16'b1111111111111100;
        weights1[28191] <= 16'b1111111111111011;
        weights1[28192] <= 16'b1111111111111010;
        weights1[28193] <= 16'b1111111111111011;
        weights1[28194] <= 16'b1111111111111111;
        weights1[28195] <= 16'b0000000000000000;
        weights1[28196] <= 16'b0000000000000000;
        weights1[28197] <= 16'b0000000000000000;
        weights1[28198] <= 16'b0000000000000001;
        weights1[28199] <= 16'b0000000000000001;
        weights1[28200] <= 16'b1111111111111100;
        weights1[28201] <= 16'b1111111111111101;
        weights1[28202] <= 16'b0000000000000000;
        weights1[28203] <= 16'b1111111111110010;
        weights1[28204] <= 16'b1111111111110010;
        weights1[28205] <= 16'b1111111111111100;
        weights1[28206] <= 16'b1111111111110111;
        weights1[28207] <= 16'b1111111111111001;
        weights1[28208] <= 16'b1111111111111100;
        weights1[28209] <= 16'b1111111111111111;
        weights1[28210] <= 16'b1111111111111010;
        weights1[28211] <= 16'b1111111111110111;
        weights1[28212] <= 16'b1111111111111001;
        weights1[28213] <= 16'b0000000000000000;
        weights1[28214] <= 16'b1111111111111111;
        weights1[28215] <= 16'b0000000000000000;
        weights1[28216] <= 16'b0000000000000000;
        weights1[28217] <= 16'b0000000000000000;
        weights1[28218] <= 16'b0000000000000000;
        weights1[28219] <= 16'b1111111111111110;
        weights1[28220] <= 16'b1111111111111100;
        weights1[28221] <= 16'b1111111111111110;
        weights1[28222] <= 16'b0000000000000001;
        weights1[28223] <= 16'b0000000000000000;
        weights1[28224] <= 16'b0000000000000000;
        weights1[28225] <= 16'b0000000000000000;
        weights1[28226] <= 16'b0000000000000000;
        weights1[28227] <= 16'b0000000000000010;
        weights1[28228] <= 16'b0000000000000000;
        weights1[28229] <= 16'b1111111111111101;
        weights1[28230] <= 16'b1111111111111011;
        weights1[28231] <= 16'b1111111111111111;
        weights1[28232] <= 16'b1111111111111101;
        weights1[28233] <= 16'b1111111111111101;
        weights1[28234] <= 16'b1111111111111010;
        weights1[28235] <= 16'b0000000000000010;
        weights1[28236] <= 16'b1111111111111110;
        weights1[28237] <= 16'b1111111111111010;
        weights1[28238] <= 16'b1111111111111101;
        weights1[28239] <= 16'b1111111111111011;
        weights1[28240] <= 16'b1111111111110110;
        weights1[28241] <= 16'b1111111111110011;
        weights1[28242] <= 16'b1111111111101101;
        weights1[28243] <= 16'b1111111111101101;
        weights1[28244] <= 16'b1111111111110001;
        weights1[28245] <= 16'b1111111111111010;
        weights1[28246] <= 16'b0000000000000000;
        weights1[28247] <= 16'b0000000000000000;
        weights1[28248] <= 16'b0000000000000001;
        weights1[28249] <= 16'b0000000000000000;
        weights1[28250] <= 16'b0000000000000000;
        weights1[28251] <= 16'b0000000000000000;
        weights1[28252] <= 16'b0000000000000000;
        weights1[28253] <= 16'b0000000000000000;
        weights1[28254] <= 16'b1111111111111100;
        weights1[28255] <= 16'b1111111111111101;
        weights1[28256] <= 16'b1111111111111100;
        weights1[28257] <= 16'b1111111111110111;
        weights1[28258] <= 16'b1111111111111010;
        weights1[28259] <= 16'b1111111111111111;
        weights1[28260] <= 16'b1111111111111011;
        weights1[28261] <= 16'b1111111111111101;
        weights1[28262] <= 16'b1111111111111100;
        weights1[28263] <= 16'b0000000000000011;
        weights1[28264] <= 16'b1111111111111101;
        weights1[28265] <= 16'b1111111111111100;
        weights1[28266] <= 16'b0000000000000000;
        weights1[28267] <= 16'b1111111111111010;
        weights1[28268] <= 16'b1111111111111101;
        weights1[28269] <= 16'b1111111111100011;
        weights1[28270] <= 16'b1111111111111100;
        weights1[28271] <= 16'b1111111111101110;
        weights1[28272] <= 16'b1111111111111101;
        weights1[28273] <= 16'b1111111111111110;
        weights1[28274] <= 16'b1111111111111101;
        weights1[28275] <= 16'b0000000000000000;
        weights1[28276] <= 16'b1111111111111110;
        weights1[28277] <= 16'b0000000000000011;
        weights1[28278] <= 16'b1111111111111101;
        weights1[28279] <= 16'b0000000000000000;
        weights1[28280] <= 16'b0000000000000001;
        weights1[28281] <= 16'b1111111111111100;
        weights1[28282] <= 16'b1111111111111001;
        weights1[28283] <= 16'b1111111111111000;
        weights1[28284] <= 16'b1111111111110010;
        weights1[28285] <= 16'b1111111111110001;
        weights1[28286] <= 16'b1111111111110100;
        weights1[28287] <= 16'b1111111111111110;
        weights1[28288] <= 16'b1111111111110111;
        weights1[28289] <= 16'b1111111111111100;
        weights1[28290] <= 16'b0000000000001111;
        weights1[28291] <= 16'b0000000000000001;
        weights1[28292] <= 16'b1111111111111110;
        weights1[28293] <= 16'b0000000000000111;
        weights1[28294] <= 16'b0000000000000110;
        weights1[28295] <= 16'b1111111111111111;
        weights1[28296] <= 16'b0000000000000000;
        weights1[28297] <= 16'b0000000000001001;
        weights1[28298] <= 16'b0000000000000100;
        weights1[28299] <= 16'b0000000000001011;
        weights1[28300] <= 16'b1111111111111100;
        weights1[28301] <= 16'b1111111111111100;
        weights1[28302] <= 16'b1111111111110110;
        weights1[28303] <= 16'b1111111111110010;
        weights1[28304] <= 16'b1111111111111011;
        weights1[28305] <= 16'b0000000000000011;
        weights1[28306] <= 16'b0000000000000000;
        weights1[28307] <= 16'b1111111111111011;
        weights1[28308] <= 16'b0000000000000001;
        weights1[28309] <= 16'b0000000000000000;
        weights1[28310] <= 16'b1111111111111011;
        weights1[28311] <= 16'b1111111111110110;
        weights1[28312] <= 16'b1111111111110001;
        weights1[28313] <= 16'b1111111111110100;
        weights1[28314] <= 16'b1111111111110001;
        weights1[28315] <= 16'b1111111111111000;
        weights1[28316] <= 16'b1111111111111001;
        weights1[28317] <= 16'b1111111111111001;
        weights1[28318] <= 16'b1111111111111111;
        weights1[28319] <= 16'b1111111111111100;
        weights1[28320] <= 16'b0000000000000110;
        weights1[28321] <= 16'b0000000000000011;
        weights1[28322] <= 16'b0000000000000110;
        weights1[28323] <= 16'b1111111111111001;
        weights1[28324] <= 16'b1111111111110011;
        weights1[28325] <= 16'b1111111111111110;
        weights1[28326] <= 16'b0000000000000111;
        weights1[28327] <= 16'b0000000000001001;
        weights1[28328] <= 16'b0000000000001000;
        weights1[28329] <= 16'b1111111111111001;
        weights1[28330] <= 16'b1111111111110001;
        weights1[28331] <= 16'b1111111111110011;
        weights1[28332] <= 16'b1111111111110110;
        weights1[28333] <= 16'b0000000000000101;
        weights1[28334] <= 16'b0000000000000010;
        weights1[28335] <= 16'b1111111111111110;
        weights1[28336] <= 16'b1111111111111110;
        weights1[28337] <= 16'b1111111111111100;
        weights1[28338] <= 16'b1111111111110101;
        weights1[28339] <= 16'b1111111111101011;
        weights1[28340] <= 16'b1111111111101111;
        weights1[28341] <= 16'b1111111111100110;
        weights1[28342] <= 16'b1111111111110101;
        weights1[28343] <= 16'b1111111111101101;
        weights1[28344] <= 16'b1111111111111100;
        weights1[28345] <= 16'b1111111111111111;
        weights1[28346] <= 16'b0000000000000001;
        weights1[28347] <= 16'b1111111111111000;
        weights1[28348] <= 16'b1111111111110011;
        weights1[28349] <= 16'b1111111111111010;
        weights1[28350] <= 16'b1111111111111111;
        weights1[28351] <= 16'b0000000000000001;
        weights1[28352] <= 16'b0000000000000001;
        weights1[28353] <= 16'b0000000000000110;
        weights1[28354] <= 16'b1111111111111001;
        weights1[28355] <= 16'b1111111111110111;
        weights1[28356] <= 16'b1111111111110110;
        weights1[28357] <= 16'b1111111111110101;
        weights1[28358] <= 16'b1111111111110111;
        weights1[28359] <= 16'b1111111111110010;
        weights1[28360] <= 16'b1111111111101110;
        weights1[28361] <= 16'b0000000000001001;
        weights1[28362] <= 16'b0000000000000001;
        weights1[28363] <= 16'b0000000000000011;
        weights1[28364] <= 16'b1111111111111101;
        weights1[28365] <= 16'b1111111111111100;
        weights1[28366] <= 16'b1111111111110111;
        weights1[28367] <= 16'b1111111111101111;
        weights1[28368] <= 16'b1111111111100110;
        weights1[28369] <= 16'b1111111111110100;
        weights1[28370] <= 16'b1111111111110111;
        weights1[28371] <= 16'b0000000000000011;
        weights1[28372] <= 16'b1111111111110101;
        weights1[28373] <= 16'b1111111111111000;
        weights1[28374] <= 16'b1111111111100010;
        weights1[28375] <= 16'b1111111111110110;
        weights1[28376] <= 16'b1111111111111110;
        weights1[28377] <= 16'b1111111111011010;
        weights1[28378] <= 16'b0000000000010010;
        weights1[28379] <= 16'b0000000000000001;
        weights1[28380] <= 16'b1111111111111000;
        weights1[28381] <= 16'b1111111111101000;
        weights1[28382] <= 16'b1111111111111001;
        weights1[28383] <= 16'b1111111111111001;
        weights1[28384] <= 16'b0000000000000111;
        weights1[28385] <= 16'b1111111111111110;
        weights1[28386] <= 16'b0000000000010110;
        weights1[28387] <= 16'b1111111111110001;
        weights1[28388] <= 16'b1111111111110111;
        weights1[28389] <= 16'b0000000000000011;
        weights1[28390] <= 16'b1111111111111000;
        weights1[28391] <= 16'b0000000000000000;
        weights1[28392] <= 16'b1111111111111110;
        weights1[28393] <= 16'b1111111111111111;
        weights1[28394] <= 16'b1111111111111011;
        weights1[28395] <= 16'b1111111111110011;
        weights1[28396] <= 16'b1111111111100101;
        weights1[28397] <= 16'b1111111111101010;
        weights1[28398] <= 16'b0000000000000000;
        weights1[28399] <= 16'b1111111111110000;
        weights1[28400] <= 16'b0000000000001100;
        weights1[28401] <= 16'b1111111111111100;
        weights1[28402] <= 16'b1111111111110111;
        weights1[28403] <= 16'b1111111111110000;
        weights1[28404] <= 16'b1111111111101111;
        weights1[28405] <= 16'b1111111111111101;
        weights1[28406] <= 16'b1111111111101111;
        weights1[28407] <= 16'b0000000000000000;
        weights1[28408] <= 16'b1111111111111100;
        weights1[28409] <= 16'b0000000000000001;
        weights1[28410] <= 16'b0000000000001000;
        weights1[28411] <= 16'b0000000000000010;
        weights1[28412] <= 16'b0000000000001000;
        weights1[28413] <= 16'b1111111111111101;
        weights1[28414] <= 16'b1111111111111111;
        weights1[28415] <= 16'b1111111111110011;
        weights1[28416] <= 16'b0000000000001101;
        weights1[28417] <= 16'b0000000000000111;
        weights1[28418] <= 16'b1111111111111101;
        weights1[28419] <= 16'b0000000000000000;
        weights1[28420] <= 16'b1111111111111110;
        weights1[28421] <= 16'b1111111111110111;
        weights1[28422] <= 16'b1111111111111010;
        weights1[28423] <= 16'b1111111111110001;
        weights1[28424] <= 16'b1111111111101001;
        weights1[28425] <= 16'b1111111111110001;
        weights1[28426] <= 16'b1111111111110111;
        weights1[28427] <= 16'b0000000000001100;
        weights1[28428] <= 16'b0000000000001101;
        weights1[28429] <= 16'b0000000000000001;
        weights1[28430] <= 16'b0000000000001000;
        weights1[28431] <= 16'b1111111111110101;
        weights1[28432] <= 16'b1111111111110100;
        weights1[28433] <= 16'b0000000000000000;
        weights1[28434] <= 16'b1111111111110010;
        weights1[28435] <= 16'b0000000000010010;
        weights1[28436] <= 16'b0000000000010100;
        weights1[28437] <= 16'b0000000000010111;
        weights1[28438] <= 16'b1111111111111101;
        weights1[28439] <= 16'b0000000000000110;
        weights1[28440] <= 16'b0000000000000111;
        weights1[28441] <= 16'b1111111111110010;
        weights1[28442] <= 16'b1111111111111010;
        weights1[28443] <= 16'b0000000000000110;
        weights1[28444] <= 16'b1111111111110101;
        weights1[28445] <= 16'b0000000000001010;
        weights1[28446] <= 16'b1111111111101111;
        weights1[28447] <= 16'b1111111111111110;
        weights1[28448] <= 16'b1111111111111001;
        weights1[28449] <= 16'b1111111111110010;
        weights1[28450] <= 16'b1111111111111101;
        weights1[28451] <= 16'b1111111111110010;
        weights1[28452] <= 16'b1111111111111110;
        weights1[28453] <= 16'b1111111111111000;
        weights1[28454] <= 16'b1111111111111100;
        weights1[28455] <= 16'b0000000000000001;
        weights1[28456] <= 16'b0000000000000001;
        weights1[28457] <= 16'b0000000000000100;
        weights1[28458] <= 16'b0000000000001011;
        weights1[28459] <= 16'b0000000000001100;
        weights1[28460] <= 16'b1111111111110101;
        weights1[28461] <= 16'b0000000000001011;
        weights1[28462] <= 16'b1111111111110101;
        weights1[28463] <= 16'b1111111111111101;
        weights1[28464] <= 16'b1111111111111111;
        weights1[28465] <= 16'b1111111111101011;
        weights1[28466] <= 16'b0000000000000010;
        weights1[28467] <= 16'b0000000000100001;
        weights1[28468] <= 16'b0000000000000010;
        weights1[28469] <= 16'b1111111111101001;
        weights1[28470] <= 16'b1111111111110000;
        weights1[28471] <= 16'b0000000000000100;
        weights1[28472] <= 16'b0000000000000100;
        weights1[28473] <= 16'b1111111111110001;
        weights1[28474] <= 16'b0000000000001010;
        weights1[28475] <= 16'b0000000000001110;
        weights1[28476] <= 16'b1111111111110100;
        weights1[28477] <= 16'b0000000000000000;
        weights1[28478] <= 16'b0000000000000101;
        weights1[28479] <= 16'b1111111111110111;
        weights1[28480] <= 16'b1111111111101001;
        weights1[28481] <= 16'b1111111111100110;
        weights1[28482] <= 16'b1111111111110110;
        weights1[28483] <= 16'b1111111111110000;
        weights1[28484] <= 16'b1111111111111000;
        weights1[28485] <= 16'b0000000000001111;
        weights1[28486] <= 16'b0000000000000101;
        weights1[28487] <= 16'b0000000000000011;
        weights1[28488] <= 16'b0000000000000001;
        weights1[28489] <= 16'b1111111111101011;
        weights1[28490] <= 16'b1111111111101100;
        weights1[28491] <= 16'b1111111111111110;
        weights1[28492] <= 16'b0000000000001111;
        weights1[28493] <= 16'b0000000000010011;
        weights1[28494] <= 16'b0000000000001100;
        weights1[28495] <= 16'b0000000000001001;
        weights1[28496] <= 16'b0000000000011000;
        weights1[28497] <= 16'b0000000000011100;
        weights1[28498] <= 16'b1111111111111011;
        weights1[28499] <= 16'b0000000000010100;
        weights1[28500] <= 16'b1111111111111110;
        weights1[28501] <= 16'b1111111111111010;
        weights1[28502] <= 16'b0000000000000001;
        weights1[28503] <= 16'b0000000000000000;
        weights1[28504] <= 16'b1111111111111011;
        weights1[28505] <= 16'b0000000000000111;
        weights1[28506] <= 16'b1111111111111011;
        weights1[28507] <= 16'b1111111111110101;
        weights1[28508] <= 16'b1111111111110000;
        weights1[28509] <= 16'b1111111111110101;
        weights1[28510] <= 16'b1111111111101001;
        weights1[28511] <= 16'b1111111111111100;
        weights1[28512] <= 16'b1111111111110000;
        weights1[28513] <= 16'b1111111111110110;
        weights1[28514] <= 16'b1111111111111111;
        weights1[28515] <= 16'b0000000000010011;
        weights1[28516] <= 16'b1111111111101001;
        weights1[28517] <= 16'b1111111111011001;
        weights1[28518] <= 16'b0000000000000011;
        weights1[28519] <= 16'b0000000000000000;
        weights1[28520] <= 16'b0000000000000010;
        weights1[28521] <= 16'b0000000000001110;
        weights1[28522] <= 16'b0000000000000111;
        weights1[28523] <= 16'b0000000000000110;
        weights1[28524] <= 16'b0000000000001100;
        weights1[28525] <= 16'b0000000000010011;
        weights1[28526] <= 16'b0000000000010111;
        weights1[28527] <= 16'b0000000000011101;
        weights1[28528] <= 16'b0000000000010100;
        weights1[28529] <= 16'b0000000000001110;
        weights1[28530] <= 16'b0000000000001011;
        weights1[28531] <= 16'b0000000000001100;
        weights1[28532] <= 16'b1111111111111101;
        weights1[28533] <= 16'b1111111111111101;
        weights1[28534] <= 16'b0000000000000000;
        weights1[28535] <= 16'b1111111111101100;
        weights1[28536] <= 16'b1111111111100011;
        weights1[28537] <= 16'b1111111111100110;
        weights1[28538] <= 16'b0000000000001001;
        weights1[28539] <= 16'b1111111111110111;
        weights1[28540] <= 16'b0000000000000111;
        weights1[28541] <= 16'b0000000000010110;
        weights1[28542] <= 16'b0000000000010111;
        weights1[28543] <= 16'b0000000000001000;
        weights1[28544] <= 16'b0000000000000001;
        weights1[28545] <= 16'b1111111111101011;
        weights1[28546] <= 16'b1111111111110101;
        weights1[28547] <= 16'b1111111111100101;
        weights1[28548] <= 16'b0000000000000000;
        weights1[28549] <= 16'b0000000000000101;
        weights1[28550] <= 16'b0000000000000110;
        weights1[28551] <= 16'b0000000000001110;
        weights1[28552] <= 16'b0000000000000100;
        weights1[28553] <= 16'b0000000000000111;
        weights1[28554] <= 16'b0000000000011100;
        weights1[28555] <= 16'b0000000000100011;
        weights1[28556] <= 16'b0000000000100110;
        weights1[28557] <= 16'b0000000000011000;
        weights1[28558] <= 16'b0000000000011000;
        weights1[28559] <= 16'b0000000000010000;
        weights1[28560] <= 16'b1111111111111111;
        weights1[28561] <= 16'b0000000000001011;
        weights1[28562] <= 16'b1111111111111100;
        weights1[28563] <= 16'b1111111111111000;
        weights1[28564] <= 16'b1111111111110010;
        weights1[28565] <= 16'b1111111111100011;
        weights1[28566] <= 16'b1111111111110001;
        weights1[28567] <= 16'b1111111111111100;
        weights1[28568] <= 16'b0000000000000111;
        weights1[28569] <= 16'b0000000000001000;
        weights1[28570] <= 16'b0000000000010111;
        weights1[28571] <= 16'b0000000000001000;
        weights1[28572] <= 16'b0000000000001010;
        weights1[28573] <= 16'b1111111111110110;
        weights1[28574] <= 16'b1111111111001101;
        weights1[28575] <= 16'b1111111111101101;
        weights1[28576] <= 16'b1111111111101010;
        weights1[28577] <= 16'b0000000000000100;
        weights1[28578] <= 16'b0000000000000101;
        weights1[28579] <= 16'b0000000000011101;
        weights1[28580] <= 16'b0000000000010101;
        weights1[28581] <= 16'b0000000000000000;
        weights1[28582] <= 16'b0000000000000101;
        weights1[28583] <= 16'b0000000000011110;
        weights1[28584] <= 16'b0000000000100011;
        weights1[28585] <= 16'b0000000000001111;
        weights1[28586] <= 16'b0000000000010110;
        weights1[28587] <= 16'b0000000000001001;
        weights1[28588] <= 16'b1111111111111100;
        weights1[28589] <= 16'b0000000000001100;
        weights1[28590] <= 16'b0000000000010000;
        weights1[28591] <= 16'b0000000000000010;
        weights1[28592] <= 16'b1111111111110011;
        weights1[28593] <= 16'b1111111111111110;
        weights1[28594] <= 16'b1111111111110101;
        weights1[28595] <= 16'b1111111111100110;
        weights1[28596] <= 16'b0000000000001100;
        weights1[28597] <= 16'b0000000000001010;
        weights1[28598] <= 16'b0000000000100001;
        weights1[28599] <= 16'b0000000000101000;
        weights1[28600] <= 16'b1111111111111111;
        weights1[28601] <= 16'b1111111111010000;
        weights1[28602] <= 16'b1111111111001101;
        weights1[28603] <= 16'b1111111111011000;
        weights1[28604] <= 16'b1111111111110101;
        weights1[28605] <= 16'b0000000000011001;
        weights1[28606] <= 16'b0000000000100001;
        weights1[28607] <= 16'b0000000000010000;
        weights1[28608] <= 16'b0000000000100001;
        weights1[28609] <= 16'b0000000000110000;
        weights1[28610] <= 16'b0000000000110111;
        weights1[28611] <= 16'b0000000000111010;
        weights1[28612] <= 16'b0000000000011110;
        weights1[28613] <= 16'b0000000000001100;
        weights1[28614] <= 16'b0000000000001000;
        weights1[28615] <= 16'b1111111111111000;
        weights1[28616] <= 16'b0000000000001001;
        weights1[28617] <= 16'b0000000000000111;
        weights1[28618] <= 16'b0000000000010001;
        weights1[28619] <= 16'b0000000000000100;
        weights1[28620] <= 16'b1111111111111100;
        weights1[28621] <= 16'b1111111111110010;
        weights1[28622] <= 16'b1111111111110110;
        weights1[28623] <= 16'b0000000000001100;
        weights1[28624] <= 16'b0000000000010000;
        weights1[28625] <= 16'b0000000000011001;
        weights1[28626] <= 16'b0000000000011010;
        weights1[28627] <= 16'b0000000000001100;
        weights1[28628] <= 16'b1111111111110110;
        weights1[28629] <= 16'b1111111111101001;
        weights1[28630] <= 16'b1111111110100110;
        weights1[28631] <= 16'b1111111110110110;
        weights1[28632] <= 16'b1111111111101000;
        weights1[28633] <= 16'b1111111111101100;
        weights1[28634] <= 16'b1111111111111001;
        weights1[28635] <= 16'b0000000000100010;
        weights1[28636] <= 16'b0000000000100111;
        weights1[28637] <= 16'b0000000000110001;
        weights1[28638] <= 16'b0000000000010110;
        weights1[28639] <= 16'b0000000000011111;
        weights1[28640] <= 16'b0000000000001101;
        weights1[28641] <= 16'b1111111111111100;
        weights1[28642] <= 16'b1111111111110001;
        weights1[28643] <= 16'b1111111111101110;
        weights1[28644] <= 16'b0000000000010010;
        weights1[28645] <= 16'b0000000000000100;
        weights1[28646] <= 16'b0000000000010000;
        weights1[28647] <= 16'b0000000000010111;
        weights1[28648] <= 16'b0000000000000111;
        weights1[28649] <= 16'b0000000000001110;
        weights1[28650] <= 16'b1111111111110101;
        weights1[28651] <= 16'b0000000000000111;
        weights1[28652] <= 16'b1111111111111001;
        weights1[28653] <= 16'b0000000000010111;
        weights1[28654] <= 16'b0000000000010100;
        weights1[28655] <= 16'b0000000000100010;
        weights1[28656] <= 16'b0000000000001010;
        weights1[28657] <= 16'b1111111111110100;
        weights1[28658] <= 16'b1111111110111100;
        weights1[28659] <= 16'b1111111110010010;
        weights1[28660] <= 16'b1111111111001000;
        weights1[28661] <= 16'b1111111111011000;
        weights1[28662] <= 16'b0000000000000110;
        weights1[28663] <= 16'b1111111111111010;
        weights1[28664] <= 16'b0000000000001000;
        weights1[28665] <= 16'b0000000000001011;
        weights1[28666] <= 16'b1111111111110000;
        weights1[28667] <= 16'b0000000000000110;
        weights1[28668] <= 16'b1111111111101011;
        weights1[28669] <= 16'b1111111111101101;
        weights1[28670] <= 16'b1111111111101101;
        weights1[28671] <= 16'b1111111111100101;
        weights1[28672] <= 16'b0000000000000101;
        weights1[28673] <= 16'b1111111111111010;
        weights1[28674] <= 16'b0000000000011001;
        weights1[28675] <= 16'b0000000000010011;
        weights1[28676] <= 16'b0000000000000010;
        weights1[28677] <= 16'b0000000000000011;
        weights1[28678] <= 16'b0000000000001111;
        weights1[28679] <= 16'b0000000000010011;
        weights1[28680] <= 16'b0000000000000110;
        weights1[28681] <= 16'b0000000000001101;
        weights1[28682] <= 16'b0000000000011100;
        weights1[28683] <= 16'b0000000000010110;
        weights1[28684] <= 16'b0000000000011011;
        weights1[28685] <= 16'b0000000000000101;
        weights1[28686] <= 16'b1111111111001111;
        weights1[28687] <= 16'b1111111110000111;
        weights1[28688] <= 16'b1111111110001111;
        weights1[28689] <= 16'b1111111110100000;
        weights1[28690] <= 16'b1111111110100111;
        weights1[28691] <= 16'b1111111110111100;
        weights1[28692] <= 16'b1111111110111101;
        weights1[28693] <= 16'b1111111110111000;
        weights1[28694] <= 16'b1111111111001011;
        weights1[28695] <= 16'b1111111111001111;
        weights1[28696] <= 16'b1111111111011010;
        weights1[28697] <= 16'b1111111111010101;
        weights1[28698] <= 16'b1111111111100100;
        weights1[28699] <= 16'b1111111111100110;
        weights1[28700] <= 16'b0000000000000100;
        weights1[28701] <= 16'b0000000000001100;
        weights1[28702] <= 16'b0000000000011010;
        weights1[28703] <= 16'b0000000000010001;
        weights1[28704] <= 16'b0000000000010001;
        weights1[28705] <= 16'b0000000000011010;
        weights1[28706] <= 16'b0000000000001011;
        weights1[28707] <= 16'b0000000000001110;
        weights1[28708] <= 16'b0000000000010111;
        weights1[28709] <= 16'b0000000000010000;
        weights1[28710] <= 16'b0000000000010110;
        weights1[28711] <= 16'b0000000000011011;
        weights1[28712] <= 16'b0000000000000110;
        weights1[28713] <= 16'b0000000000010010;
        weights1[28714] <= 16'b1111111111100101;
        weights1[28715] <= 16'b1111111110010100;
        weights1[28716] <= 16'b1111111101110110;
        weights1[28717] <= 16'b1111111101101111;
        weights1[28718] <= 16'b1111111101111111;
        weights1[28719] <= 16'b1111111110011001;
        weights1[28720] <= 16'b1111111110100001;
        weights1[28721] <= 16'b1111111110101010;
        weights1[28722] <= 16'b1111111111000111;
        weights1[28723] <= 16'b1111111111001010;
        weights1[28724] <= 16'b1111111111001101;
        weights1[28725] <= 16'b1111111111010001;
        weights1[28726] <= 16'b1111111111100001;
        weights1[28727] <= 16'b1111111111100111;
        weights1[28728] <= 16'b1111111111111000;
        weights1[28729] <= 16'b0000000000010111;
        weights1[28730] <= 16'b0000000000100100;
        weights1[28731] <= 16'b0000000000001011;
        weights1[28732] <= 16'b0000000000000000;
        weights1[28733] <= 16'b0000000000010011;
        weights1[28734] <= 16'b0000000000000101;
        weights1[28735] <= 16'b1111111111111110;
        weights1[28736] <= 16'b0000000000000110;
        weights1[28737] <= 16'b0000000000001100;
        weights1[28738] <= 16'b0000000000001100;
        weights1[28739] <= 16'b0000000000011001;
        weights1[28740] <= 16'b0000000000010001;
        weights1[28741] <= 16'b0000000000011001;
        weights1[28742] <= 16'b1111111111101010;
        weights1[28743] <= 16'b1111111111001000;
        weights1[28744] <= 16'b1111111101110111;
        weights1[28745] <= 16'b1111111101001110;
        weights1[28746] <= 16'b1111111110000001;
        weights1[28747] <= 16'b1111111110011100;
        weights1[28748] <= 16'b1111111110101010;
        weights1[28749] <= 16'b1111111111001000;
        weights1[28750] <= 16'b1111111111000100;
        weights1[28751] <= 16'b1111111111010010;
        weights1[28752] <= 16'b1111111111010001;
        weights1[28753] <= 16'b1111111111011011;
        weights1[28754] <= 16'b1111111111100001;
        weights1[28755] <= 16'b1111111111101000;
        weights1[28756] <= 16'b1111111111111001;
        weights1[28757] <= 16'b0000000000000000;
        weights1[28758] <= 16'b0000000000000100;
        weights1[28759] <= 16'b0000000000000100;
        weights1[28760] <= 16'b1111111111111100;
        weights1[28761] <= 16'b1111111111111110;
        weights1[28762] <= 16'b0000000000001010;
        weights1[28763] <= 16'b0000000000010001;
        weights1[28764] <= 16'b0000000000010011;
        weights1[28765] <= 16'b0000000000000110;
        weights1[28766] <= 16'b0000000000010000;
        weights1[28767] <= 16'b0000000000001111;
        weights1[28768] <= 16'b0000000000010000;
        weights1[28769] <= 16'b0000000000100101;
        weights1[28770] <= 16'b0000000000100010;
        weights1[28771] <= 16'b0000000000001001;
        weights1[28772] <= 16'b1111111110101111;
        weights1[28773] <= 16'b1111111101110101;
        weights1[28774] <= 16'b1111111110000010;
        weights1[28775] <= 16'b1111111110011110;
        weights1[28776] <= 16'b1111111110110010;
        weights1[28777] <= 16'b1111111111000001;
        weights1[28778] <= 16'b1111111111001011;
        weights1[28779] <= 16'b1111111111010000;
        weights1[28780] <= 16'b1111111111010110;
        weights1[28781] <= 16'b1111111111011101;
        weights1[28782] <= 16'b1111111111100101;
        weights1[28783] <= 16'b1111111111101101;
        weights1[28784] <= 16'b1111111111111100;
        weights1[28785] <= 16'b0000000000000011;
        weights1[28786] <= 16'b1111111111111111;
        weights1[28787] <= 16'b0000000000011001;
        weights1[28788] <= 16'b0000000000010010;
        weights1[28789] <= 16'b0000000000001011;
        weights1[28790] <= 16'b1111111111110101;
        weights1[28791] <= 16'b0000000000011010;
        weights1[28792] <= 16'b0000000000000011;
        weights1[28793] <= 16'b0000000000001100;
        weights1[28794] <= 16'b0000000000001111;
        weights1[28795] <= 16'b0000000000001000;
        weights1[28796] <= 16'b0000000000100011;
        weights1[28797] <= 16'b0000000000011111;
        weights1[28798] <= 16'b0000000000101101;
        weights1[28799] <= 16'b0000000000101110;
        weights1[28800] <= 16'b1111111111110100;
        weights1[28801] <= 16'b1111111110011101;
        weights1[28802] <= 16'b1111111110001011;
        weights1[28803] <= 16'b1111111110011100;
        weights1[28804] <= 16'b1111111110111001;
        weights1[28805] <= 16'b1111111111001000;
        weights1[28806] <= 16'b1111111111010100;
        weights1[28807] <= 16'b1111111111011010;
        weights1[28808] <= 16'b1111111111011101;
        weights1[28809] <= 16'b1111111111011111;
        weights1[28810] <= 16'b1111111111100110;
        weights1[28811] <= 16'b1111111111101011;
        weights1[28812] <= 16'b1111111111110111;
        weights1[28813] <= 16'b0000000000001101;
        weights1[28814] <= 16'b0000000000010100;
        weights1[28815] <= 16'b0000000000001100;
        weights1[28816] <= 16'b1111111111110101;
        weights1[28817] <= 16'b0000000000011101;
        weights1[28818] <= 16'b0000000000001101;
        weights1[28819] <= 16'b0000000000011101;
        weights1[28820] <= 16'b0000000000001111;
        weights1[28821] <= 16'b0000000000010000;
        weights1[28822] <= 16'b0000000000001101;
        weights1[28823] <= 16'b0000000000001001;
        weights1[28824] <= 16'b0000000000010001;
        weights1[28825] <= 16'b0000000000011010;
        weights1[28826] <= 16'b0000000000010001;
        weights1[28827] <= 16'b0000000000111000;
        weights1[28828] <= 16'b0000000000000100;
        weights1[28829] <= 16'b1111111110111000;
        weights1[28830] <= 16'b1111111110011010;
        weights1[28831] <= 16'b1111111110100010;
        weights1[28832] <= 16'b1111111110111110;
        weights1[28833] <= 16'b1111111111001111;
        weights1[28834] <= 16'b1111111111010111;
        weights1[28835] <= 16'b1111111111011010;
        weights1[28836] <= 16'b1111111111100001;
        weights1[28837] <= 16'b1111111111100011;
        weights1[28838] <= 16'b1111111111101110;
        weights1[28839] <= 16'b1111111111100110;
        weights1[28840] <= 16'b1111111111111001;
        weights1[28841] <= 16'b0000000000000101;
        weights1[28842] <= 16'b0000000000010011;
        weights1[28843] <= 16'b0000000000010001;
        weights1[28844] <= 16'b0000000000001000;
        weights1[28845] <= 16'b0000000000000100;
        weights1[28846] <= 16'b0000000000010100;
        weights1[28847] <= 16'b0000000000001101;
        weights1[28848] <= 16'b1111111111110100;
        weights1[28849] <= 16'b0000000000001001;
        weights1[28850] <= 16'b0000000000000101;
        weights1[28851] <= 16'b0000000000000111;
        weights1[28852] <= 16'b0000000000011001;
        weights1[28853] <= 16'b0000000000000010;
        weights1[28854] <= 16'b0000000000010111;
        weights1[28855] <= 16'b0000000000100101;
        weights1[28856] <= 16'b0000000000101010;
        weights1[28857] <= 16'b1111111111010111;
        weights1[28858] <= 16'b1111111110111000;
        weights1[28859] <= 16'b1111111110101101;
        weights1[28860] <= 16'b1111111111001010;
        weights1[28861] <= 16'b1111111111010000;
        weights1[28862] <= 16'b1111111111011010;
        weights1[28863] <= 16'b1111111111011110;
        weights1[28864] <= 16'b1111111111100100;
        weights1[28865] <= 16'b1111111111100101;
        weights1[28866] <= 16'b1111111111100110;
        weights1[28867] <= 16'b1111111111101101;
        weights1[28868] <= 16'b1111111111111101;
        weights1[28869] <= 16'b0000000000010000;
        weights1[28870] <= 16'b0000000000001100;
        weights1[28871] <= 16'b0000000000001011;
        weights1[28872] <= 16'b0000000000010001;
        weights1[28873] <= 16'b0000000000010111;
        weights1[28874] <= 16'b1111111111111101;
        weights1[28875] <= 16'b0000000000001001;
        weights1[28876] <= 16'b1111111111111010;
        weights1[28877] <= 16'b0000000000010110;
        weights1[28878] <= 16'b0000000000010110;
        weights1[28879] <= 16'b0000000000010000;
        weights1[28880] <= 16'b0000000000000011;
        weights1[28881] <= 16'b0000000000000111;
        weights1[28882] <= 16'b0000000000011110;
        weights1[28883] <= 16'b0000000000010100;
        weights1[28884] <= 16'b0000000000101001;
        weights1[28885] <= 16'b1111111111011000;
        weights1[28886] <= 16'b1111111110111001;
        weights1[28887] <= 16'b1111111110111001;
        weights1[28888] <= 16'b1111111111001100;
        weights1[28889] <= 16'b1111111111001111;
        weights1[28890] <= 16'b1111111111011011;
        weights1[28891] <= 16'b1111111111100000;
        weights1[28892] <= 16'b1111111111100001;
        weights1[28893] <= 16'b1111111111100101;
        weights1[28894] <= 16'b1111111111101011;
        weights1[28895] <= 16'b1111111111110000;
        weights1[28896] <= 16'b1111111111111000;
        weights1[28897] <= 16'b0000000000000101;
        weights1[28898] <= 16'b0000000000010001;
        weights1[28899] <= 16'b0000000000010100;
        weights1[28900] <= 16'b0000000000010101;
        weights1[28901] <= 16'b0000000000011011;
        weights1[28902] <= 16'b0000000000001000;
        weights1[28903] <= 16'b0000000000010100;
        weights1[28904] <= 16'b0000000000000101;
        weights1[28905] <= 16'b0000000000001001;
        weights1[28906] <= 16'b0000000000011101;
        weights1[28907] <= 16'b0000000000010111;
        weights1[28908] <= 16'b0000000000010110;
        weights1[28909] <= 16'b0000000000010110;
        weights1[28910] <= 16'b0000000000100000;
        weights1[28911] <= 16'b0000000000111101;
        weights1[28912] <= 16'b0000000000011111;
        weights1[28913] <= 16'b1111111111110110;
        weights1[28914] <= 16'b1111111111010001;
        weights1[28915] <= 16'b1111111111001000;
        weights1[28916] <= 16'b1111111111010010;
        weights1[28917] <= 16'b1111111111100000;
        weights1[28918] <= 16'b1111111111100101;
        weights1[28919] <= 16'b1111111111100011;
        weights1[28920] <= 16'b1111111111100100;
        weights1[28921] <= 16'b1111111111101010;
        weights1[28922] <= 16'b1111111111110000;
        weights1[28923] <= 16'b1111111111111001;
        weights1[28924] <= 16'b0000000000000011;
        weights1[28925] <= 16'b0000000000001001;
        weights1[28926] <= 16'b0000000000001001;
        weights1[28927] <= 16'b0000000000001100;
        weights1[28928] <= 16'b0000000000000111;
        weights1[28929] <= 16'b0000000000010001;
        weights1[28930] <= 16'b0000000000000000;
        weights1[28931] <= 16'b0000000000001010;
        weights1[28932] <= 16'b0000000000010000;
        weights1[28933] <= 16'b1111111111111101;
        weights1[28934] <= 16'b0000000000011110;
        weights1[28935] <= 16'b0000000000010001;
        weights1[28936] <= 16'b0000000000001101;
        weights1[28937] <= 16'b0000000000010000;
        weights1[28938] <= 16'b0000000000010000;
        weights1[28939] <= 16'b0000000000001010;
        weights1[28940] <= 16'b0000000000000001;
        weights1[28941] <= 16'b1111111111100011;
        weights1[28942] <= 16'b1111111111001100;
        weights1[28943] <= 16'b1111111111001010;
        weights1[28944] <= 16'b1111111111011010;
        weights1[28945] <= 16'b1111111111100011;
        weights1[28946] <= 16'b1111111111100000;
        weights1[28947] <= 16'b1111111111011111;
        weights1[28948] <= 16'b1111111111101101;
        weights1[28949] <= 16'b1111111111110101;
        weights1[28950] <= 16'b1111111111111010;
        weights1[28951] <= 16'b1111111111111111;
        weights1[28952] <= 16'b0000000000000010;
        weights1[28953] <= 16'b0000000000001000;
        weights1[28954] <= 16'b0000000000010010;
        weights1[28955] <= 16'b0000000000001011;
        weights1[28956] <= 16'b1111111111111101;
        weights1[28957] <= 16'b0000000000010000;
        weights1[28958] <= 16'b0000000000000101;
        weights1[28959] <= 16'b0000000000001111;
        weights1[28960] <= 16'b0000000000011000;
        weights1[28961] <= 16'b0000000000010000;
        weights1[28962] <= 16'b0000000000011111;
        weights1[28963] <= 16'b0000000000000101;
        weights1[28964] <= 16'b0000000000010110;
        weights1[28965] <= 16'b0000000000011011;
        weights1[28966] <= 16'b0000000000001111;
        weights1[28967] <= 16'b0000000000010001;
        weights1[28968] <= 16'b1111111111111111;
        weights1[28969] <= 16'b1111111111011110;
        weights1[28970] <= 16'b1111111111100000;
        weights1[28971] <= 16'b1111111111010010;
        weights1[28972] <= 16'b1111111111011100;
        weights1[28973] <= 16'b1111111111011111;
        weights1[28974] <= 16'b1111111111100101;
        weights1[28975] <= 16'b1111111111101101;
        weights1[28976] <= 16'b1111111111110011;
        weights1[28977] <= 16'b1111111111111000;
        weights1[28978] <= 16'b1111111111111101;
        weights1[28979] <= 16'b0000000000000000;
        weights1[28980] <= 16'b0000000000000010;
        weights1[28981] <= 16'b0000000000000000;
        weights1[28982] <= 16'b0000000000000111;
        weights1[28983] <= 16'b0000000000001010;
        weights1[28984] <= 16'b0000000000001110;
        weights1[28985] <= 16'b0000000000001111;
        weights1[28986] <= 16'b0000000000011001;
        weights1[28987] <= 16'b0000000000011010;
        weights1[28988] <= 16'b0000000000010110;
        weights1[28989] <= 16'b0000000000011001;
        weights1[28990] <= 16'b0000000000011011;
        weights1[28991] <= 16'b0000000000100100;
        weights1[28992] <= 16'b0000000000100001;
        weights1[28993] <= 16'b0000000000010111;
        weights1[28994] <= 16'b0000000000000011;
        weights1[28995] <= 16'b1111111111111100;
        weights1[28996] <= 16'b1111111111110001;
        weights1[28997] <= 16'b1111111111100101;
        weights1[28998] <= 16'b1111111111100000;
        weights1[28999] <= 16'b1111111111011111;
        weights1[29000] <= 16'b1111111111100100;
        weights1[29001] <= 16'b1111111111100111;
        weights1[29002] <= 16'b1111111111101111;
        weights1[29003] <= 16'b1111111111110111;
        weights1[29004] <= 16'b1111111111111001;
        weights1[29005] <= 16'b1111111111111110;
        weights1[29006] <= 16'b0000000000000000;
        weights1[29007] <= 16'b0000000000000000;
        weights1[29008] <= 16'b0000000000000000;
        weights1[29009] <= 16'b0000000000000001;
        weights1[29010] <= 16'b0000000000000001;
        weights1[29011] <= 16'b1111111111111110;
        weights1[29012] <= 16'b1111111111111010;
        weights1[29013] <= 16'b1111111111111011;
        weights1[29014] <= 16'b1111111111111100;
        weights1[29015] <= 16'b1111111111111110;
        weights1[29016] <= 16'b1111111111111111;
        weights1[29017] <= 16'b1111111111110001;
        weights1[29018] <= 16'b1111111111101110;
        weights1[29019] <= 16'b1111111111110111;
        weights1[29020] <= 16'b1111111111110110;
        weights1[29021] <= 16'b0000000000000100;
        weights1[29022] <= 16'b0000000000000011;
        weights1[29023] <= 16'b0000000000000101;
        weights1[29024] <= 16'b1111111111111111;
        weights1[29025] <= 16'b1111111111110000;
        weights1[29026] <= 16'b1111111111111010;
        weights1[29027] <= 16'b1111111111111100;
        weights1[29028] <= 16'b0000000000000000;
        weights1[29029] <= 16'b1111111111111101;
        weights1[29030] <= 16'b1111111111111000;
        weights1[29031] <= 16'b1111111111110101;
        weights1[29032] <= 16'b1111111111111110;
        weights1[29033] <= 16'b0000000000000111;
        weights1[29034] <= 16'b0000000000000010;
        weights1[29035] <= 16'b1111111111111110;
        weights1[29036] <= 16'b1111111111111111;
        weights1[29037] <= 16'b0000000000000001;
        weights1[29038] <= 16'b0000000000000000;
        weights1[29039] <= 16'b1111111111111111;
        weights1[29040] <= 16'b1111111111111101;
        weights1[29041] <= 16'b1111111111110111;
        weights1[29042] <= 16'b1111111111111001;
        weights1[29043] <= 16'b1111111111111111;
        weights1[29044] <= 16'b1111111111111111;
        weights1[29045] <= 16'b1111111111110011;
        weights1[29046] <= 16'b1111111111111011;
        weights1[29047] <= 16'b1111111111110010;
        weights1[29048] <= 16'b0000000000000001;
        weights1[29049] <= 16'b0000000000000110;
        weights1[29050] <= 16'b0000000000000100;
        weights1[29051] <= 16'b1111111111111001;
        weights1[29052] <= 16'b1111111111111110;
        weights1[29053] <= 16'b1111111111111000;
        weights1[29054] <= 16'b1111111111110101;
        weights1[29055] <= 16'b0000000000000010;
        weights1[29056] <= 16'b0000000000000110;
        weights1[29057] <= 16'b0000000000000101;
        weights1[29058] <= 16'b1111111111110101;
        weights1[29059] <= 16'b1111111111110111;
        weights1[29060] <= 16'b0000000000000010;
        weights1[29061] <= 16'b0000000000001001;
        weights1[29062] <= 16'b0000000000000000;
        weights1[29063] <= 16'b0000000000000001;
        weights1[29064] <= 16'b0000000000000000;
        weights1[29065] <= 16'b1111111111111101;
        weights1[29066] <= 16'b1111111111111110;
        weights1[29067] <= 16'b0000000000000111;
        weights1[29068] <= 16'b1111111111111001;
        weights1[29069] <= 16'b0000000000000000;
        weights1[29070] <= 16'b1111111111101100;
        weights1[29071] <= 16'b1111111111110010;
        weights1[29072] <= 16'b1111111111111111;
        weights1[29073] <= 16'b0000000000001000;
        weights1[29074] <= 16'b1111111111111110;
        weights1[29075] <= 16'b0000000000000010;
        weights1[29076] <= 16'b1111111111110101;
        weights1[29077] <= 16'b0000000000000110;
        weights1[29078] <= 16'b1111111111110110;
        weights1[29079] <= 16'b0000000000001001;
        weights1[29080] <= 16'b0000000000000000;
        weights1[29081] <= 16'b1111111111111000;
        weights1[29082] <= 16'b1111111111111101;
        weights1[29083] <= 16'b1111111111110101;
        weights1[29084] <= 16'b0000000000000100;
        weights1[29085] <= 16'b1111111111110101;
        weights1[29086] <= 16'b1111111111101110;
        weights1[29087] <= 16'b0000000000000010;
        weights1[29088] <= 16'b0000000000000001;
        weights1[29089] <= 16'b0000000000000001;
        weights1[29090] <= 16'b0000000000001001;
        weights1[29091] <= 16'b1111111111111110;
        weights1[29092] <= 16'b1111111111111111;
        weights1[29093] <= 16'b1111111111111100;
        weights1[29094] <= 16'b0000000000000000;
        weights1[29095] <= 16'b0000000000000000;
        weights1[29096] <= 16'b1111111111110110;
        weights1[29097] <= 16'b1111111111111010;
        weights1[29098] <= 16'b1111111111111110;
        weights1[29099] <= 16'b1111111111111000;
        weights1[29100] <= 16'b1111111111111100;
        weights1[29101] <= 16'b0000000000000000;
        weights1[29102] <= 16'b0000000000001111;
        weights1[29103] <= 16'b1111111111111101;
        weights1[29104] <= 16'b0000000000000110;
        weights1[29105] <= 16'b1111111111110110;
        weights1[29106] <= 16'b0000000000000111;
        weights1[29107] <= 16'b0000000000000111;
        weights1[29108] <= 16'b1111111111110011;
        weights1[29109] <= 16'b0000000000000100;
        weights1[29110] <= 16'b1111111111111101;
        weights1[29111] <= 16'b0000000000001001;
        weights1[29112] <= 16'b1111111111111011;
        weights1[29113] <= 16'b1111111111111100;
        weights1[29114] <= 16'b0000000000000010;
        weights1[29115] <= 16'b0000000000001000;
        weights1[29116] <= 16'b0000000000000111;
        weights1[29117] <= 16'b1111111111111010;
        weights1[29118] <= 16'b0000000000000001;
        weights1[29119] <= 16'b1111111111111110;
        weights1[29120] <= 16'b1111111111111110;
        weights1[29121] <= 16'b1111111111111011;
        weights1[29122] <= 16'b1111111111111110;
        weights1[29123] <= 16'b1111111111111110;
        weights1[29124] <= 16'b0000000000000011;
        weights1[29125] <= 16'b0000000000000001;
        weights1[29126] <= 16'b0000000000000101;
        weights1[29127] <= 16'b1111111111111011;
        weights1[29128] <= 16'b0000000000000100;
        weights1[29129] <= 16'b1111111111111110;
        weights1[29130] <= 16'b1111111111111101;
        weights1[29131] <= 16'b1111111111111101;
        weights1[29132] <= 16'b0000000000000100;
        weights1[29133] <= 16'b0000000000000011;
        weights1[29134] <= 16'b0000000000001000;
        weights1[29135] <= 16'b0000000000000110;
        weights1[29136] <= 16'b0000000000001011;
        weights1[29137] <= 16'b1111111111101101;
        weights1[29138] <= 16'b0000000000000010;
        weights1[29139] <= 16'b0000000000000000;
        weights1[29140] <= 16'b0000000000001110;
        weights1[29141] <= 16'b0000000000000011;
        weights1[29142] <= 16'b1111111111110011;
        weights1[29143] <= 16'b1111111111111101;
        weights1[29144] <= 16'b1111111111110110;
        weights1[29145] <= 16'b1111111111111110;
        weights1[29146] <= 16'b1111111111111100;
        weights1[29147] <= 16'b1111111111110100;
        weights1[29148] <= 16'b0000000000000010;
        weights1[29149] <= 16'b0000000000000000;
        weights1[29150] <= 16'b1111111111111101;
        weights1[29151] <= 16'b1111111111110101;
        weights1[29152] <= 16'b1111111111111001;
        weights1[29153] <= 16'b0000000000000000;
        weights1[29154] <= 16'b0000000000000000;
        weights1[29155] <= 16'b1111111111110011;
        weights1[29156] <= 16'b1111111111111010;
        weights1[29157] <= 16'b1111111111111110;
        weights1[29158] <= 16'b1111111111111100;
        weights1[29159] <= 16'b1111111111111111;
        weights1[29160] <= 16'b1111111111110000;
        weights1[29161] <= 16'b1111111111110010;
        weights1[29162] <= 16'b0000000000001011;
        weights1[29163] <= 16'b0000000000000100;
        weights1[29164] <= 16'b1111111111111111;
        weights1[29165] <= 16'b1111111111111010;
        weights1[29166] <= 16'b1111111111110110;
        weights1[29167] <= 16'b0000000000001001;
        weights1[29168] <= 16'b1111111111110100;
        weights1[29169] <= 16'b0000000000011010;
        weights1[29170] <= 16'b0000000000000001;
        weights1[29171] <= 16'b0000000000001011;
        weights1[29172] <= 16'b0000000000000100;
        weights1[29173] <= 16'b0000000000000010;
        weights1[29174] <= 16'b1111111111111111;
        weights1[29175] <= 16'b0000000000000100;
        weights1[29176] <= 16'b0000000000000111;
        weights1[29177] <= 16'b0000000000000010;
        weights1[29178] <= 16'b0000000000001011;
        weights1[29179] <= 16'b0000000000000011;
        weights1[29180] <= 16'b0000000000000101;
        weights1[29181] <= 16'b1111111111111010;
        weights1[29182] <= 16'b1111111111110010;
        weights1[29183] <= 16'b1111111111111101;
        weights1[29184] <= 16'b1111111111111101;
        weights1[29185] <= 16'b1111111111111100;
        weights1[29186] <= 16'b0000000000000000;
        weights1[29187] <= 16'b1111111111111000;
        weights1[29188] <= 16'b0000000000000101;
        weights1[29189] <= 16'b1111111111110011;
        weights1[29190] <= 16'b1111111111101111;
        weights1[29191] <= 16'b1111111111111101;
        weights1[29192] <= 16'b1111111111111110;
        weights1[29193] <= 16'b0000000000000100;
        weights1[29194] <= 16'b1111111111111011;
        weights1[29195] <= 16'b1111111111110111;
        weights1[29196] <= 16'b1111111111111000;
        weights1[29197] <= 16'b0000000000001011;
        weights1[29198] <= 16'b0000000000000011;
        weights1[29199] <= 16'b1111111111111110;
        weights1[29200] <= 16'b1111111111101110;
        weights1[29201] <= 16'b1111111111111011;
        weights1[29202] <= 16'b1111111111111111;
        weights1[29203] <= 16'b0000000000000110;
        weights1[29204] <= 16'b0000000000001011;
        weights1[29205] <= 16'b0000000000010001;
        weights1[29206] <= 16'b0000000000001100;
        weights1[29207] <= 16'b0000000000000011;
        weights1[29208] <= 16'b0000000000000101;
        weights1[29209] <= 16'b1111111111110101;
        weights1[29210] <= 16'b0000000000001110;
        weights1[29211] <= 16'b1111111111111100;
        weights1[29212] <= 16'b1111111111111100;
        weights1[29213] <= 16'b0000000000000000;
        weights1[29214] <= 16'b1111111111101000;
        weights1[29215] <= 16'b0000000000000010;
        weights1[29216] <= 16'b0000000000000011;
        weights1[29217] <= 16'b0000000000000010;
        weights1[29218] <= 16'b0000000000010100;
        weights1[29219] <= 16'b1111111111110000;
        weights1[29220] <= 16'b0000000000000100;
        weights1[29221] <= 16'b0000000000000111;
        weights1[29222] <= 16'b0000000000000010;
        weights1[29223] <= 16'b0000000000000011;
        weights1[29224] <= 16'b0000000000000011;
        weights1[29225] <= 16'b1111111111111100;
        weights1[29226] <= 16'b0000000000000101;
        weights1[29227] <= 16'b0000000000000001;
        weights1[29228] <= 16'b1111111111111011;
        weights1[29229] <= 16'b0000000000000001;
        weights1[29230] <= 16'b0000000000001001;
        weights1[29231] <= 16'b0000000000001001;
        weights1[29232] <= 16'b0000000000001100;
        weights1[29233] <= 16'b0000000000010110;
        weights1[29234] <= 16'b0000000000000000;
        weights1[29235] <= 16'b0000000000010001;
        weights1[29236] <= 16'b1111111111111010;
        weights1[29237] <= 16'b1111111111111110;
        weights1[29238] <= 16'b0000000000000000;
        weights1[29239] <= 16'b0000000000000001;
        weights1[29240] <= 16'b1111111111110101;
        weights1[29241] <= 16'b1111111111110111;
        weights1[29242] <= 16'b1111111111111101;
        weights1[29243] <= 16'b1111111111110011;
        weights1[29244] <= 16'b0000000000001000;
        weights1[29245] <= 16'b1111111111111001;
        weights1[29246] <= 16'b1111111111111010;
        weights1[29247] <= 16'b1111111111111100;
        weights1[29248] <= 16'b0000000000000000;
        weights1[29249] <= 16'b1111111111111001;
        weights1[29250] <= 16'b0000000000001101;
        weights1[29251] <= 16'b0000000000001111;
        weights1[29252] <= 16'b0000000000001000;
        weights1[29253] <= 16'b1111111111110111;
        weights1[29254] <= 16'b1111111111111000;
        weights1[29255] <= 16'b1111111111111110;
        weights1[29256] <= 16'b0000000000000101;
        weights1[29257] <= 16'b0000000000010001;
        weights1[29258] <= 16'b1111111111101111;
        weights1[29259] <= 16'b1111111111110111;
        weights1[29260] <= 16'b0000000000001110;
        weights1[29261] <= 16'b0000000000001101;
        weights1[29262] <= 16'b1111111111111000;
        weights1[29263] <= 16'b0000000000000000;
        weights1[29264] <= 16'b1111111111111010;
        weights1[29265] <= 16'b1111111111111011;
        weights1[29266] <= 16'b0000000000000100;
        weights1[29267] <= 16'b0000000000000010;
        weights1[29268] <= 16'b0000000000001100;
        weights1[29269] <= 16'b0000000000001000;
        weights1[29270] <= 16'b1111111111110000;
        weights1[29271] <= 16'b1111111111111001;
        weights1[29272] <= 16'b1111111111110101;
        weights1[29273] <= 16'b1111111111111000;
        weights1[29274] <= 16'b0000000000001111;
        weights1[29275] <= 16'b1111111111111010;
        weights1[29276] <= 16'b1111111111111000;
        weights1[29277] <= 16'b0000000000001011;
        weights1[29278] <= 16'b1111111111111010;
        weights1[29279] <= 16'b0000000000000000;
        weights1[29280] <= 16'b1111111111110110;
        weights1[29281] <= 16'b0000000000001001;
        weights1[29282] <= 16'b0000000000001010;
        weights1[29283] <= 16'b1111111111111110;
        weights1[29284] <= 16'b1111111111111110;
        weights1[29285] <= 16'b1111111111111001;
        weights1[29286] <= 16'b0000000000000100;
        weights1[29287] <= 16'b0000000000000000;
        weights1[29288] <= 16'b0000000000000110;
        weights1[29289] <= 16'b1111111111111100;
        weights1[29290] <= 16'b1111111111110011;
        weights1[29291] <= 16'b0000000000000011;
        weights1[29292] <= 16'b1111111111111000;
        weights1[29293] <= 16'b1111111111111001;
        weights1[29294] <= 16'b1111111111110001;
        weights1[29295] <= 16'b0000000000000000;
        weights1[29296] <= 16'b1111111111111000;
        weights1[29297] <= 16'b1111111111111111;
        weights1[29298] <= 16'b0000000000001011;
        weights1[29299] <= 16'b1111111111110001;
        weights1[29300] <= 16'b0000000000001101;
        weights1[29301] <= 16'b1111111111101101;
        weights1[29302] <= 16'b1111111111110111;
        weights1[29303] <= 16'b1111111111111000;
        weights1[29304] <= 16'b1111111111111110;
        weights1[29305] <= 16'b1111111111111011;
        weights1[29306] <= 16'b0000000000000110;
        weights1[29307] <= 16'b0000000000000101;
        weights1[29308] <= 16'b0000000000000111;
        weights1[29309] <= 16'b0000000000000001;
        weights1[29310] <= 16'b1111111111110011;
        weights1[29311] <= 16'b0000000000001111;
        weights1[29312] <= 16'b1111111111111111;
        weights1[29313] <= 16'b0000000000010100;
        weights1[29314] <= 16'b1111111111110100;
        weights1[29315] <= 16'b1111111111111011;
        weights1[29316] <= 16'b0000000000000111;
        weights1[29317] <= 16'b0000000000000111;
        weights1[29318] <= 16'b1111111111111110;
        weights1[29319] <= 16'b0000000000010011;
        weights1[29320] <= 16'b0000000000011011;
        weights1[29321] <= 16'b1111111111111111;
        weights1[29322] <= 16'b0000000000001001;
        weights1[29323] <= 16'b0000000000000111;
        weights1[29324] <= 16'b0000000000000011;
        weights1[29325] <= 16'b0000000000000101;
        weights1[29326] <= 16'b0000000000001000;
        weights1[29327] <= 16'b1111111111110110;
        weights1[29328] <= 16'b0000000000000111;
        weights1[29329] <= 16'b1111111111111101;
        weights1[29330] <= 16'b0000000000000101;
        weights1[29331] <= 16'b1111111111111110;
        weights1[29332] <= 16'b1111111111111101;
        weights1[29333] <= 16'b0000000000000001;
        weights1[29334] <= 16'b0000000000000000;
        weights1[29335] <= 16'b0000000000000111;
        weights1[29336] <= 16'b1111111111111010;
        weights1[29337] <= 16'b0000000000000111;
        weights1[29338] <= 16'b0000000000001000;
        weights1[29339] <= 16'b1111111111111001;
        weights1[29340] <= 16'b0000000000000001;
        weights1[29341] <= 16'b1111111111110000;
        weights1[29342] <= 16'b1111111111111000;
        weights1[29343] <= 16'b0000000000000100;
        weights1[29344] <= 16'b0000000000001000;
        weights1[29345] <= 16'b1111111111110111;
        weights1[29346] <= 16'b0000000000000010;
        weights1[29347] <= 16'b0000000000001100;
        weights1[29348] <= 16'b1111111111111101;
        weights1[29349] <= 16'b0000000000001011;
        weights1[29350] <= 16'b0000000000000101;
        weights1[29351] <= 16'b0000000000001011;
        weights1[29352] <= 16'b0000000000001011;
        weights1[29353] <= 16'b1111111111111011;
        weights1[29354] <= 16'b1111111111110101;
        weights1[29355] <= 16'b0000000000001010;
        weights1[29356] <= 16'b1111111111110101;
        weights1[29357] <= 16'b0000000000000111;
        weights1[29358] <= 16'b1111111111110000;
        weights1[29359] <= 16'b0000000000000100;
        weights1[29360] <= 16'b1111111111111111;
        weights1[29361] <= 16'b0000000000000110;
        weights1[29362] <= 16'b0000000000000000;
        weights1[29363] <= 16'b1111111111110110;
        weights1[29364] <= 16'b0000000000001110;
        weights1[29365] <= 16'b0000000000000110;
        weights1[29366] <= 16'b0000000000000000;
        weights1[29367] <= 16'b0000000000000011;
        weights1[29368] <= 16'b1111111111101110;
        weights1[29369] <= 16'b1111111111111100;
        weights1[29370] <= 16'b1111111111110110;
        weights1[29371] <= 16'b1111111111111110;
        weights1[29372] <= 16'b1111111111111101;
        weights1[29373] <= 16'b1111111111111000;
        weights1[29374] <= 16'b0000000000001010;
        weights1[29375] <= 16'b0000000000000011;
        weights1[29376] <= 16'b1111111111110101;
        weights1[29377] <= 16'b1111111111111001;
        weights1[29378] <= 16'b0000000000000011;
        weights1[29379] <= 16'b0000000000000000;
        weights1[29380] <= 16'b1111111111110111;
        weights1[29381] <= 16'b0000000000001101;
        weights1[29382] <= 16'b0000000000001001;
        weights1[29383] <= 16'b0000000000001001;
        weights1[29384] <= 16'b1111111111110010;
        weights1[29385] <= 16'b1111111111111010;
        weights1[29386] <= 16'b0000000000000011;
        weights1[29387] <= 16'b1111111111101101;
        weights1[29388] <= 16'b1111111111111110;
        weights1[29389] <= 16'b0000000000000100;
        weights1[29390] <= 16'b1111111111111111;
        weights1[29391] <= 16'b0000000000000110;
        weights1[29392] <= 16'b0000000000010010;
        weights1[29393] <= 16'b1111111111111001;
        weights1[29394] <= 16'b1111111111111010;
        weights1[29395] <= 16'b1111111111110100;
        weights1[29396] <= 16'b0000000000001001;
        weights1[29397] <= 16'b1111111111111000;
        weights1[29398] <= 16'b0000000000000100;
        weights1[29399] <= 16'b1111111111111100;
        weights1[29400] <= 16'b1111111111110100;
        weights1[29401] <= 16'b1111111111101111;
        weights1[29402] <= 16'b1111111111111110;
        weights1[29403] <= 16'b1111111111101110;
        weights1[29404] <= 16'b1111111111110101;
        weights1[29405] <= 16'b0000000000001000;
        weights1[29406] <= 16'b1111111111111000;
        weights1[29407] <= 16'b0000000000001000;
        weights1[29408] <= 16'b0000000000001000;
        weights1[29409] <= 16'b1111111111111110;
        weights1[29410] <= 16'b1111111111111100;
        weights1[29411] <= 16'b0000000000000010;
        weights1[29412] <= 16'b0000000000001011;
        weights1[29413] <= 16'b0000000000000000;
        weights1[29414] <= 16'b0000000000000001;
        weights1[29415] <= 16'b1111111111110100;
        weights1[29416] <= 16'b0000000000000011;
        weights1[29417] <= 16'b1111111111111010;
        weights1[29418] <= 16'b0000000000010001;
        weights1[29419] <= 16'b0000000000000001;
        weights1[29420] <= 16'b0000000000001000;
        weights1[29421] <= 16'b1111111111111110;
        weights1[29422] <= 16'b0000000000001100;
        weights1[29423] <= 16'b0000000000001000;
        weights1[29424] <= 16'b1111111111111011;
        weights1[29425] <= 16'b0000000000000001;
        weights1[29426] <= 16'b0000000000000110;
        weights1[29427] <= 16'b0000000000000110;
        weights1[29428] <= 16'b1111111111110011;
        weights1[29429] <= 16'b1111111111110101;
        weights1[29430] <= 16'b1111111111111000;
        weights1[29431] <= 16'b1111111111110110;
        weights1[29432] <= 16'b0000000000000101;
        weights1[29433] <= 16'b0000000000001010;
        weights1[29434] <= 16'b0000000000000011;
        weights1[29435] <= 16'b0000000000011001;
        weights1[29436] <= 16'b0000000000001011;
        weights1[29437] <= 16'b0000000000001110;
        weights1[29438] <= 16'b1111111111101110;
        weights1[29439] <= 16'b0000000000001010;
        weights1[29440] <= 16'b1111111111110100;
        weights1[29441] <= 16'b1111111111111001;
        weights1[29442] <= 16'b0000000000000011;
        weights1[29443] <= 16'b0000000000000010;
        weights1[29444] <= 16'b1111111111110000;
        weights1[29445] <= 16'b0000000000000000;
        weights1[29446] <= 16'b0000000000000010;
        weights1[29447] <= 16'b0000000000000111;
        weights1[29448] <= 16'b0000000000010000;
        weights1[29449] <= 16'b0000000000000100;
        weights1[29450] <= 16'b0000000000001001;
        weights1[29451] <= 16'b1111111111110001;
        weights1[29452] <= 16'b1111111111111110;
        weights1[29453] <= 16'b0000000000001000;
        weights1[29454] <= 16'b0000000000000000;
        weights1[29455] <= 16'b0000000000000101;
        weights1[29456] <= 16'b1111111111110011;
        weights1[29457] <= 16'b1111111111110110;
        weights1[29458] <= 16'b0000000000000000;
        weights1[29459] <= 16'b1111111111110100;
        weights1[29460] <= 16'b1111111111111111;
        weights1[29461] <= 16'b0000000000011000;
        weights1[29462] <= 16'b0000000000010110;
        weights1[29463] <= 16'b0000000000000110;
        weights1[29464] <= 16'b0000000000001100;
        weights1[29465] <= 16'b1111111111110111;
        weights1[29466] <= 16'b1111111111101001;
        weights1[29467] <= 16'b1111111111110001;
        weights1[29468] <= 16'b0000000000000000;
        weights1[29469] <= 16'b1111111111111100;
        weights1[29470] <= 16'b1111111111101011;
        weights1[29471] <= 16'b1111111111100000;
        weights1[29472] <= 16'b1111111111110111;
        weights1[29473] <= 16'b1111111111110011;
        weights1[29474] <= 16'b0000000000011010;
        weights1[29475] <= 16'b0000000000011010;
        weights1[29476] <= 16'b0000000000001011;
        weights1[29477] <= 16'b0000000000001010;
        weights1[29478] <= 16'b0000000000001100;
        weights1[29479] <= 16'b1111111111111110;
        weights1[29480] <= 16'b1111111111101001;
        weights1[29481] <= 16'b1111111111111111;
        weights1[29482] <= 16'b0000000000000010;
        weights1[29483] <= 16'b1111111111111111;
        weights1[29484] <= 16'b1111111111111101;
        weights1[29485] <= 16'b0000000000000111;
        weights1[29486] <= 16'b0000000000001110;
        weights1[29487] <= 16'b0000000000000010;
        weights1[29488] <= 16'b0000000000000110;
        weights1[29489] <= 16'b0000000000011001;
        weights1[29490] <= 16'b0000000000001011;
        weights1[29491] <= 16'b1111111111111011;
        weights1[29492] <= 16'b1111111111111001;
        weights1[29493] <= 16'b1111111111011100;
        weights1[29494] <= 16'b1111111111101110;
        weights1[29495] <= 16'b0000000000000011;
        weights1[29496] <= 16'b0000000000010111;
        weights1[29497] <= 16'b0000000000001001;
        weights1[29498] <= 16'b1111111111111111;
        weights1[29499] <= 16'b1111111111101111;
        weights1[29500] <= 16'b1111111111011011;
        weights1[29501] <= 16'b1111111111100101;
        weights1[29502] <= 16'b0000000000000010;
        weights1[29503] <= 16'b0000000000010011;
        weights1[29504] <= 16'b0000000000010000;
        weights1[29505] <= 16'b0000000000001110;
        weights1[29506] <= 16'b1111111111111000;
        weights1[29507] <= 16'b1111111111101011;
        weights1[29508] <= 16'b1111111111101001;
        weights1[29509] <= 16'b1111111111011011;
        weights1[29510] <= 16'b1111111111110010;
        weights1[29511] <= 16'b1111111111111100;
        weights1[29512] <= 16'b0000000000001010;
        weights1[29513] <= 16'b0000000000010000;
        weights1[29514] <= 16'b0000000000010100;
        weights1[29515] <= 16'b0000000000010010;
        weights1[29516] <= 16'b0000000000101011;
        weights1[29517] <= 16'b0000000000100111;
        weights1[29518] <= 16'b1111111111111101;
        weights1[29519] <= 16'b0000000000010101;
        weights1[29520] <= 16'b1111111111101110;
        weights1[29521] <= 16'b1111111111001101;
        weights1[29522] <= 16'b1111111111110111;
        weights1[29523] <= 16'b1111111111110101;
        weights1[29524] <= 16'b0000000000100111;
        weights1[29525] <= 16'b0000000000100000;
        weights1[29526] <= 16'b1111111111110101;
        weights1[29527] <= 16'b1111111111100110;
        weights1[29528] <= 16'b1111111111011010;
        weights1[29529] <= 16'b1111111111010111;
        weights1[29530] <= 16'b0000000000001110;
        weights1[29531] <= 16'b0000000000101100;
        weights1[29532] <= 16'b0000000000000110;
        weights1[29533] <= 16'b0000000000100110;
        weights1[29534] <= 16'b0000000000010000;
        weights1[29535] <= 16'b1111111111111111;
        weights1[29536] <= 16'b1111111111100001;
        weights1[29537] <= 16'b1111111111100111;
        weights1[29538] <= 16'b1111111111100101;
        weights1[29539] <= 16'b1111111111111100;
        weights1[29540] <= 16'b0000000000010001;
        weights1[29541] <= 16'b0000000000010010;
        weights1[29542] <= 16'b0000000000011110;
        weights1[29543] <= 16'b0000000000101001;
        weights1[29544] <= 16'b0000000000101110;
        weights1[29545] <= 16'b0000000000100101;
        weights1[29546] <= 16'b1111111111111001;
        weights1[29547] <= 16'b1111111111011000;
        weights1[29548] <= 16'b1111111111011100;
        weights1[29549] <= 16'b1111111111011011;
        weights1[29550] <= 16'b1111111111110110;
        weights1[29551] <= 16'b0000000000001111;
        weights1[29552] <= 16'b0000000000100001;
        weights1[29553] <= 16'b0000000000011100;
        weights1[29554] <= 16'b1111111111110100;
        weights1[29555] <= 16'b1111111111011011;
        weights1[29556] <= 16'b1111111110111111;
        weights1[29557] <= 16'b1111111111001010;
        weights1[29558] <= 16'b0000000000001101;
        weights1[29559] <= 16'b0000000000100101;
        weights1[29560] <= 16'b0000000000000111;
        weights1[29561] <= 16'b0000000000101100;
        weights1[29562] <= 16'b0000000000001101;
        weights1[29563] <= 16'b0000000000001001;
        weights1[29564] <= 16'b0000000000000111;
        weights1[29565] <= 16'b1111111111010110;
        weights1[29566] <= 16'b1111111111100111;
        weights1[29567] <= 16'b1111111111110001;
        weights1[29568] <= 16'b0000000000001100;
        weights1[29569] <= 16'b0000000000011001;
        weights1[29570] <= 16'b0000000000100000;
        weights1[29571] <= 16'b0000000000011100;
        weights1[29572] <= 16'b0000000000010010;
        weights1[29573] <= 16'b0000000000000000;
        weights1[29574] <= 16'b1111111111101110;
        weights1[29575] <= 16'b1111111111001100;
        weights1[29576] <= 16'b1111111110110111;
        weights1[29577] <= 16'b1111111111010001;
        weights1[29578] <= 16'b1111111111101000;
        weights1[29579] <= 16'b0000000000100000;
        weights1[29580] <= 16'b0000000000111111;
        weights1[29581] <= 16'b0000000000001000;
        weights1[29582] <= 16'b1111111111111000;
        weights1[29583] <= 16'b1111111111000111;
        weights1[29584] <= 16'b1111111111000110;
        weights1[29585] <= 16'b1111111110110100;
        weights1[29586] <= 16'b0000000000001010;
        weights1[29587] <= 16'b0000000001000100;
        weights1[29588] <= 16'b0000000000010011;
        weights1[29589] <= 16'b0000000000010000;
        weights1[29590] <= 16'b0000000000100100;
        weights1[29591] <= 16'b0000000000010000;
        weights1[29592] <= 16'b1111111111111111;
        weights1[29593] <= 16'b1111111111011010;
        weights1[29594] <= 16'b1111111111101100;
        weights1[29595] <= 16'b1111111111101110;
        weights1[29596] <= 16'b0000000000000111;
        weights1[29597] <= 16'b0000000000001100;
        weights1[29598] <= 16'b0000000000011000;
        weights1[29599] <= 16'b0000000000000010;
        weights1[29600] <= 16'b0000000000000000;
        weights1[29601] <= 16'b1111111111011011;
        weights1[29602] <= 16'b1111111111001100;
        weights1[29603] <= 16'b1111111110011001;
        weights1[29604] <= 16'b1111111110010110;
        weights1[29605] <= 16'b1111111111111101;
        weights1[29606] <= 16'b0000000000011101;
        weights1[29607] <= 16'b0000000000110100;
        weights1[29608] <= 16'b0000000001010100;
        weights1[29609] <= 16'b0000000000000000;
        weights1[29610] <= 16'b1111111111011110;
        weights1[29611] <= 16'b1111111111010000;
        weights1[29612] <= 16'b1111111110000110;
        weights1[29613] <= 16'b1111111110010111;
        weights1[29614] <= 16'b0000000000101101;
        weights1[29615] <= 16'b0000000001001110;
        weights1[29616] <= 16'b0000000000011110;
        weights1[29617] <= 16'b0000000000001110;
        weights1[29618] <= 16'b0000000000010111;
        weights1[29619] <= 16'b0000000000001001;
        weights1[29620] <= 16'b0000000000011001;
        weights1[29621] <= 16'b1111111111011111;
        weights1[29622] <= 16'b1111111111111001;
        weights1[29623] <= 16'b1111111111101110;
        weights1[29624] <= 16'b1111111111111110;
        weights1[29625] <= 16'b1111111111111111;
        weights1[29626] <= 16'b1111111111111011;
        weights1[29627] <= 16'b1111111111010111;
        weights1[29628] <= 16'b1111111110111110;
        weights1[29629] <= 16'b1111111110110000;
        weights1[29630] <= 16'b1111111110000010;
        weights1[29631] <= 16'b1111111101011101;
        weights1[29632] <= 16'b1111111111011100;
        weights1[29633] <= 16'b1111111111111110;
        weights1[29634] <= 16'b0000000000110100;
        weights1[29635] <= 16'b0000000000110100;
        weights1[29636] <= 16'b0000000000111111;
        weights1[29637] <= 16'b1111111111110110;
        weights1[29638] <= 16'b1111111111001011;
        weights1[29639] <= 16'b1111111110110000;
        weights1[29640] <= 16'b1111111101001010;
        weights1[29641] <= 16'b1111111101110110;
        weights1[29642] <= 16'b0000000000100100;
        weights1[29643] <= 16'b0000000001100100;
        weights1[29644] <= 16'b0000000000010111;
        weights1[29645] <= 16'b0000000000100111;
        weights1[29646] <= 16'b0000000000100011;
        weights1[29647] <= 16'b0000000000001110;
        weights1[29648] <= 16'b1111111111110110;
        weights1[29649] <= 16'b1111111111111001;
        weights1[29650] <= 16'b1111111111101101;
        weights1[29651] <= 16'b1111111111111001;
        weights1[29652] <= 16'b1111111111111000;
        weights1[29653] <= 16'b1111111111101010;
        weights1[29654] <= 16'b1111111111011100;
        weights1[29655] <= 16'b1111111111001011;
        weights1[29656] <= 16'b1111111110111000;
        weights1[29657] <= 16'b1111111110010101;
        weights1[29658] <= 16'b1111111101110110;
        weights1[29659] <= 16'b1111111110100101;
        weights1[29660] <= 16'b0000000000000000;
        weights1[29661] <= 16'b0000000000011101;
        weights1[29662] <= 16'b0000000000100101;
        weights1[29663] <= 16'b0000000000111001;
        weights1[29664] <= 16'b0000000000110111;
        weights1[29665] <= 16'b0000000000001101;
        weights1[29666] <= 16'b1111111110110010;
        weights1[29667] <= 16'b1111111101111011;
        weights1[29668] <= 16'b1111111101001101;
        weights1[29669] <= 16'b1111111110100100;
        weights1[29670] <= 16'b0000000001000111;
        weights1[29671] <= 16'b0000000001000111;
        weights1[29672] <= 16'b0000000000011110;
        weights1[29673] <= 16'b0000000000101111;
        weights1[29674] <= 16'b0000000000001010;
        weights1[29675] <= 16'b0000000000000110;
        weights1[29676] <= 16'b0000000000010001;
        weights1[29677] <= 16'b0000000000000011;
        weights1[29678] <= 16'b1111111111110110;
        weights1[29679] <= 16'b1111111111111100;
        weights1[29680] <= 16'b1111111111110101;
        weights1[29681] <= 16'b1111111111100111;
        weights1[29682] <= 16'b1111111111011001;
        weights1[29683] <= 16'b1111111111000011;
        weights1[29684] <= 16'b1111111110101100;
        weights1[29685] <= 16'b1111111110000110;
        weights1[29686] <= 16'b1111111110100110;
        weights1[29687] <= 16'b1111111111101100;
        weights1[29688] <= 16'b0000000001000111;
        weights1[29689] <= 16'b0000000000101010;
        weights1[29690] <= 16'b0000000000010010;
        weights1[29691] <= 16'b0000000000100011;
        weights1[29692] <= 16'b0000000000100101;
        weights1[29693] <= 16'b1111111110110010;
        weights1[29694] <= 16'b1111111110100100;
        weights1[29695] <= 16'b1111111101100101;
        weights1[29696] <= 16'b1111111101010001;
        weights1[29697] <= 16'b1111111110101011;
        weights1[29698] <= 16'b0000000000010110;
        weights1[29699] <= 16'b0000000000111001;
        weights1[29700] <= 16'b0000000000011100;
        weights1[29701] <= 16'b1111111111111010;
        weights1[29702] <= 16'b0000000000011101;
        weights1[29703] <= 16'b0000000000101011;
        weights1[29704] <= 16'b0000000000011101;
        weights1[29705] <= 16'b0000000000000110;
        weights1[29706] <= 16'b1111111111111100;
        weights1[29707] <= 16'b1111111111111010;
        weights1[29708] <= 16'b1111111111111100;
        weights1[29709] <= 16'b1111111111101101;
        weights1[29710] <= 16'b1111111111100010;
        weights1[29711] <= 16'b1111111111000001;
        weights1[29712] <= 16'b1111111110100011;
        weights1[29713] <= 16'b1111111110100011;
        weights1[29714] <= 16'b1111111111011001;
        weights1[29715] <= 16'b1111111111111101;
        weights1[29716] <= 16'b0000000000111100;
        weights1[29717] <= 16'b0000000001000111;
        weights1[29718] <= 16'b0000000000101011;
        weights1[29719] <= 16'b0000000000111111;
        weights1[29720] <= 16'b0000000000011101;
        weights1[29721] <= 16'b1111111111000000;
        weights1[29722] <= 16'b1111111110010001;
        weights1[29723] <= 16'b1111111101010100;
        weights1[29724] <= 16'b1111111100101110;
        weights1[29725] <= 16'b1111111110111011;
        weights1[29726] <= 16'b0000000000000000;
        weights1[29727] <= 16'b0000000000111111;
        weights1[29728] <= 16'b0000000000101100;
        weights1[29729] <= 16'b0000000000011000;
        weights1[29730] <= 16'b0000000000011001;
        weights1[29731] <= 16'b0000000000100101;
        weights1[29732] <= 16'b0000000000011000;
        weights1[29733] <= 16'b0000000000001000;
        weights1[29734] <= 16'b1111111111111011;
        weights1[29735] <= 16'b1111111111111011;
        weights1[29736] <= 16'b1111111111111011;
        weights1[29737] <= 16'b1111111111110001;
        weights1[29738] <= 16'b1111111111100001;
        weights1[29739] <= 16'b1111111111001101;
        weights1[29740] <= 16'b1111111111001000;
        weights1[29741] <= 16'b1111111111001110;
        weights1[29742] <= 16'b1111111111111001;
        weights1[29743] <= 16'b0000000000100101;
        weights1[29744] <= 16'b0000000000011100;
        weights1[29745] <= 16'b0000000000001111;
        weights1[29746] <= 16'b0000000000011110;
        weights1[29747] <= 16'b0000000000010011;
        weights1[29748] <= 16'b1111111111100111;
        weights1[29749] <= 16'b1111111111010010;
        weights1[29750] <= 16'b1111111110000101;
        weights1[29751] <= 16'b1111111101101011;
        weights1[29752] <= 16'b1111111101110001;
        weights1[29753] <= 16'b1111111111000110;
        weights1[29754] <= 16'b1111111111111010;
        weights1[29755] <= 16'b0000000000001100;
        weights1[29756] <= 16'b0000000000010010;
        weights1[29757] <= 16'b0000000000001110;
        weights1[29758] <= 16'b0000000000011010;
        weights1[29759] <= 16'b0000000000100011;
        weights1[29760] <= 16'b0000000000010110;
        weights1[29761] <= 16'b0000000000001111;
        weights1[29762] <= 16'b0000000000000111;
        weights1[29763] <= 16'b0000000000000000;
        weights1[29764] <= 16'b1111111111111110;
        weights1[29765] <= 16'b1111111111110110;
        weights1[29766] <= 16'b1111111111101011;
        weights1[29767] <= 16'b1111111111100101;
        weights1[29768] <= 16'b1111111111110000;
        weights1[29769] <= 16'b1111111111111001;
        weights1[29770] <= 16'b0000000000100000;
        weights1[29771] <= 16'b0000000000101100;
        weights1[29772] <= 16'b0000000000101000;
        weights1[29773] <= 16'b0000000000101010;
        weights1[29774] <= 16'b1111111111111011;
        weights1[29775] <= 16'b1111111111110011;
        weights1[29776] <= 16'b1111111111010111;
        weights1[29777] <= 16'b1111111110100101;
        weights1[29778] <= 16'b1111111101101100;
        weights1[29779] <= 16'b1111111101001101;
        weights1[29780] <= 16'b1111111101011101;
        weights1[29781] <= 16'b1111111110100001;
        weights1[29782] <= 16'b1111111111010011;
        weights1[29783] <= 16'b1111111111101110;
        weights1[29784] <= 16'b0000000000001100;
        weights1[29785] <= 16'b0000000000011011;
        weights1[29786] <= 16'b0000000000011110;
        weights1[29787] <= 16'b0000000000100100;
        weights1[29788] <= 16'b0000000000100111;
        weights1[29789] <= 16'b0000000000001101;
        weights1[29790] <= 16'b0000000000001001;
        weights1[29791] <= 16'b0000000000000011;
        weights1[29792] <= 16'b0000000000000000;
        weights1[29793] <= 16'b0000000000000000;
        weights1[29794] <= 16'b0000000000000000;
        weights1[29795] <= 16'b0000000000000000;
        weights1[29796] <= 16'b1111111111111111;
        weights1[29797] <= 16'b1111111111111111;
        weights1[29798] <= 16'b0000000000000000;
        weights1[29799] <= 16'b1111111111111111;
        weights1[29800] <= 16'b0000000000000010;
        weights1[29801] <= 16'b0000000000000001;
        weights1[29802] <= 16'b1111111111111111;
        weights1[29803] <= 16'b0000000000000100;
        weights1[29804] <= 16'b0000000000001100;
        weights1[29805] <= 16'b0000000000001010;
        weights1[29806] <= 16'b0000000000010110;
        weights1[29807] <= 16'b0000000000011011;
        weights1[29808] <= 16'b0000000000010111;
        weights1[29809] <= 16'b0000000000001001;
        weights1[29810] <= 16'b0000000000001000;
        weights1[29811] <= 16'b0000000000001100;
        weights1[29812] <= 16'b0000000000001001;
        weights1[29813] <= 16'b1111111111111110;
        weights1[29814] <= 16'b1111111111111010;
        weights1[29815] <= 16'b1111111111111111;
        weights1[29816] <= 16'b1111111111111101;
        weights1[29817] <= 16'b1111111111111111;
        weights1[29818] <= 16'b1111111111111111;
        weights1[29819] <= 16'b0000000000000000;
        weights1[29820] <= 16'b0000000000000000;
        weights1[29821] <= 16'b0000000000000000;
        weights1[29822] <= 16'b0000000000000000;
        weights1[29823] <= 16'b1111111111111110;
        weights1[29824] <= 16'b1111111111111111;
        weights1[29825] <= 16'b1111111111111100;
        weights1[29826] <= 16'b0000000000000000;
        weights1[29827] <= 16'b1111111111111110;
        weights1[29828] <= 16'b1111111111111110;
        weights1[29829] <= 16'b1111111111111100;
        weights1[29830] <= 16'b0000000000000000;
        weights1[29831] <= 16'b0000000000001000;
        weights1[29832] <= 16'b0000000000001100;
        weights1[29833] <= 16'b0000000000001111;
        weights1[29834] <= 16'b0000000000001011;
        weights1[29835] <= 16'b0000000000011000;
        weights1[29836] <= 16'b0000000000010010;
        weights1[29837] <= 16'b0000000000001010;
        weights1[29838] <= 16'b0000000000001000;
        weights1[29839] <= 16'b0000000000000101;
        weights1[29840] <= 16'b0000000000001001;
        weights1[29841] <= 16'b0000000000000100;
        weights1[29842] <= 16'b0000000000000011;
        weights1[29843] <= 16'b1111111111111110;
        weights1[29844] <= 16'b1111111111111010;
        weights1[29845] <= 16'b1111111111111100;
        weights1[29846] <= 16'b1111111111111111;
        weights1[29847] <= 16'b0000000000000000;
        weights1[29848] <= 16'b0000000000000000;
        weights1[29849] <= 16'b0000000000000000;
        weights1[29850] <= 16'b1111111111111110;
        weights1[29851] <= 16'b1111111111111011;
        weights1[29852] <= 16'b1111111111111101;
        weights1[29853] <= 16'b1111111111111101;
        weights1[29854] <= 16'b1111111111111100;
        weights1[29855] <= 16'b1111111111111101;
        weights1[29856] <= 16'b1111111111111001;
        weights1[29857] <= 16'b1111111111110101;
        weights1[29858] <= 16'b1111111111110110;
        weights1[29859] <= 16'b0000000000000000;
        weights1[29860] <= 16'b0000000000000111;
        weights1[29861] <= 16'b0000000000010100;
        weights1[29862] <= 16'b0000000000011000;
        weights1[29863] <= 16'b0000000000011100;
        weights1[29864] <= 16'b0000000000010000;
        weights1[29865] <= 16'b0000000000001010;
        weights1[29866] <= 16'b0000000000001011;
        weights1[29867] <= 16'b0000000000000100;
        weights1[29868] <= 16'b0000000000000000;
        weights1[29869] <= 16'b1111111111111010;
        weights1[29870] <= 16'b1111111111101110;
        weights1[29871] <= 16'b1111111111101110;
        weights1[29872] <= 16'b1111111111110010;
        weights1[29873] <= 16'b1111111111111011;
        weights1[29874] <= 16'b1111111111111110;
        weights1[29875] <= 16'b1111111111111111;
        weights1[29876] <= 16'b0000000000000000;
        weights1[29877] <= 16'b0000000000000000;
        weights1[29878] <= 16'b1111111111111101;
        weights1[29879] <= 16'b1111111111111101;
        weights1[29880] <= 16'b1111111111111010;
        weights1[29881] <= 16'b1111111111111101;
        weights1[29882] <= 16'b1111111111110110;
        weights1[29883] <= 16'b1111111111110100;
        weights1[29884] <= 16'b1111111111110100;
        weights1[29885] <= 16'b1111111111101101;
        weights1[29886] <= 16'b1111111111101010;
        weights1[29887] <= 16'b1111111111111000;
        weights1[29888] <= 16'b1111111111111111;
        weights1[29889] <= 16'b0000000000001011;
        weights1[29890] <= 16'b0000000000001011;
        weights1[29891] <= 16'b0000000000001101;
        weights1[29892] <= 16'b0000000000001001;
        weights1[29893] <= 16'b0000000000000011;
        weights1[29894] <= 16'b0000000000000011;
        weights1[29895] <= 16'b1111111111111100;
        weights1[29896] <= 16'b1111111111111101;
        weights1[29897] <= 16'b1111111111111100;
        weights1[29898] <= 16'b1111111111100111;
        weights1[29899] <= 16'b1111111111100110;
        weights1[29900] <= 16'b1111111111101111;
        weights1[29901] <= 16'b1111111111110101;
        weights1[29902] <= 16'b1111111111111010;
        weights1[29903] <= 16'b1111111111111111;
        weights1[29904] <= 16'b0000000000000000;
        weights1[29905] <= 16'b0000000000000001;
        weights1[29906] <= 16'b1111111111111110;
        weights1[29907] <= 16'b1111111111111000;
        weights1[29908] <= 16'b1111111111111011;
        weights1[29909] <= 16'b1111111111111000;
        weights1[29910] <= 16'b1111111111101110;
        weights1[29911] <= 16'b1111111111101001;
        weights1[29912] <= 16'b1111111111101010;
        weights1[29913] <= 16'b1111111111100111;
        weights1[29914] <= 16'b1111111111101011;
        weights1[29915] <= 16'b1111111111110100;
        weights1[29916] <= 16'b1111111111111101;
        weights1[29917] <= 16'b1111111111111100;
        weights1[29918] <= 16'b0000000000001000;
        weights1[29919] <= 16'b1111111111111111;
        weights1[29920] <= 16'b1111111111110111;
        weights1[29921] <= 16'b0000000000000100;
        weights1[29922] <= 16'b1111111111111010;
        weights1[29923] <= 16'b1111111111110100;
        weights1[29924] <= 16'b1111111111101101;
        weights1[29925] <= 16'b1111111111101001;
        weights1[29926] <= 16'b1111111111101011;
        weights1[29927] <= 16'b1111111111101001;
        weights1[29928] <= 16'b1111111111101100;
        weights1[29929] <= 16'b1111111111110111;
        weights1[29930] <= 16'b1111111111111001;
        weights1[29931] <= 16'b1111111111111110;
        weights1[29932] <= 16'b0000000000000001;
        weights1[29933] <= 16'b0000000000000010;
        weights1[29934] <= 16'b1111111111111101;
        weights1[29935] <= 16'b1111111111111100;
        weights1[29936] <= 16'b1111111111110110;
        weights1[29937] <= 16'b1111111111111100;
        weights1[29938] <= 16'b1111111111111000;
        weights1[29939] <= 16'b1111111111110111;
        weights1[29940] <= 16'b1111111111101100;
        weights1[29941] <= 16'b1111111111100110;
        weights1[29942] <= 16'b1111111111101000;
        weights1[29943] <= 16'b1111111111110100;
        weights1[29944] <= 16'b1111111111110011;
        weights1[29945] <= 16'b0000000000000001;
        weights1[29946] <= 16'b1111111111111100;
        weights1[29947] <= 16'b0000000000000111;
        weights1[29948] <= 16'b0000000000000101;
        weights1[29949] <= 16'b0000000000001011;
        weights1[29950] <= 16'b0000000000000001;
        weights1[29951] <= 16'b1111111111110101;
        weights1[29952] <= 16'b1111111111110101;
        weights1[29953] <= 16'b1111111111101100;
        weights1[29954] <= 16'b1111111111011001;
        weights1[29955] <= 16'b1111111111100011;
        weights1[29956] <= 16'b1111111111110010;
        weights1[29957] <= 16'b1111111111110101;
        weights1[29958] <= 16'b1111111111111100;
        weights1[29959] <= 16'b0000000000000000;
        weights1[29960] <= 16'b0000000000000000;
        weights1[29961] <= 16'b0000000000000000;
        weights1[29962] <= 16'b0000000000000001;
        weights1[29963] <= 16'b1111111111111101;
        weights1[29964] <= 16'b1111111111111001;
        weights1[29965] <= 16'b1111111111111101;
        weights1[29966] <= 16'b1111111111110100;
        weights1[29967] <= 16'b1111111111110000;
        weights1[29968] <= 16'b1111111111101101;
        weights1[29969] <= 16'b1111111111101110;
        weights1[29970] <= 16'b1111111111101010;
        weights1[29971] <= 16'b1111111111100111;
        weights1[29972] <= 16'b1111111111101111;
        weights1[29973] <= 16'b1111111111110100;
        weights1[29974] <= 16'b1111111111111111;
        weights1[29975] <= 16'b0000000000001011;
        weights1[29976] <= 16'b0000000000010110;
        weights1[29977] <= 16'b0000000000000111;
        weights1[29978] <= 16'b1111111111111000;
        weights1[29979] <= 16'b1111111111110010;
        weights1[29980] <= 16'b1111111111101100;
        weights1[29981] <= 16'b1111111111100011;
        weights1[29982] <= 16'b1111111111011011;
        weights1[29983] <= 16'b1111111111101000;
        weights1[29984] <= 16'b1111111111101100;
        weights1[29985] <= 16'b1111111111110111;
        weights1[29986] <= 16'b1111111111111100;
        weights1[29987] <= 16'b1111111111111111;
        weights1[29988] <= 16'b0000000000000001;
        weights1[29989] <= 16'b0000000000000000;
        weights1[29990] <= 16'b0000000000000000;
        weights1[29991] <= 16'b1111111111111101;
        weights1[29992] <= 16'b0000000000000000;
        weights1[29993] <= 16'b1111111111111101;
        weights1[29994] <= 16'b1111111111110001;
        weights1[29995] <= 16'b1111111111110110;
        weights1[29996] <= 16'b1111111111101101;
        weights1[29997] <= 16'b1111111111100011;
        weights1[29998] <= 16'b1111111111100000;
        weights1[29999] <= 16'b1111111111011011;
        weights1[30000] <= 16'b1111111111011101;
        weights1[30001] <= 16'b1111111111100110;
        weights1[30002] <= 16'b1111111111100111;
        weights1[30003] <= 16'b1111111111111111;
        weights1[30004] <= 16'b0000000000001101;
        weights1[30005] <= 16'b0000000000001111;
        weights1[30006] <= 16'b1111111111111100;
        weights1[30007] <= 16'b1111111111101111;
        weights1[30008] <= 16'b1111111111100111;
        weights1[30009] <= 16'b1111111111011010;
        weights1[30010] <= 16'b1111111111010111;
        weights1[30011] <= 16'b1111111111100111;
        weights1[30012] <= 16'b1111111111101100;
        weights1[30013] <= 16'b1111111111111000;
        weights1[30014] <= 16'b1111111111111110;
        weights1[30015] <= 16'b1111111111111111;
        weights1[30016] <= 16'b0000000000000000;
        weights1[30017] <= 16'b0000000000000000;
        weights1[30018] <= 16'b0000000000000000;
        weights1[30019] <= 16'b0000000000000000;
        weights1[30020] <= 16'b0000000000000011;
        weights1[30021] <= 16'b0000000000000010;
        weights1[30022] <= 16'b1111111111111010;
        weights1[30023] <= 16'b1111111111111100;
        weights1[30024] <= 16'b1111111111101101;
        weights1[30025] <= 16'b1111111111100001;
        weights1[30026] <= 16'b1111111111011100;
        weights1[30027] <= 16'b1111111111011000;
        weights1[30028] <= 16'b1111111111100101;
        weights1[30029] <= 16'b1111111111101011;
        weights1[30030] <= 16'b1111111111110011;
        weights1[30031] <= 16'b0000000000000100;
        weights1[30032] <= 16'b0000000000010011;
        weights1[30033] <= 16'b0000000000010011;
        weights1[30034] <= 16'b0000000000000110;
        weights1[30035] <= 16'b0000000000000001;
        weights1[30036] <= 16'b1111111111101011;
        weights1[30037] <= 16'b1111111111101101;
        weights1[30038] <= 16'b1111111111011100;
        weights1[30039] <= 16'b1111111111100101;
        weights1[30040] <= 16'b1111111111101100;
        weights1[30041] <= 16'b1111111111110010;
        weights1[30042] <= 16'b1111111111111000;
        weights1[30043] <= 16'b1111111111111100;
        weights1[30044] <= 16'b1111111111111110;
        weights1[30045] <= 16'b0000000000000010;
        weights1[30046] <= 16'b0000000000001001;
        weights1[30047] <= 16'b0000000000000010;
        weights1[30048] <= 16'b0000000000000100;
        weights1[30049] <= 16'b0000000000000111;
        weights1[30050] <= 16'b1111111111111111;
        weights1[30051] <= 16'b1111111111110101;
        weights1[30052] <= 16'b1111111111101100;
        weights1[30053] <= 16'b1111111111011011;
        weights1[30054] <= 16'b1111111111011011;
        weights1[30055] <= 16'b1111111111101010;
        weights1[30056] <= 16'b0000000000000000;
        weights1[30057] <= 16'b1111111111111010;
        weights1[30058] <= 16'b1111111111111001;
        weights1[30059] <= 16'b0000000000000100;
        weights1[30060] <= 16'b0000000000000111;
        weights1[30061] <= 16'b0000000000011000;
        weights1[30062] <= 16'b0000000000001000;
        weights1[30063] <= 16'b1111111111111101;
        weights1[30064] <= 16'b1111111111101011;
        weights1[30065] <= 16'b1111111111100101;
        weights1[30066] <= 16'b1111111111011011;
        weights1[30067] <= 16'b1111111111010101;
        weights1[30068] <= 16'b1111111111100101;
        weights1[30069] <= 16'b1111111111110101;
        weights1[30070] <= 16'b1111111111111000;
        weights1[30071] <= 16'b1111111111111100;
        weights1[30072] <= 16'b0000000000000010;
        weights1[30073] <= 16'b0000000000000011;
        weights1[30074] <= 16'b0000000000000110;
        weights1[30075] <= 16'b0000000000000011;
        weights1[30076] <= 16'b0000000000000110;
        weights1[30077] <= 16'b1111111111111000;
        weights1[30078] <= 16'b1111111111111000;
        weights1[30079] <= 16'b1111111111101111;
        weights1[30080] <= 16'b1111111111101101;
        weights1[30081] <= 16'b1111111111101100;
        weights1[30082] <= 16'b1111111111100000;
        weights1[30083] <= 16'b1111111111111011;
        weights1[30084] <= 16'b1111111111111001;
        weights1[30085] <= 16'b1111111111111000;
        weights1[30086] <= 16'b1111111111100111;
        weights1[30087] <= 16'b1111111111110010;
        weights1[30088] <= 16'b1111111111111111;
        weights1[30089] <= 16'b0000000000010100;
        weights1[30090] <= 16'b0000000000001001;
        weights1[30091] <= 16'b1111111111110100;
        weights1[30092] <= 16'b1111111111101010;
        weights1[30093] <= 16'b1111111111011001;
        weights1[30094] <= 16'b1111111111010001;
        weights1[30095] <= 16'b1111111111010010;
        weights1[30096] <= 16'b1111111111100010;
        weights1[30097] <= 16'b1111111111101001;
        weights1[30098] <= 16'b1111111111110010;
        weights1[30099] <= 16'b1111111111111100;
        weights1[30100] <= 16'b0000000000000001;
        weights1[30101] <= 16'b1111111111111111;
        weights1[30102] <= 16'b0000000000000100;
        weights1[30103] <= 16'b0000000000000101;
        weights1[30104] <= 16'b1111111111111111;
        weights1[30105] <= 16'b1111111111111101;
        weights1[30106] <= 16'b1111111111111010;
        weights1[30107] <= 16'b1111111111101100;
        weights1[30108] <= 16'b1111111111100000;
        weights1[30109] <= 16'b1111111111101010;
        weights1[30110] <= 16'b1111111111100010;
        weights1[30111] <= 16'b1111111111111100;
        weights1[30112] <= 16'b1111111111111010;
        weights1[30113] <= 16'b1111111111110011;
        weights1[30114] <= 16'b1111111111101011;
        weights1[30115] <= 16'b1111111111110110;
        weights1[30116] <= 16'b0000000000010101;
        weights1[30117] <= 16'b0000000000100001;
        weights1[30118] <= 16'b0000000000001011;
        weights1[30119] <= 16'b0000000000000010;
        weights1[30120] <= 16'b1111111111110110;
        weights1[30121] <= 16'b1111111111011011;
        weights1[30122] <= 16'b1111111111001000;
        weights1[30123] <= 16'b1111111111010100;
        weights1[30124] <= 16'b1111111111100001;
        weights1[30125] <= 16'b1111111111101101;
        weights1[30126] <= 16'b1111111111110101;
        weights1[30127] <= 16'b1111111111111000;
        weights1[30128] <= 16'b0000000000000001;
        weights1[30129] <= 16'b1111111111111011;
        weights1[30130] <= 16'b1111111111111111;
        weights1[30131] <= 16'b0000000000001000;
        weights1[30132] <= 16'b0000000000000010;
        weights1[30133] <= 16'b0000000000000101;
        weights1[30134] <= 16'b1111111111111000;
        weights1[30135] <= 16'b1111111111101101;
        weights1[30136] <= 16'b1111111111101000;
        weights1[30137] <= 16'b1111111111101110;
        weights1[30138] <= 16'b1111111111111001;
        weights1[30139] <= 16'b1111111111111110;
        weights1[30140] <= 16'b1111111111110010;
        weights1[30141] <= 16'b1111111111100011;
        weights1[30142] <= 16'b1111111111101010;
        weights1[30143] <= 16'b0000000000000100;
        weights1[30144] <= 16'b0000000000011100;
        weights1[30145] <= 16'b0000000000011000;
        weights1[30146] <= 16'b0000000000000110;
        weights1[30147] <= 16'b0000000000000000;
        weights1[30148] <= 16'b1111111111110011;
        weights1[30149] <= 16'b1111111111100010;
        weights1[30150] <= 16'b1111111111010001;
        weights1[30151] <= 16'b1111111111010100;
        weights1[30152] <= 16'b1111111111100110;
        weights1[30153] <= 16'b1111111111101110;
        weights1[30154] <= 16'b1111111111110100;
        weights1[30155] <= 16'b1111111111111010;
        weights1[30156] <= 16'b1111111111111111;
        weights1[30157] <= 16'b0000000000000000;
        weights1[30158] <= 16'b0000000000000011;
        weights1[30159] <= 16'b0000000000000001;
        weights1[30160] <= 16'b0000000000000001;
        weights1[30161] <= 16'b0000000000000111;
        weights1[30162] <= 16'b1111111111111111;
        weights1[30163] <= 16'b1111111111110010;
        weights1[30164] <= 16'b1111111111111011;
        weights1[30165] <= 16'b1111111111110101;
        weights1[30166] <= 16'b0000000000000000;
        weights1[30167] <= 16'b1111111111111010;
        weights1[30168] <= 16'b1111111111110000;
        weights1[30169] <= 16'b1111111111101000;
        weights1[30170] <= 16'b1111111111101011;
        weights1[30171] <= 16'b0000000000000111;
        weights1[30172] <= 16'b0000000000011001;
        weights1[30173] <= 16'b0000000000011000;
        weights1[30174] <= 16'b0000000000010000;
        weights1[30175] <= 16'b0000000000000100;
        weights1[30176] <= 16'b1111111111101110;
        weights1[30177] <= 16'b1111111111100000;
        weights1[30178] <= 16'b1111111111011110;
        weights1[30179] <= 16'b1111111111101010;
        weights1[30180] <= 16'b1111111111101100;
        weights1[30181] <= 16'b1111111111110111;
        weights1[30182] <= 16'b1111111111111001;
        weights1[30183] <= 16'b1111111111111111;
        weights1[30184] <= 16'b0000000000000001;
        weights1[30185] <= 16'b0000000000000010;
        weights1[30186] <= 16'b0000000000000000;
        weights1[30187] <= 16'b0000000000000011;
        weights1[30188] <= 16'b1111111111111101;
        weights1[30189] <= 16'b0000000000000101;
        weights1[30190] <= 16'b1111111111111011;
        weights1[30191] <= 16'b0000000000000000;
        weights1[30192] <= 16'b1111111111111110;
        weights1[30193] <= 16'b0000000000000110;
        weights1[30194] <= 16'b0000000000000000;
        weights1[30195] <= 16'b1111111111111010;
        weights1[30196] <= 16'b1111111111101010;
        weights1[30197] <= 16'b1111111111010111;
        weights1[30198] <= 16'b1111111111100100;
        weights1[30199] <= 16'b0000000000000000;
        weights1[30200] <= 16'b0000000000011010;
        weights1[30201] <= 16'b0000000000011011;
        weights1[30202] <= 16'b0000000000001100;
        weights1[30203] <= 16'b0000000000000111;
        weights1[30204] <= 16'b1111111111111011;
        weights1[30205] <= 16'b1111111111101100;
        weights1[30206] <= 16'b1111111111100001;
        weights1[30207] <= 16'b1111111111110110;
        weights1[30208] <= 16'b1111111111111000;
        weights1[30209] <= 16'b1111111111111100;
        weights1[30210] <= 16'b1111111111111110;
        weights1[30211] <= 16'b1111111111111100;
        weights1[30212] <= 16'b0000000000000011;
        weights1[30213] <= 16'b1111111111111110;
        weights1[30214] <= 16'b0000000000000010;
        weights1[30215] <= 16'b1111111111111100;
        weights1[30216] <= 16'b1111111111111100;
        weights1[30217] <= 16'b0000000000000011;
        weights1[30218] <= 16'b0000000000000100;
        weights1[30219] <= 16'b1111111111111110;
        weights1[30220] <= 16'b0000000000000101;
        weights1[30221] <= 16'b0000000000000001;
        weights1[30222] <= 16'b0000000000000011;
        weights1[30223] <= 16'b1111111111110101;
        weights1[30224] <= 16'b1111111111100100;
        weights1[30225] <= 16'b1111111111010001;
        weights1[30226] <= 16'b1111111111101011;
        weights1[30227] <= 16'b0000000000001011;
        weights1[30228] <= 16'b0000000000011111;
        weights1[30229] <= 16'b0000000000011110;
        weights1[30230] <= 16'b0000000000001110;
        weights1[30231] <= 16'b0000000000000001;
        weights1[30232] <= 16'b1111111111110010;
        weights1[30233] <= 16'b1111111111100101;
        weights1[30234] <= 16'b1111111111110001;
        weights1[30235] <= 16'b1111111111111011;
        weights1[30236] <= 16'b1111111111111000;
        weights1[30237] <= 16'b0000000000000001;
        weights1[30238] <= 16'b0000000000000001;
        weights1[30239] <= 16'b1111111111111011;
        weights1[30240] <= 16'b0000000000000101;
        weights1[30241] <= 16'b1111111111111011;
        weights1[30242] <= 16'b0000000000000011;
        weights1[30243] <= 16'b1111111111111001;
        weights1[30244] <= 16'b1111111111111111;
        weights1[30245] <= 16'b0000000000000000;
        weights1[30246] <= 16'b0000000000001011;
        weights1[30247] <= 16'b0000000000010000;
        weights1[30248] <= 16'b1111111111111100;
        weights1[30249] <= 16'b1111111111111001;
        weights1[30250] <= 16'b1111111111111001;
        weights1[30251] <= 16'b1111111111011100;
        weights1[30252] <= 16'b1111111111100100;
        weights1[30253] <= 16'b1111111111010100;
        weights1[30254] <= 16'b1111111111100010;
        weights1[30255] <= 16'b0000000000010011;
        weights1[30256] <= 16'b0000000000010010;
        weights1[30257] <= 16'b0000000000011001;
        weights1[30258] <= 16'b0000000000010110;
        weights1[30259] <= 16'b0000000000001000;
        weights1[30260] <= 16'b1111111111111110;
        weights1[30261] <= 16'b1111111111110010;
        weights1[30262] <= 16'b1111111111110100;
        weights1[30263] <= 16'b1111111111111111;
        weights1[30264] <= 16'b0000000000000011;
        weights1[30265] <= 16'b0000000000001000;
        weights1[30266] <= 16'b0000000000000000;
        weights1[30267] <= 16'b1111111111111101;
        weights1[30268] <= 16'b0000000000000001;
        weights1[30269] <= 16'b0000000000000000;
        weights1[30270] <= 16'b1111111111111111;
        weights1[30271] <= 16'b1111111111111101;
        weights1[30272] <= 16'b0000000000000110;
        weights1[30273] <= 16'b0000000000000010;
        weights1[30274] <= 16'b0000000000000001;
        weights1[30275] <= 16'b0000000000000011;
        weights1[30276] <= 16'b1111111111111011;
        weights1[30277] <= 16'b1111111111111000;
        weights1[30278] <= 16'b1111111111101111;
        weights1[30279] <= 16'b1111111111100100;
        weights1[30280] <= 16'b1111111111100000;
        weights1[30281] <= 16'b1111111111001001;
        weights1[30282] <= 16'b1111111111101001;
        weights1[30283] <= 16'b0000000000010110;
        weights1[30284] <= 16'b0000000000010010;
        weights1[30285] <= 16'b0000000000010110;
        weights1[30286] <= 16'b0000000000001110;
        weights1[30287] <= 16'b1111111111111010;
        weights1[30288] <= 16'b1111111111111001;
        weights1[30289] <= 16'b1111111111110001;
        weights1[30290] <= 16'b1111111111111110;
        weights1[30291] <= 16'b0000000000001010;
        weights1[30292] <= 16'b0000000000001011;
        weights1[30293] <= 16'b0000000000010000;
        weights1[30294] <= 16'b0000000000000011;
        weights1[30295] <= 16'b0000000000000000;
        weights1[30296] <= 16'b1111111111111111;
        weights1[30297] <= 16'b0000000000000001;
        weights1[30298] <= 16'b1111111111111111;
        weights1[30299] <= 16'b1111111111111101;
        weights1[30300] <= 16'b0000000000000011;
        weights1[30301] <= 16'b0000000000000010;
        weights1[30302] <= 16'b1111111111111100;
        weights1[30303] <= 16'b1111111111110101;
        weights1[30304] <= 16'b1111111111110010;
        weights1[30305] <= 16'b1111111111101010;
        weights1[30306] <= 16'b1111111111100010;
        weights1[30307] <= 16'b1111111111100000;
        weights1[30308] <= 16'b1111111111010100;
        weights1[30309] <= 16'b1111111111001011;
        weights1[30310] <= 16'b1111111111101010;
        weights1[30311] <= 16'b0000000000001010;
        weights1[30312] <= 16'b0000000000010010;
        weights1[30313] <= 16'b0000000000010011;
        weights1[30314] <= 16'b0000000000000110;
        weights1[30315] <= 16'b0000000000000010;
        weights1[30316] <= 16'b1111111111111011;
        weights1[30317] <= 16'b0000000000000100;
        weights1[30318] <= 16'b0000000000011000;
        weights1[30319] <= 16'b0000000000010001;
        weights1[30320] <= 16'b0000000000010110;
        weights1[30321] <= 16'b0000000000001101;
        weights1[30322] <= 16'b0000000000001000;
        weights1[30323] <= 16'b0000000000000000;
        weights1[30324] <= 16'b1111111111111110;
        weights1[30325] <= 16'b0000000000000001;
        weights1[30326] <= 16'b1111111111111011;
        weights1[30327] <= 16'b1111111111111100;
        weights1[30328] <= 16'b0000000000000001;
        weights1[30329] <= 16'b1111111111110100;
        weights1[30330] <= 16'b1111111111110110;
        weights1[30331] <= 16'b1111111111101110;
        weights1[30332] <= 16'b1111111111100111;
        weights1[30333] <= 16'b1111111111011111;
        weights1[30334] <= 16'b1111111111010011;
        weights1[30335] <= 16'b1111111111011000;
        weights1[30336] <= 16'b1111111111011011;
        weights1[30337] <= 16'b1111111111011111;
        weights1[30338] <= 16'b1111111111110001;
        weights1[30339] <= 16'b1111111111111111;
        weights1[30340] <= 16'b0000000000010100;
        weights1[30341] <= 16'b0000000000010010;
        weights1[30342] <= 16'b0000000000001010;
        weights1[30343] <= 16'b1111111111111101;
        weights1[30344] <= 16'b0000000000000011;
        weights1[30345] <= 16'b0000000000000101;
        weights1[30346] <= 16'b0000000000011001;
        weights1[30347] <= 16'b0000000000010010;
        weights1[30348] <= 16'b0000000000010101;
        weights1[30349] <= 16'b0000000000010000;
        weights1[30350] <= 16'b0000000000001100;
        weights1[30351] <= 16'b0000000000000011;
        weights1[30352] <= 16'b1111111111111100;
        weights1[30353] <= 16'b1111111111111110;
        weights1[30354] <= 16'b1111111111111011;
        weights1[30355] <= 16'b1111111111111000;
        weights1[30356] <= 16'b1111111111111101;
        weights1[30357] <= 16'b1111111111101111;
        weights1[30358] <= 16'b1111111111110001;
        weights1[30359] <= 16'b1111111111110100;
        weights1[30360] <= 16'b1111111111100110;
        weights1[30361] <= 16'b1111111111011010;
        weights1[30362] <= 16'b1111111111010101;
        weights1[30363] <= 16'b1111111111001111;
        weights1[30364] <= 16'b1111111111100111;
        weights1[30365] <= 16'b1111111111101001;
        weights1[30366] <= 16'b1111111111111100;
        weights1[30367] <= 16'b0000000000000011;
        weights1[30368] <= 16'b0000000000010011;
        weights1[30369] <= 16'b0000000000010001;
        weights1[30370] <= 16'b0000000000001101;
        weights1[30371] <= 16'b0000000000001000;
        weights1[30372] <= 16'b0000000000001110;
        weights1[30373] <= 16'b0000000000001000;
        weights1[30374] <= 16'b0000000000010010;
        weights1[30375] <= 16'b0000000000010110;
        weights1[30376] <= 16'b0000000000001101;
        weights1[30377] <= 16'b0000000000000100;
        weights1[30378] <= 16'b0000000000001001;
        weights1[30379] <= 16'b0000000000000110;
        weights1[30380] <= 16'b1111111111111111;
        weights1[30381] <= 16'b1111111111111110;
        weights1[30382] <= 16'b1111111111111001;
        weights1[30383] <= 16'b1111111111111010;
        weights1[30384] <= 16'b1111111111110110;
        weights1[30385] <= 16'b1111111111111001;
        weights1[30386] <= 16'b1111111111110110;
        weights1[30387] <= 16'b1111111111110100;
        weights1[30388] <= 16'b1111111111101101;
        weights1[30389] <= 16'b1111111111100110;
        weights1[30390] <= 16'b1111111111011001;
        weights1[30391] <= 16'b1111111111010110;
        weights1[30392] <= 16'b1111111111100000;
        weights1[30393] <= 16'b1111111111111001;
        weights1[30394] <= 16'b0000000000001000;
        weights1[30395] <= 16'b0000000000010000;
        weights1[30396] <= 16'b0000000000010011;
        weights1[30397] <= 16'b0000000000011001;
        weights1[30398] <= 16'b0000000000000111;
        weights1[30399] <= 16'b0000000000000111;
        weights1[30400] <= 16'b0000000000001110;
        weights1[30401] <= 16'b0000000000001011;
        weights1[30402] <= 16'b0000000000001110;
        weights1[30403] <= 16'b0000000000001000;
        weights1[30404] <= 16'b0000000000001101;
        weights1[30405] <= 16'b1111111111111100;
        weights1[30406] <= 16'b0000000000000010;
        weights1[30407] <= 16'b1111111111111111;
        weights1[30408] <= 16'b1111111111111110;
        weights1[30409] <= 16'b1111111111111101;
        weights1[30410] <= 16'b1111111111111000;
        weights1[30411] <= 16'b1111111111110101;
        weights1[30412] <= 16'b1111111111110011;
        weights1[30413] <= 16'b1111111111110011;
        weights1[30414] <= 16'b1111111111111001;
        weights1[30415] <= 16'b1111111111110110;
        weights1[30416] <= 16'b1111111111110010;
        weights1[30417] <= 16'b1111111111110000;
        weights1[30418] <= 16'b1111111111101110;
        weights1[30419] <= 16'b1111111111111011;
        weights1[30420] <= 16'b1111111111111011;
        weights1[30421] <= 16'b0000000000000001;
        weights1[30422] <= 16'b0000000000000101;
        weights1[30423] <= 16'b0000000000010001;
        weights1[30424] <= 16'b0000000000001110;
        weights1[30425] <= 16'b0000000000011011;
        weights1[30426] <= 16'b0000000000010001;
        weights1[30427] <= 16'b0000000000000110;
        weights1[30428] <= 16'b0000000000001010;
        weights1[30429] <= 16'b0000000000001011;
        weights1[30430] <= 16'b0000000000010000;
        weights1[30431] <= 16'b0000000000001100;
        weights1[30432] <= 16'b0000000000001101;
        weights1[30433] <= 16'b0000000000000111;
        weights1[30434] <= 16'b0000000000000011;
        weights1[30435] <= 16'b0000000000000001;
        weights1[30436] <= 16'b1111111111111110;
        weights1[30437] <= 16'b1111111111111110;
        weights1[30438] <= 16'b1111111111111001;
        weights1[30439] <= 16'b1111111111110110;
        weights1[30440] <= 16'b1111111111101110;
        weights1[30441] <= 16'b1111111111110011;
        weights1[30442] <= 16'b1111111111101110;
        weights1[30443] <= 16'b1111111111110001;
        weights1[30444] <= 16'b1111111111110000;
        weights1[30445] <= 16'b1111111111110000;
        weights1[30446] <= 16'b0000000000000001;
        weights1[30447] <= 16'b0000000000000101;
        weights1[30448] <= 16'b0000000000001010;
        weights1[30449] <= 16'b1111111111111110;
        weights1[30450] <= 16'b1111111111111000;
        weights1[30451] <= 16'b0000000000001100;
        weights1[30452] <= 16'b0000000000000000;
        weights1[30453] <= 16'b0000000000000111;
        weights1[30454] <= 16'b0000000000010100;
        weights1[30455] <= 16'b0000000000000010;
        weights1[30456] <= 16'b0000000000000111;
        weights1[30457] <= 16'b0000000000000111;
        weights1[30458] <= 16'b0000000000001010;
        weights1[30459] <= 16'b0000000000001001;
        weights1[30460] <= 16'b0000000000000001;
        weights1[30461] <= 16'b0000000000000011;
        weights1[30462] <= 16'b0000000000000011;
        weights1[30463] <= 16'b0000000000000010;
        weights1[30464] <= 16'b1111111111111111;
        weights1[30465] <= 16'b1111111111111110;
        weights1[30466] <= 16'b1111111111111001;
        weights1[30467] <= 16'b1111111111111000;
        weights1[30468] <= 16'b1111111111101111;
        weights1[30469] <= 16'b1111111111110001;
        weights1[30470] <= 16'b1111111111110001;
        weights1[30471] <= 16'b1111111111111000;
        weights1[30472] <= 16'b1111111111101110;
        weights1[30473] <= 16'b1111111111110110;
        weights1[30474] <= 16'b0000000000000000;
        weights1[30475] <= 16'b0000000000000011;
        weights1[30476] <= 16'b0000000000001011;
        weights1[30477] <= 16'b0000000000000111;
        weights1[30478] <= 16'b0000000000000001;
        weights1[30479] <= 16'b0000000000000011;
        weights1[30480] <= 16'b0000000000010010;
        weights1[30481] <= 16'b0000000000001100;
        weights1[30482] <= 16'b0000000000001011;
        weights1[30483] <= 16'b0000000000000001;
        weights1[30484] <= 16'b0000000000000111;
        weights1[30485] <= 16'b0000000000000100;
        weights1[30486] <= 16'b0000000000000110;
        weights1[30487] <= 16'b0000000000000110;
        weights1[30488] <= 16'b0000000000000011;
        weights1[30489] <= 16'b1111111111111111;
        weights1[30490] <= 16'b1111111111111101;
        weights1[30491] <= 16'b0000000000000001;
        weights1[30492] <= 16'b1111111111111111;
        weights1[30493] <= 16'b1111111111111110;
        weights1[30494] <= 16'b1111111111111100;
        weights1[30495] <= 16'b1111111111111110;
        weights1[30496] <= 16'b1111111111110100;
        weights1[30497] <= 16'b1111111111101101;
        weights1[30498] <= 16'b1111111111101111;
        weights1[30499] <= 16'b1111111111110101;
        weights1[30500] <= 16'b1111111111111001;
        weights1[30501] <= 16'b0000000000000100;
        weights1[30502] <= 16'b0000000000001010;
        weights1[30503] <= 16'b0000000000001101;
        weights1[30504] <= 16'b1111111111111010;
        weights1[30505] <= 16'b1111111111111110;
        weights1[30506] <= 16'b1111111111111101;
        weights1[30507] <= 16'b1111111111111110;
        weights1[30508] <= 16'b0000000000001011;
        weights1[30509] <= 16'b0000000000010010;
        weights1[30510] <= 16'b0000000000000110;
        weights1[30511] <= 16'b0000000000001000;
        weights1[30512] <= 16'b0000000000001101;
        weights1[30513] <= 16'b0000000000010000;
        weights1[30514] <= 16'b0000000000001010;
        weights1[30515] <= 16'b0000000000000100;
        weights1[30516] <= 16'b0000000000000010;
        weights1[30517] <= 16'b0000000000000000;
        weights1[30518] <= 16'b1111111111111111;
        weights1[30519] <= 16'b1111111111111111;
        weights1[30520] <= 16'b1111111111111101;
        weights1[30521] <= 16'b1111111111111101;
        weights1[30522] <= 16'b1111111111111111;
        weights1[30523] <= 16'b1111111111111110;
        weights1[30524] <= 16'b1111111111111001;
        weights1[30525] <= 16'b1111111111110101;
        weights1[30526] <= 16'b1111111111110101;
        weights1[30527] <= 16'b1111111111111001;
        weights1[30528] <= 16'b1111111111111100;
        weights1[30529] <= 16'b0000000000000111;
        weights1[30530] <= 16'b0000000000001011;
        weights1[30531] <= 16'b0000000000001001;
        weights1[30532] <= 16'b0000000000000001;
        weights1[30533] <= 16'b1111111111111110;
        weights1[30534] <= 16'b0000000000000110;
        weights1[30535] <= 16'b0000000000010001;
        weights1[30536] <= 16'b0000000000001101;
        weights1[30537] <= 16'b0000000000001000;
        weights1[30538] <= 16'b1111111111111010;
        weights1[30539] <= 16'b0000000000000000;
        weights1[30540] <= 16'b0000000000000110;
        weights1[30541] <= 16'b0000000000001101;
        weights1[30542] <= 16'b0000000000001001;
        weights1[30543] <= 16'b1111111111111111;
        weights1[30544] <= 16'b0000000000000000;
        weights1[30545] <= 16'b1111111111111111;
        weights1[30546] <= 16'b1111111111111111;
        weights1[30547] <= 16'b0000000000000000;
        weights1[30548] <= 16'b1111111111111110;
        weights1[30549] <= 16'b1111111111111110;
        weights1[30550] <= 16'b1111111111111110;
        weights1[30551] <= 16'b1111111111111111;
        weights1[30552] <= 16'b1111111111111101;
        weights1[30553] <= 16'b1111111111111101;
        weights1[30554] <= 16'b1111111111111110;
        weights1[30555] <= 16'b0000000000000101;
        weights1[30556] <= 16'b0000000000000100;
        weights1[30557] <= 16'b0000000000000110;
        weights1[30558] <= 16'b0000000000001000;
        weights1[30559] <= 16'b0000000000001111;
        weights1[30560] <= 16'b0000000000001100;
        weights1[30561] <= 16'b0000000000001010;
        weights1[30562] <= 16'b0000000000001011;
        weights1[30563] <= 16'b0000000000001010;
        weights1[30564] <= 16'b0000000000011010;
        weights1[30565] <= 16'b0000000000001111;
        weights1[30566] <= 16'b0000000000001001;
        weights1[30567] <= 16'b0000000000010010;
        weights1[30568] <= 16'b0000000000001000;
        weights1[30569] <= 16'b0000000000001001;
        weights1[30570] <= 16'b0000000000000100;
        weights1[30571] <= 16'b0000000000000011;
        weights1[30572] <= 16'b0000000000000010;
        weights1[30573] <= 16'b1111111111111111;
        weights1[30574] <= 16'b1111111111111111;
        weights1[30575] <= 16'b0000000000000000;
        weights1[30576] <= 16'b0000000000000001;
        weights1[30577] <= 16'b0000000000000001;
        weights1[30578] <= 16'b0000000000000001;
        weights1[30579] <= 16'b0000000000000000;
        weights1[30580] <= 16'b1111111111111101;
        weights1[30581] <= 16'b1111111111110111;
        weights1[30582] <= 16'b1111111111110110;
        weights1[30583] <= 16'b1111111111101110;
        weights1[30584] <= 16'b1111111111101011;
        weights1[30585] <= 16'b1111111111111101;
        weights1[30586] <= 16'b0000000000000001;
        weights1[30587] <= 16'b1111111111110101;
        weights1[30588] <= 16'b1111111111110101;
        weights1[30589] <= 16'b1111111111111111;
        weights1[30590] <= 16'b1111111111110110;
        weights1[30591] <= 16'b1111111111110000;
        weights1[30592] <= 16'b1111111111110000;
        weights1[30593] <= 16'b1111111111110011;
        weights1[30594] <= 16'b1111111111111101;
        weights1[30595] <= 16'b1111111111111111;
        weights1[30596] <= 16'b1111111111110110;
        weights1[30597] <= 16'b0000000000000101;
        weights1[30598] <= 16'b1111111111111111;
        weights1[30599] <= 16'b0000000000001101;
        weights1[30600] <= 16'b0000000000001000;
        weights1[30601] <= 16'b0000000000001000;
        weights1[30602] <= 16'b0000000000001000;
        weights1[30603] <= 16'b1111111111111110;
        weights1[30604] <= 16'b0000000000000001;
        weights1[30605] <= 16'b0000000000000000;
        weights1[30606] <= 16'b0000000000000000;
        weights1[30607] <= 16'b1111111111111111;
        weights1[30608] <= 16'b1111111111111101;
        weights1[30609] <= 16'b1111111111111111;
        weights1[30610] <= 16'b1111111111111100;
        weights1[30611] <= 16'b1111111111111110;
        weights1[30612] <= 16'b0000000000000011;
        weights1[30613] <= 16'b1111111111111001;
        weights1[30614] <= 16'b1111111111111100;
        weights1[30615] <= 16'b1111111111101110;
        weights1[30616] <= 16'b1111111111111011;
        weights1[30617] <= 16'b1111111111110100;
        weights1[30618] <= 16'b1111111111111001;
        weights1[30619] <= 16'b1111111111110111;
        weights1[30620] <= 16'b1111111111110001;
        weights1[30621] <= 16'b1111111111110001;
        weights1[30622] <= 16'b1111111111110001;
        weights1[30623] <= 16'b0000000000001001;
        weights1[30624] <= 16'b1111111111110001;
        weights1[30625] <= 16'b1111111111110100;
        weights1[30626] <= 16'b0000000000000110;
        weights1[30627] <= 16'b1111111111111101;
        weights1[30628] <= 16'b0000000000000101;
        weights1[30629] <= 16'b0000000000010000;
        weights1[30630] <= 16'b0000000000001101;
        weights1[30631] <= 16'b0000000000000110;
        weights1[30632] <= 16'b0000000000000011;
        weights1[30633] <= 16'b0000000000000011;
        weights1[30634] <= 16'b0000000000000111;
        weights1[30635] <= 16'b0000000000000001;
        weights1[30636] <= 16'b0000000000000011;
        weights1[30637] <= 16'b1111111111111111;
        weights1[30638] <= 16'b0000000000000010;
        weights1[30639] <= 16'b0000000000000011;
        weights1[30640] <= 16'b1111111111110010;
        weights1[30641] <= 16'b1111111111111110;
        weights1[30642] <= 16'b0000000000000111;
        weights1[30643] <= 16'b1111111111111111;
        weights1[30644] <= 16'b0000000000000001;
        weights1[30645] <= 16'b1111111111111011;
        weights1[30646] <= 16'b1111111111111000;
        weights1[30647] <= 16'b0000000000000100;
        weights1[30648] <= 16'b0000000000000010;
        weights1[30649] <= 16'b0000000000000100;
        weights1[30650] <= 16'b0000000000001011;
        weights1[30651] <= 16'b0000000000000111;
        weights1[30652] <= 16'b0000000000001100;
        weights1[30653] <= 16'b0000000000000111;
        weights1[30654] <= 16'b1111111111111010;
        weights1[30655] <= 16'b0000000000000111;
        weights1[30656] <= 16'b0000000000010010;
        weights1[30657] <= 16'b0000000000001111;
        weights1[30658] <= 16'b0000000000010010;
        weights1[30659] <= 16'b0000000000001100;
        weights1[30660] <= 16'b0000000000001001;
        weights1[30661] <= 16'b0000000000000101;
        weights1[30662] <= 16'b0000000000000110;
        weights1[30663] <= 16'b0000000000001010;
        weights1[30664] <= 16'b0000000000000011;
        weights1[30665] <= 16'b0000000000001010;
        weights1[30666] <= 16'b0000000000000000;
        weights1[30667] <= 16'b0000000000000010;
        weights1[30668] <= 16'b0000000000000101;
        weights1[30669] <= 16'b0000000000010001;
        weights1[30670] <= 16'b1111111111111000;
        weights1[30671] <= 16'b0000000000001011;
        weights1[30672] <= 16'b1111111111111001;
        weights1[30673] <= 16'b1111111111111101;
        weights1[30674] <= 16'b0000000000000001;
        weights1[30675] <= 16'b1111111111110101;
        weights1[30676] <= 16'b0000000000000001;
        weights1[30677] <= 16'b1111111111110000;
        weights1[30678] <= 16'b1111111111110110;
        weights1[30679] <= 16'b1111111111111010;
        weights1[30680] <= 16'b0000000000000000;
        weights1[30681] <= 16'b0000000000000101;
        weights1[30682] <= 16'b0000000000000111;
        weights1[30683] <= 16'b0000000000001101;
        weights1[30684] <= 16'b0000000000010111;
        weights1[30685] <= 16'b0000000000000010;
        weights1[30686] <= 16'b0000000000010000;
        weights1[30687] <= 16'b0000000000001001;
        weights1[30688] <= 16'b0000000000001100;
        weights1[30689] <= 16'b0000000000000101;
        weights1[30690] <= 16'b0000000000010000;
        weights1[30691] <= 16'b0000000000010100;
        weights1[30692] <= 16'b0000000000100000;
        weights1[30693] <= 16'b0000000000010101;
        weights1[30694] <= 16'b0000000000000010;
        weights1[30695] <= 16'b0000000000000001;
        weights1[30696] <= 16'b1111111111110001;
        weights1[30697] <= 16'b1111111111111010;
        weights1[30698] <= 16'b1111111111100111;
        weights1[30699] <= 16'b1111111111111001;
        weights1[30700] <= 16'b0000000000001100;
        weights1[30701] <= 16'b0000000000000011;
        weights1[30702] <= 16'b1111111111111110;
        weights1[30703] <= 16'b1111111111111110;
        weights1[30704] <= 16'b0000000000001001;
        weights1[30705] <= 16'b0000000000011001;
        weights1[30706] <= 16'b0000000000010001;
        weights1[30707] <= 16'b0000000000010100;
        weights1[30708] <= 16'b1111111111111011;
        weights1[30709] <= 16'b0000000000000101;
        weights1[30710] <= 16'b1111111111111110;
        weights1[30711] <= 16'b1111111111110110;
        weights1[30712] <= 16'b1111111111111111;
        weights1[30713] <= 16'b0000000000010011;
        weights1[30714] <= 16'b0000000000001010;
        weights1[30715] <= 16'b0000000000001101;
        weights1[30716] <= 16'b0000000000010100;
        weights1[30717] <= 16'b0000000000010100;
        weights1[30718] <= 16'b0000000000010010;
        weights1[30719] <= 16'b0000000000011011;
        weights1[30720] <= 16'b0000000000011011;
        weights1[30721] <= 16'b0000000000011001;
        weights1[30722] <= 16'b0000000000001001;
        weights1[30723] <= 16'b0000000000011001;
        weights1[30724] <= 16'b0000000000000011;
        weights1[30725] <= 16'b1111111111111101;
        weights1[30726] <= 16'b0000000000000000;
        weights1[30727] <= 16'b0000000000001010;
        weights1[30728] <= 16'b1111111111111111;
        weights1[30729] <= 16'b0000000000001001;
        weights1[30730] <= 16'b1111111111111101;
        weights1[30731] <= 16'b0000000000010111;
        weights1[30732] <= 16'b0000000000001001;
        weights1[30733] <= 16'b0000000000011011;
        weights1[30734] <= 16'b0000000000010101;
        weights1[30735] <= 16'b0000000000000100;
        weights1[30736] <= 16'b0000000000001110;
        weights1[30737] <= 16'b0000000000001011;
        weights1[30738] <= 16'b0000000000010000;
        weights1[30739] <= 16'b0000000000000011;
        weights1[30740] <= 16'b0000000000001010;
        weights1[30741] <= 16'b0000000000001101;
        weights1[30742] <= 16'b0000000000011101;
        weights1[30743] <= 16'b0000000000010101;
        weights1[30744] <= 16'b0000000000010010;
        weights1[30745] <= 16'b0000000000010001;
        weights1[30746] <= 16'b0000000000010101;
        weights1[30747] <= 16'b0000000000101010;
        weights1[30748] <= 16'b0000000000101010;
        weights1[30749] <= 16'b0000000000101100;
        weights1[30750] <= 16'b0000000000101001;
        weights1[30751] <= 16'b0000000000011011;
        weights1[30752] <= 16'b0000000000011010;
        weights1[30753] <= 16'b0000000000010101;
        weights1[30754] <= 16'b0000000000001000;
        weights1[30755] <= 16'b0000000000000111;
        weights1[30756] <= 16'b0000000000001000;
        weights1[30757] <= 16'b0000000000001100;
        weights1[30758] <= 16'b0000000000001111;
        weights1[30759] <= 16'b0000000000001011;
        weights1[30760] <= 16'b0000000000001110;
        weights1[30761] <= 16'b0000000000001000;
        weights1[30762] <= 16'b0000000000010101;
        weights1[30763] <= 16'b0000000000000101;
        weights1[30764] <= 16'b1111111111110010;
        weights1[30765] <= 16'b0000000000001111;
        weights1[30766] <= 16'b0000000000010101;
        weights1[30767] <= 16'b0000000000001111;
        weights1[30768] <= 16'b0000000000011000;
        weights1[30769] <= 16'b0000000000000100;
        weights1[30770] <= 16'b0000000000010101;
        weights1[30771] <= 16'b0000000000011100;
        weights1[30772] <= 16'b0000000000001100;
        weights1[30773] <= 16'b0000000000001100;
        weights1[30774] <= 16'b0000000000010011;
        weights1[30775] <= 16'b0000000000101111;
        weights1[30776] <= 16'b0000000000000000;
        weights1[30777] <= 16'b0000000000001111;
        weights1[30778] <= 16'b0000000000010101;
        weights1[30779] <= 16'b0000000001001001;
        weights1[30780] <= 16'b0000000000001110;
        weights1[30781] <= 16'b0000000000100010;
        weights1[30782] <= 16'b0000000000100011;
        weights1[30783] <= 16'b0000000000001111;
        weights1[30784] <= 16'b0000000000010111;
        weights1[30785] <= 16'b0000000000010111;
        weights1[30786] <= 16'b0000000000010110;
        weights1[30787] <= 16'b0000000000010011;
        weights1[30788] <= 16'b0000000000011001;
        weights1[30789] <= 16'b0000000000000010;
        weights1[30790] <= 16'b0000000000001101;
        weights1[30791] <= 16'b0000000000011001;
        weights1[30792] <= 16'b0000000000011001;
        weights1[30793] <= 16'b0000000000011001;
        weights1[30794] <= 16'b0000000000000001;
        weights1[30795] <= 16'b0000000000010000;
        weights1[30796] <= 16'b0000000000010011;
        weights1[30797] <= 16'b0000000000001100;
        weights1[30798] <= 16'b1111111111111010;
        weights1[30799] <= 16'b0000000000100000;
        weights1[30800] <= 16'b0000000000010010;
        weights1[30801] <= 16'b0000000000011011;
        weights1[30802] <= 16'b0000000000011011;
        weights1[30803] <= 16'b0000000000100100;
        weights1[30804] <= 16'b0000000000100111;
        weights1[30805] <= 16'b0000000000011100;
        weights1[30806] <= 16'b0000000000010110;
        weights1[30807] <= 16'b0000000000100111;
        weights1[30808] <= 16'b0000000000100101;
        weights1[30809] <= 16'b0000000000101000;
        weights1[30810] <= 16'b0000000000011010;
        weights1[30811] <= 16'b0000000000110101;
        weights1[30812] <= 16'b0000000000001010;
        weights1[30813] <= 16'b0000000000011110;
        weights1[30814] <= 16'b0000000000010100;
        weights1[30815] <= 16'b0000000000100110;
        weights1[30816] <= 16'b0000000000001011;
        weights1[30817] <= 16'b0000000000001011;
        weights1[30818] <= 16'b0000000000001001;
        weights1[30819] <= 16'b0000000000001011;
        weights1[30820] <= 16'b0000000000001011;
        weights1[30821] <= 16'b0000000000011100;
        weights1[30822] <= 16'b0000000000000110;
        weights1[30823] <= 16'b0000000000000001;
        weights1[30824] <= 16'b0000000000010101;
        weights1[30825] <= 16'b0000000000000011;
        weights1[30826] <= 16'b0000000000001010;
        weights1[30827] <= 16'b0000000000010000;
        weights1[30828] <= 16'b0000000000001100;
        weights1[30829] <= 16'b0000000000011000;
        weights1[30830] <= 16'b0000000000100101;
        weights1[30831] <= 16'b0000000000011111;
        weights1[30832] <= 16'b0000000000101100;
        weights1[30833] <= 16'b0000000000011111;
        weights1[30834] <= 16'b0000000000100110;
        weights1[30835] <= 16'b0000000000010111;
        weights1[30836] <= 16'b0000000000100100;
        weights1[30837] <= 16'b0000000000011000;
        weights1[30838] <= 16'b0000000000011100;
        weights1[30839] <= 16'b0000000000101001;
        weights1[30840] <= 16'b0000000000011101;
        weights1[30841] <= 16'b0000000000011001;
        weights1[30842] <= 16'b0000000000011001;
        weights1[30843] <= 16'b0000000000001101;
        weights1[30844] <= 16'b0000000000100100;
        weights1[30845] <= 16'b0000000000101101;
        weights1[30846] <= 16'b0000000000001111;
        weights1[30847] <= 16'b0000000000001110;
        weights1[30848] <= 16'b0000000000001011;
        weights1[30849] <= 16'b1111111111111110;
        weights1[30850] <= 16'b0000000000011001;
        weights1[30851] <= 16'b0000000000000100;
        weights1[30852] <= 16'b0000000000001101;
        weights1[30853] <= 16'b0000000000010001;
        weights1[30854] <= 16'b0000000000001111;
        weights1[30855] <= 16'b0000000000001101;
        weights1[30856] <= 16'b0000000000001110;
        weights1[30857] <= 16'b0000000000011000;
        weights1[30858] <= 16'b0000000000101010;
        weights1[30859] <= 16'b0000000000100101;
        weights1[30860] <= 16'b0000000000010100;
        weights1[30861] <= 16'b0000000000101100;
        weights1[30862] <= 16'b0000000000010011;
        weights1[30863] <= 16'b0000000000011011;
        weights1[30864] <= 16'b0000000000100111;
        weights1[30865] <= 16'b0000000000011110;
        weights1[30866] <= 16'b0000000000101001;
        weights1[30867] <= 16'b0000000000011000;
        weights1[30868] <= 16'b0000000000011010;
        weights1[30869] <= 16'b0000000000010001;
        weights1[30870] <= 16'b0000000000100011;
        weights1[30871] <= 16'b0000000000110111;
        weights1[30872] <= 16'b0000000000010000;
        weights1[30873] <= 16'b0000000000110001;
        weights1[30874] <= 16'b0000000000011000;
        weights1[30875] <= 16'b0000000000110100;
        weights1[30876] <= 16'b0000000000010101;
        weights1[30877] <= 16'b0000000000011000;
        weights1[30878] <= 16'b0000000000010011;
        weights1[30879] <= 16'b0000000000000110;
        weights1[30880] <= 16'b1111111111111110;
        weights1[30881] <= 16'b0000000000100110;
        weights1[30882] <= 16'b0000000000011010;
        weights1[30883] <= 16'b0000000000000101;
        weights1[30884] <= 16'b0000000000001010;
        weights1[30885] <= 16'b0000000000001110;
        weights1[30886] <= 16'b0000000000010101;
        weights1[30887] <= 16'b0000000000011111;
        weights1[30888] <= 16'b0000000000100001;
        weights1[30889] <= 16'b0000000000011100;
        weights1[30890] <= 16'b0000000000101001;
        weights1[30891] <= 16'b0000000000110010;
        weights1[30892] <= 16'b0000000000100001;
        weights1[30893] <= 16'b0000000000001001;
        weights1[30894] <= 16'b0000000000011011;
        weights1[30895] <= 16'b0000000000100100;
        weights1[30896] <= 16'b0000000000010101;
        weights1[30897] <= 16'b0000000000011001;
        weights1[30898] <= 16'b0000000000101001;
        weights1[30899] <= 16'b0000000000101001;
        weights1[30900] <= 16'b0000000000011010;
        weights1[30901] <= 16'b0000000000100010;
        weights1[30902] <= 16'b0000000000011111;
        weights1[30903] <= 16'b0000000000101100;
        weights1[30904] <= 16'b0000000000100001;
        weights1[30905] <= 16'b0000000000100110;
        weights1[30906] <= 16'b0000000000111011;
        weights1[30907] <= 16'b0000000000111001;
        weights1[30908] <= 16'b0000000000110111;
        weights1[30909] <= 16'b0000000000100011;
        weights1[30910] <= 16'b0000000000101100;
        weights1[30911] <= 16'b0000000000011010;
        weights1[30912] <= 16'b1111111111111101;
        weights1[30913] <= 16'b1111111111110000;
        weights1[30914] <= 16'b0000000000001110;
        weights1[30915] <= 16'b0000000000011010;
        weights1[30916] <= 16'b0000000000100111;
        weights1[30917] <= 16'b0000000000101000;
        weights1[30918] <= 16'b0000000000001000;
        weights1[30919] <= 16'b0000000000010010;
        weights1[30920] <= 16'b0000000000110000;
        weights1[30921] <= 16'b0000000000010001;
        weights1[30922] <= 16'b0000000000011101;
        weights1[30923] <= 16'b0000000000101110;
        weights1[30924] <= 16'b0000000000011111;
        weights1[30925] <= 16'b0000000000011010;
        weights1[30926] <= 16'b0000000000011000;
        weights1[30927] <= 16'b0000000000001100;
        weights1[30928] <= 16'b0000000000100100;
        weights1[30929] <= 16'b0000000000011110;
        weights1[30930] <= 16'b0000000000100110;
        weights1[30931] <= 16'b0000000000101011;
        weights1[30932] <= 16'b0000000000101011;
        weights1[30933] <= 16'b0000000000110011;
        weights1[30934] <= 16'b0000000000110010;
        weights1[30935] <= 16'b0000000000100010;
        weights1[30936] <= 16'b0000000000111000;
        weights1[30937] <= 16'b0000000000100011;
        weights1[30938] <= 16'b0000000000100001;
        weights1[30939] <= 16'b0000000000001111;
        weights1[30940] <= 16'b1111111111110110;
        weights1[30941] <= 16'b1111111111100100;
        weights1[30942] <= 16'b1111111111110010;
        weights1[30943] <= 16'b0000000000011100;
        weights1[30944] <= 16'b0000000000101001;
        weights1[30945] <= 16'b0000000000010111;
        weights1[30946] <= 16'b0000000000001001;
        weights1[30947] <= 16'b0000000000010111;
        weights1[30948] <= 16'b0000000000011101;
        weights1[30949] <= 16'b0000000000001110;
        weights1[30950] <= 16'b0000000000010110;
        weights1[30951] <= 16'b1111111111111100;
        weights1[30952] <= 16'b0000000000011001;
        weights1[30953] <= 16'b0000000000010011;
        weights1[30954] <= 16'b1111111111111101;
        weights1[30955] <= 16'b0000000000001010;
        weights1[30956] <= 16'b1111111111111101;
        weights1[30957] <= 16'b0000000000001011;
        weights1[30958] <= 16'b0000000000001101;
        weights1[30959] <= 16'b0000000000011001;
        weights1[30960] <= 16'b0000000000011110;
        weights1[30961] <= 16'b0000000000001010;
        weights1[30962] <= 16'b0000000000001101;
        weights1[30963] <= 16'b0000000000100111;
        weights1[30964] <= 16'b0000000000100000;
        weights1[30965] <= 16'b0000000000010100;
        weights1[30966] <= 16'b0000000000011010;
        weights1[30967] <= 16'b0000000000000110;
        weights1[30968] <= 16'b1111111111100010;
        weights1[30969] <= 16'b1111111111011000;
        weights1[30970] <= 16'b1111111111010000;
        weights1[30971] <= 16'b1111111111011000;
        weights1[30972] <= 16'b1111111111101111;
        weights1[30973] <= 16'b1111111111100101;
        weights1[30974] <= 16'b1111111111101111;
        weights1[30975] <= 16'b1111111111111001;
        weights1[30976] <= 16'b1111111111111111;
        weights1[30977] <= 16'b1111111111011100;
        weights1[30978] <= 16'b1111111110110101;
        weights1[30979] <= 16'b1111111110111100;
        weights1[30980] <= 16'b1111111111000000;
        weights1[30981] <= 16'b1111111111001100;
        weights1[30982] <= 16'b1111111111010110;
        weights1[30983] <= 16'b1111111111011000;
        weights1[30984] <= 16'b1111111111110100;
        weights1[30985] <= 16'b1111111111100011;
        weights1[30986] <= 16'b1111111111011001;
        weights1[30987] <= 16'b1111111111111000;
        weights1[30988] <= 16'b0000000000000010;
        weights1[30989] <= 16'b0000000000000100;
        weights1[30990] <= 16'b1111111111110111;
        weights1[30991] <= 16'b0000000000000101;
        weights1[30992] <= 16'b1111111111110111;
        weights1[30993] <= 16'b0000000000000010;
        weights1[30994] <= 16'b0000000000000111;
        weights1[30995] <= 16'b0000000000001001;
        weights1[30996] <= 16'b1111111111010111;
        weights1[30997] <= 16'b1111111111001010;
        weights1[30998] <= 16'b1111111110110001;
        weights1[30999] <= 16'b1111111110101100;
        weights1[31000] <= 16'b1111111110111101;
        weights1[31001] <= 16'b1111111110110100;
        weights1[31002] <= 16'b1111111110110000;
        weights1[31003] <= 16'b1111111110110110;
        weights1[31004] <= 16'b1111111110000100;
        weights1[31005] <= 16'b1111111101110010;
        weights1[31006] <= 16'b1111111110001000;
        weights1[31007] <= 16'b1111111110000110;
        weights1[31008] <= 16'b1111111110001101;
        weights1[31009] <= 16'b1111111110001111;
        weights1[31010] <= 16'b1111111110001111;
        weights1[31011] <= 16'b1111111110101100;
        weights1[31012] <= 16'b1111111110110011;
        weights1[31013] <= 16'b1111111110111111;
        weights1[31014] <= 16'b1111111111001001;
        weights1[31015] <= 16'b1111111111000110;
        weights1[31016] <= 16'b1111111110111100;
        weights1[31017] <= 16'b1111111111011100;
        weights1[31018] <= 16'b1111111111010011;
        weights1[31019] <= 16'b1111111111101001;
        weights1[31020] <= 16'b1111111111011011;
        weights1[31021] <= 16'b1111111111111011;
        weights1[31022] <= 16'b1111111111111001;
        weights1[31023] <= 16'b1111111111111010;
        weights1[31024] <= 16'b1111111111011010;
        weights1[31025] <= 16'b1111111111001000;
        weights1[31026] <= 16'b1111111110111001;
        weights1[31027] <= 16'b1111111110110000;
        weights1[31028] <= 16'b1111111110011001;
        weights1[31029] <= 16'b1111111110000111;
        weights1[31030] <= 16'b1111111101111110;
        weights1[31031] <= 16'b1111111101100111;
        weights1[31032] <= 16'b1111111101110100;
        weights1[31033] <= 16'b1111111101111011;
        weights1[31034] <= 16'b1111111110101100;
        weights1[31035] <= 16'b1111111110110100;
        weights1[31036] <= 16'b1111111110110010;
        weights1[31037] <= 16'b1111111110111000;
        weights1[31038] <= 16'b1111111110111000;
        weights1[31039] <= 16'b1111111110101111;
        weights1[31040] <= 16'b1111111110111000;
        weights1[31041] <= 16'b1111111110111001;
        weights1[31042] <= 16'b1111111110111010;
        weights1[31043] <= 16'b1111111111001001;
        weights1[31044] <= 16'b1111111110101111;
        weights1[31045] <= 16'b1111111111010110;
        weights1[31046] <= 16'b1111111111010001;
        weights1[31047] <= 16'b1111111111001001;
        weights1[31048] <= 16'b1111111111011010;
        weights1[31049] <= 16'b1111111111111011;
        weights1[31050] <= 16'b1111111111101100;
        weights1[31051] <= 16'b1111111111110010;
        weights1[31052] <= 16'b1111111111011110;
        weights1[31053] <= 16'b1111111111000101;
        weights1[31054] <= 16'b1111111111000111;
        weights1[31055] <= 16'b1111111110110011;
        weights1[31056] <= 16'b1111111110011001;
        weights1[31057] <= 16'b1111111110010100;
        weights1[31058] <= 16'b1111111101110101;
        weights1[31059] <= 16'b1111111110011000;
        weights1[31060] <= 16'b1111111111001001;
        weights1[31061] <= 16'b1111111111101011;
        weights1[31062] <= 16'b1111111111101001;
        weights1[31063] <= 16'b1111111111101001;
        weights1[31064] <= 16'b1111111111110001;
        weights1[31065] <= 16'b1111111111100110;
        weights1[31066] <= 16'b1111111111100100;
        weights1[31067] <= 16'b1111111111011100;
        weights1[31068] <= 16'b1111111111011110;
        weights1[31069] <= 16'b1111111111100011;
        weights1[31070] <= 16'b1111111111011100;
        weights1[31071] <= 16'b1111111111010011;
        weights1[31072] <= 16'b1111111111011101;
        weights1[31073] <= 16'b1111111110111000;
        weights1[31074] <= 16'b1111111111100110;
        weights1[31075] <= 16'b1111111111010101;
        weights1[31076] <= 16'b1111111111101000;
        weights1[31077] <= 16'b1111111111101100;
        weights1[31078] <= 16'b1111111111100101;
        weights1[31079] <= 16'b1111111111101101;
        weights1[31080] <= 16'b1111111111100001;
        weights1[31081] <= 16'b1111111111010101;
        weights1[31082] <= 16'b1111111111001001;
        weights1[31083] <= 16'b1111111110110000;
        weights1[31084] <= 16'b1111111111001010;
        weights1[31085] <= 16'b1111111110111001;
        weights1[31086] <= 16'b1111111111011001;
        weights1[31087] <= 16'b1111111111011111;
        weights1[31088] <= 16'b1111111111111010;
        weights1[31089] <= 16'b0000000000000010;
        weights1[31090] <= 16'b0000000000000010;
        weights1[31091] <= 16'b0000000000000000;
        weights1[31092] <= 16'b1111111111111111;
        weights1[31093] <= 16'b1111111111111000;
        weights1[31094] <= 16'b1111111111110011;
        weights1[31095] <= 16'b1111111111110010;
        weights1[31096] <= 16'b1111111111010111;
        weights1[31097] <= 16'b1111111111100100;
        weights1[31098] <= 16'b1111111111011101;
        weights1[31099] <= 16'b1111111111011100;
        weights1[31100] <= 16'b1111111111011011;
        weights1[31101] <= 16'b1111111111100101;
        weights1[31102] <= 16'b1111111111100111;
        weights1[31103] <= 16'b1111111111001011;
        weights1[31104] <= 16'b1111111111100101;
        weights1[31105] <= 16'b1111111111100011;
        weights1[31106] <= 16'b1111111111101011;
        weights1[31107] <= 16'b1111111111110001;
        weights1[31108] <= 16'b1111111111100110;
        weights1[31109] <= 16'b1111111111011110;
        weights1[31110] <= 16'b1111111111010111;
        weights1[31111] <= 16'b1111111111001110;
        weights1[31112] <= 16'b1111111111001111;
        weights1[31113] <= 16'b1111111111101011;
        weights1[31114] <= 16'b1111111111101001;
        weights1[31115] <= 16'b1111111111111000;
        weights1[31116] <= 16'b1111111111101111;
        weights1[31117] <= 16'b1111111111110100;
        weights1[31118] <= 16'b0000000000000001;
        weights1[31119] <= 16'b1111111111111100;
        weights1[31120] <= 16'b1111111111101100;
        weights1[31121] <= 16'b1111111111110001;
        weights1[31122] <= 16'b1111111111110100;
        weights1[31123] <= 16'b1111111111110110;
        weights1[31124] <= 16'b1111111111110001;
        weights1[31125] <= 16'b1111111111101101;
        weights1[31126] <= 16'b1111111111011101;
        weights1[31127] <= 16'b1111111111011011;
        weights1[31128] <= 16'b1111111111100010;
        weights1[31129] <= 16'b1111111111000011;
        weights1[31130] <= 16'b1111111111001110;
        weights1[31131] <= 16'b1111111111011111;
        weights1[31132] <= 16'b1111111111111001;
        weights1[31133] <= 16'b1111111111101001;
        weights1[31134] <= 16'b1111111111100111;
        weights1[31135] <= 16'b1111111111110000;
        weights1[31136] <= 16'b1111111111100101;
        weights1[31137] <= 16'b1111111111101010;
        weights1[31138] <= 16'b1111111111100011;
        weights1[31139] <= 16'b1111111111011001;
        weights1[31140] <= 16'b1111111111011111;
        weights1[31141] <= 16'b1111111111111111;
        weights1[31142] <= 16'b0000000000000111;
        weights1[31143] <= 16'b1111111111111101;
        weights1[31144] <= 16'b1111111111111001;
        weights1[31145] <= 16'b1111111111111100;
        weights1[31146] <= 16'b1111111111111000;
        weights1[31147] <= 16'b1111111111111000;
        weights1[31148] <= 16'b1111111111110101;
        weights1[31149] <= 16'b1111111111111011;
        weights1[31150] <= 16'b1111111111101100;
        weights1[31151] <= 16'b1111111111101010;
        weights1[31152] <= 16'b1111111111110100;
        weights1[31153] <= 16'b1111111111010111;
        weights1[31154] <= 16'b1111111111101011;
        weights1[31155] <= 16'b1111111111010111;
        weights1[31156] <= 16'b1111111111010101;
        weights1[31157] <= 16'b1111111111011010;
        weights1[31158] <= 16'b1111111111011011;
        weights1[31159] <= 16'b1111111111100100;
        weights1[31160] <= 16'b1111111111101101;
        weights1[31161] <= 16'b1111111111110001;
        weights1[31162] <= 16'b1111111111110001;
        weights1[31163] <= 16'b1111111111101111;
        weights1[31164] <= 16'b1111111111110101;
        weights1[31165] <= 16'b1111111111110011;
        weights1[31166] <= 16'b1111111111101111;
        weights1[31167] <= 16'b1111111111100100;
        weights1[31168] <= 16'b1111111111100010;
        weights1[31169] <= 16'b0000000000011010;
        weights1[31170] <= 16'b0000000000000101;
        weights1[31171] <= 16'b1111111111110011;
        weights1[31172] <= 16'b1111111111111101;
        weights1[31173] <= 16'b1111111111100101;
        weights1[31174] <= 16'b0000000000000010;
        weights1[31175] <= 16'b1111111111111111;
        weights1[31176] <= 16'b1111111111101001;
        weights1[31177] <= 16'b1111111111101110;
        weights1[31178] <= 16'b1111111111101100;
        weights1[31179] <= 16'b1111111111101100;
        weights1[31180] <= 16'b1111111111110101;
        weights1[31181] <= 16'b1111111111110001;
        weights1[31182] <= 16'b1111111111100101;
        weights1[31183] <= 16'b1111111111110001;
        weights1[31184] <= 16'b1111111111011110;
        weights1[31185] <= 16'b1111111111110100;
        weights1[31186] <= 16'b1111111111110111;
        weights1[31187] <= 16'b1111111111100100;
        weights1[31188] <= 16'b1111111111101000;
        weights1[31189] <= 16'b1111111111101100;
        weights1[31190] <= 16'b1111111111111001;
        weights1[31191] <= 16'b1111111111110100;
        weights1[31192] <= 16'b1111111111111100;
        weights1[31193] <= 16'b1111111111110100;
        weights1[31194] <= 16'b1111111111111101;
        weights1[31195] <= 16'b1111111111110100;
        weights1[31196] <= 16'b1111111111111111;
        weights1[31197] <= 16'b0000000000000001;
        weights1[31198] <= 16'b1111111111100101;
        weights1[31199] <= 16'b1111111111111011;
        weights1[31200] <= 16'b0000000000101000;
        weights1[31201] <= 16'b0000000000011100;
        weights1[31202] <= 16'b1111111111111100;
        weights1[31203] <= 16'b1111111111101011;
        weights1[31204] <= 16'b0000000000000010;
        weights1[31205] <= 16'b1111111111111101;
        weights1[31206] <= 16'b1111111111111111;
        weights1[31207] <= 16'b0000000000001000;
        weights1[31208] <= 16'b1111111111100111;
        weights1[31209] <= 16'b0000000000000101;
        weights1[31210] <= 16'b1111111111101010;
        weights1[31211] <= 16'b1111111111101011;
        weights1[31212] <= 16'b1111111111101000;
        weights1[31213] <= 16'b1111111111111001;
        weights1[31214] <= 16'b1111111111111010;
        weights1[31215] <= 16'b1111111111101000;
        weights1[31216] <= 16'b1111111111101000;
        weights1[31217] <= 16'b1111111111100110;
        weights1[31218] <= 16'b1111111111110100;
        weights1[31219] <= 16'b1111111111110100;
        weights1[31220] <= 16'b1111111111111000;
        weights1[31221] <= 16'b1111111111110011;
        weights1[31222] <= 16'b1111111111110101;
        weights1[31223] <= 16'b1111111111111110;
        weights1[31224] <= 16'b1111111111110111;
        weights1[31225] <= 16'b0000000000001110;
        weights1[31226] <= 16'b1111111111110101;
        weights1[31227] <= 16'b1111111111110101;
        weights1[31228] <= 16'b1111111111101001;
        weights1[31229] <= 16'b1111111111100100;
        weights1[31230] <= 16'b1111111111011111;
        weights1[31231] <= 16'b1111111111011101;
        weights1[31232] <= 16'b1111111111111111;
        weights1[31233] <= 16'b1111111111101110;
        weights1[31234] <= 16'b1111111111110100;
        weights1[31235] <= 16'b1111111111101010;
        weights1[31236] <= 16'b1111111111110100;
        weights1[31237] <= 16'b1111111111111111;
        weights1[31238] <= 16'b1111111111110000;
        weights1[31239] <= 16'b1111111111101001;
        weights1[31240] <= 16'b1111111111110101;
        weights1[31241] <= 16'b1111111111101101;
        weights1[31242] <= 16'b1111111111101011;
        weights1[31243] <= 16'b1111111111100010;
        weights1[31244] <= 16'b1111111111100101;
        weights1[31245] <= 16'b1111111111101001;
        weights1[31246] <= 16'b1111111111110110;
        weights1[31247] <= 16'b1111111111111001;
        weights1[31248] <= 16'b1111111111111111;
        weights1[31249] <= 16'b1111111111111110;
        weights1[31250] <= 16'b1111111111110111;
        weights1[31251] <= 16'b0000000000000000;
        weights1[31252] <= 16'b1111111111111001;
        weights1[31253] <= 16'b0000000000010010;
        weights1[31254] <= 16'b0000000000001000;
        weights1[31255] <= 16'b0000000000001100;
        weights1[31256] <= 16'b0000000000100000;
        weights1[31257] <= 16'b1111111111101100;
        weights1[31258] <= 16'b0000000000001001;
        weights1[31259] <= 16'b1111111111110110;
        weights1[31260] <= 16'b1111111111101001;
        weights1[31261] <= 16'b1111111111101001;
        weights1[31262] <= 16'b1111111111011010;
        weights1[31263] <= 16'b1111111111010100;
        weights1[31264] <= 16'b0000000000001100;
        weights1[31265] <= 16'b0000000000000101;
        weights1[31266] <= 16'b1111111111110001;
        weights1[31267] <= 16'b1111111111101111;
        weights1[31268] <= 16'b1111111111100011;
        weights1[31269] <= 16'b1111111111110010;
        weights1[31270] <= 16'b1111111111110010;
        weights1[31271] <= 16'b1111111111110000;
        weights1[31272] <= 16'b1111111111100110;
        weights1[31273] <= 16'b1111111111101100;
        weights1[31274] <= 16'b1111111111110111;
        weights1[31275] <= 16'b1111111111111110;
        weights1[31276] <= 16'b0000000000000011;
        weights1[31277] <= 16'b1111111111110110;
        weights1[31278] <= 16'b1111111111111111;
        weights1[31279] <= 16'b1111111111111010;
        weights1[31280] <= 16'b0000000000000010;
        weights1[31281] <= 16'b0000000000001100;
        weights1[31282] <= 16'b0000000000010000;
        weights1[31283] <= 16'b0000000000001000;
        weights1[31284] <= 16'b0000000000001001;
        weights1[31285] <= 16'b1111111111011110;
        weights1[31286] <= 16'b0000000000001100;
        weights1[31287] <= 16'b0000000000101100;
        weights1[31288] <= 16'b0000000000001110;
        weights1[31289] <= 16'b0000000000000101;
        weights1[31290] <= 16'b1111111111111110;
        weights1[31291] <= 16'b0000000000010001;
        weights1[31292] <= 16'b1111111111110010;
        weights1[31293] <= 16'b1111111111001011;
        weights1[31294] <= 16'b1111111111101001;
        weights1[31295] <= 16'b1111111111011001;
        weights1[31296] <= 16'b1111111111100110;
        weights1[31297] <= 16'b1111111111110100;
        weights1[31298] <= 16'b1111111111110001;
        weights1[31299] <= 16'b1111111111101101;
        weights1[31300] <= 16'b1111111111101111;
        weights1[31301] <= 16'b1111111111110110;
        weights1[31302] <= 16'b1111111111111011;
        weights1[31303] <= 16'b1111111111111111;
        weights1[31304] <= 16'b1111111111111101;
        weights1[31305] <= 16'b1111111111111010;
        weights1[31306] <= 16'b0000000000000110;
        weights1[31307] <= 16'b0000000000000100;
        weights1[31308] <= 16'b1111111111111001;
        weights1[31309] <= 16'b0000000000010100;
        weights1[31310] <= 16'b0000000000010111;
        weights1[31311] <= 16'b0000000000000111;
        weights1[31312] <= 16'b0000000000001000;
        weights1[31313] <= 16'b0000000000001010;
        weights1[31314] <= 16'b1111111111110101;
        weights1[31315] <= 16'b1111111111111011;
        weights1[31316] <= 16'b0000000000001000;
        weights1[31317] <= 16'b0000000000000110;
        weights1[31318] <= 16'b0000000000000110;
        weights1[31319] <= 16'b0000000000000010;
        weights1[31320] <= 16'b1111111111101110;
        weights1[31321] <= 16'b1111111111011100;
        weights1[31322] <= 16'b1111111111101000;
        weights1[31323] <= 16'b1111111111011010;
        weights1[31324] <= 16'b1111111111011010;
        weights1[31325] <= 16'b1111111111101000;
        weights1[31326] <= 16'b1111111111110101;
        weights1[31327] <= 16'b1111111111110101;
        weights1[31328] <= 16'b1111111111110111;
        weights1[31329] <= 16'b1111111111111010;
        weights1[31330] <= 16'b1111111111111101;
        weights1[31331] <= 16'b1111111111111111;
        weights1[31332] <= 16'b0000000000000011;
        weights1[31333] <= 16'b0000000000000011;
        weights1[31334] <= 16'b0000000000000000;
        weights1[31335] <= 16'b0000000000001001;
        weights1[31336] <= 16'b0000000000000110;
        weights1[31337] <= 16'b1111111111111101;
        weights1[31338] <= 16'b1111111111111101;
        weights1[31339] <= 16'b0000000000000100;
        weights1[31340] <= 16'b1111111111111100;
        weights1[31341] <= 16'b0000000000010000;
        weights1[31342] <= 16'b0000000000000011;
        weights1[31343] <= 16'b1111111111101000;
        weights1[31344] <= 16'b1111111111101101;
        weights1[31345] <= 16'b1111111111111100;
        weights1[31346] <= 16'b1111111111110100;
        weights1[31347] <= 16'b1111111111101111;
        weights1[31348] <= 16'b1111111111100011;
        weights1[31349] <= 16'b1111111111100011;
        weights1[31350] <= 16'b1111111111001101;
        weights1[31351] <= 16'b1111111111011111;
        weights1[31352] <= 16'b1111111111100010;
        weights1[31353] <= 16'b1111111111100101;
        weights1[31354] <= 16'b1111111111101101;
        weights1[31355] <= 16'b1111111111110101;
        weights1[31356] <= 16'b1111111111110111;
        weights1[31357] <= 16'b1111111111111111;
        weights1[31358] <= 16'b0000000000000000;
        weights1[31359] <= 16'b0000000000000000;
        weights1[31360] <= 16'b0000000000000000;
        weights1[31361] <= 16'b1111111111111111;
        weights1[31362] <= 16'b0000000000000010;
        weights1[31363] <= 16'b1111111111111110;
        weights1[31364] <= 16'b0000000000000001;
        weights1[31365] <= 16'b0000000000000101;
        weights1[31366] <= 16'b0000000000000100;
        weights1[31367] <= 16'b0000000000001011;
        weights1[31368] <= 16'b0000000000010000;
        weights1[31369] <= 16'b0000000000011000;
        weights1[31370] <= 16'b0000000000001010;
        weights1[31371] <= 16'b0000000000010101;
        weights1[31372] <= 16'b0000000000000101;
        weights1[31373] <= 16'b0000000000000011;
        weights1[31374] <= 16'b1111111111111011;
        weights1[31375] <= 16'b1111111111110110;
        weights1[31376] <= 16'b0000000000000011;
        weights1[31377] <= 16'b0000000000000011;
        weights1[31378] <= 16'b1111111111111110;
        weights1[31379] <= 16'b0000000000000001;
        weights1[31380] <= 16'b1111111111111100;
        weights1[31381] <= 16'b0000000000000011;
        weights1[31382] <= 16'b0000000000000110;
        weights1[31383] <= 16'b0000000000000001;
        weights1[31384] <= 16'b0000000000000101;
        weights1[31385] <= 16'b0000000000000010;
        weights1[31386] <= 16'b0000000000000100;
        weights1[31387] <= 16'b0000000000000000;
        weights1[31388] <= 16'b0000000000000000;
        weights1[31389] <= 16'b0000000000000001;
        weights1[31390] <= 16'b1111111111111111;
        weights1[31391] <= 16'b0000000000000010;
        weights1[31392] <= 16'b0000000000001011;
        weights1[31393] <= 16'b0000000000010111;
        weights1[31394] <= 16'b0000000000010011;
        weights1[31395] <= 16'b0000000000010000;
        weights1[31396] <= 16'b0000000000010101;
        weights1[31397] <= 16'b0000000000011110;
        weights1[31398] <= 16'b0000000000010110;
        weights1[31399] <= 16'b0000000000010111;
        weights1[31400] <= 16'b0000000000010001;
        weights1[31401] <= 16'b0000000000010010;
        weights1[31402] <= 16'b0000000000010111;
        weights1[31403] <= 16'b0000000000011011;
        weights1[31404] <= 16'b0000000000001101;
        weights1[31405] <= 16'b0000000000010101;
        weights1[31406] <= 16'b0000000000000111;
        weights1[31407] <= 16'b0000000000000101;
        weights1[31408] <= 16'b0000000000001110;
        weights1[31409] <= 16'b0000000000010000;
        weights1[31410] <= 16'b0000000000001010;
        weights1[31411] <= 16'b0000000000001101;
        weights1[31412] <= 16'b0000000000000000;
        weights1[31413] <= 16'b0000000000000100;
        weights1[31414] <= 16'b0000000000000100;
        weights1[31415] <= 16'b0000000000000010;
        weights1[31416] <= 16'b0000000000000010;
        weights1[31417] <= 16'b0000000000000010;
        weights1[31418] <= 16'b0000000000000111;
        weights1[31419] <= 16'b0000000000001110;
        weights1[31420] <= 16'b0000000000011001;
        weights1[31421] <= 16'b0000000000010101;
        weights1[31422] <= 16'b0000000000011110;
        weights1[31423] <= 16'b0000000000001101;
        weights1[31424] <= 16'b0000000000011000;
        weights1[31425] <= 16'b0000000000011100;
        weights1[31426] <= 16'b0000000000000110;
        weights1[31427] <= 16'b0000000000001110;
        weights1[31428] <= 16'b0000000000011001;
        weights1[31429] <= 16'b0000000000001011;
        weights1[31430] <= 16'b0000000000100100;
        weights1[31431] <= 16'b0000000000010111;
        weights1[31432] <= 16'b0000000000001010;
        weights1[31433] <= 16'b0000000000001110;
        weights1[31434] <= 16'b0000000000100001;
        weights1[31435] <= 16'b0000000000000101;
        weights1[31436] <= 16'b0000000000010111;
        weights1[31437] <= 16'b0000000000011110;
        weights1[31438] <= 16'b0000000000001111;
        weights1[31439] <= 16'b0000000000001011;
        weights1[31440] <= 16'b0000000000001001;
        weights1[31441] <= 16'b0000000000001100;
        weights1[31442] <= 16'b0000000000001011;
        weights1[31443] <= 16'b0000000000001000;
        weights1[31444] <= 16'b0000000000000011;
        weights1[31445] <= 16'b0000000000000100;
        weights1[31446] <= 16'b0000000000001010;
        weights1[31447] <= 16'b0000000000010110;
        weights1[31448] <= 16'b0000000000011011;
        weights1[31449] <= 16'b0000000000011110;
        weights1[31450] <= 16'b0000000000011111;
        weights1[31451] <= 16'b0000000000101011;
        weights1[31452] <= 16'b0000000000100101;
        weights1[31453] <= 16'b0000000000001001;
        weights1[31454] <= 16'b0000000000011101;
        weights1[31455] <= 16'b0000000000001111;
        weights1[31456] <= 16'b0000000000011011;
        weights1[31457] <= 16'b0000000000011010;
        weights1[31458] <= 16'b0000000000010011;
        weights1[31459] <= 16'b1111111111100101;
        weights1[31460] <= 16'b1111111111111001;
        weights1[31461] <= 16'b0000000000010101;
        weights1[31462] <= 16'b1111111111111110;
        weights1[31463] <= 16'b1111111111111101;
        weights1[31464] <= 16'b0000000000100000;
        weights1[31465] <= 16'b0000000000001101;
        weights1[31466] <= 16'b0000000000001011;
        weights1[31467] <= 16'b0000000000010110;
        weights1[31468] <= 16'b0000000000001101;
        weights1[31469] <= 16'b0000000000010010;
        weights1[31470] <= 16'b0000000000010010;
        weights1[31471] <= 16'b0000000000000110;
        weights1[31472] <= 16'b0000000000000000;
        weights1[31473] <= 16'b0000000000001011;
        weights1[31474] <= 16'b0000000000001110;
        weights1[31475] <= 16'b0000000000100000;
        weights1[31476] <= 16'b0000000000011011;
        weights1[31477] <= 16'b0000000000010001;
        weights1[31478] <= 16'b0000000000100001;
        weights1[31479] <= 16'b0000000000100000;
        weights1[31480] <= 16'b0000000000010111;
        weights1[31481] <= 16'b0000000000010101;
        weights1[31482] <= 16'b0000000000100000;
        weights1[31483] <= 16'b0000000000001011;
        weights1[31484] <= 16'b1111111111110100;
        weights1[31485] <= 16'b0000000000000011;
        weights1[31486] <= 16'b0000000000001011;
        weights1[31487] <= 16'b1111111111111001;
        weights1[31488] <= 16'b0000000000001000;
        weights1[31489] <= 16'b1111111111101110;
        weights1[31490] <= 16'b1111111111111111;
        weights1[31491] <= 16'b0000000000010010;
        weights1[31492] <= 16'b0000000000000110;
        weights1[31493] <= 16'b0000000000001000;
        weights1[31494] <= 16'b1111111111111100;
        weights1[31495] <= 16'b0000000000100000;
        weights1[31496] <= 16'b0000000000001111;
        weights1[31497] <= 16'b0000000000010010;
        weights1[31498] <= 16'b0000000000011001;
        weights1[31499] <= 16'b0000000000001100;
        weights1[31500] <= 16'b0000000000000010;
        weights1[31501] <= 16'b0000000000000111;
        weights1[31502] <= 16'b0000000000011010;
        weights1[31503] <= 16'b0000000000101100;
        weights1[31504] <= 16'b0000000000011111;
        weights1[31505] <= 16'b0000000000001110;
        weights1[31506] <= 16'b0000000000010010;
        weights1[31507] <= 16'b0000000000010110;
        weights1[31508] <= 16'b1111111111111010;
        weights1[31509] <= 16'b0000000000000101;
        weights1[31510] <= 16'b1111111111110110;
        weights1[31511] <= 16'b1111111111111101;
        weights1[31512] <= 16'b0000000000011010;
        weights1[31513] <= 16'b0000000000001100;
        weights1[31514] <= 16'b0000000000010111;
        weights1[31515] <= 16'b0000000000111011;
        weights1[31516] <= 16'b0000000000011000;
        weights1[31517] <= 16'b0000000000010010;
        weights1[31518] <= 16'b1111111111110000;
        weights1[31519] <= 16'b0000000000101000;
        weights1[31520] <= 16'b0000000000010010;
        weights1[31521] <= 16'b0000000000000110;
        weights1[31522] <= 16'b1111111111101111;
        weights1[31523] <= 16'b0000000000001110;
        weights1[31524] <= 16'b0000000000011000;
        weights1[31525] <= 16'b0000000000011100;
        weights1[31526] <= 16'b0000000000011100;
        weights1[31527] <= 16'b0000000000011010;
        weights1[31528] <= 16'b0000000000000101;
        weights1[31529] <= 16'b0000000000001011;
        weights1[31530] <= 16'b0000000000011000;
        weights1[31531] <= 16'b0000000000011111;
        weights1[31532] <= 16'b0000000000001111;
        weights1[31533] <= 16'b0000000000011000;
        weights1[31534] <= 16'b0000000000011100;
        weights1[31535] <= 16'b0000000000010110;
        weights1[31536] <= 16'b0000000000000110;
        weights1[31537] <= 16'b0000000000011101;
        weights1[31538] <= 16'b0000000000000011;
        weights1[31539] <= 16'b0000000000000001;
        weights1[31540] <= 16'b1111111111110111;
        weights1[31541] <= 16'b0000000000000010;
        weights1[31542] <= 16'b0000000000001010;
        weights1[31543] <= 16'b0000000000001100;
        weights1[31544] <= 16'b1111111111111001;
        weights1[31545] <= 16'b0000000000001101;
        weights1[31546] <= 16'b0000000000000010;
        weights1[31547] <= 16'b0000000000011001;
        weights1[31548] <= 16'b0000000000000101;
        weights1[31549] <= 16'b1111111111111000;
        weights1[31550] <= 16'b0000000000101010;
        weights1[31551] <= 16'b0000000000101010;
        weights1[31552] <= 16'b0000000000011011;
        weights1[31553] <= 16'b0000000000011011;
        weights1[31554] <= 16'b0000000000100100;
        weights1[31555] <= 16'b0000000000011010;
        weights1[31556] <= 16'b0000000000000100;
        weights1[31557] <= 16'b0000000000010010;
        weights1[31558] <= 16'b0000000000010011;
        weights1[31559] <= 16'b0000000000001100;
        weights1[31560] <= 16'b0000000000010110;
        weights1[31561] <= 16'b0000000000011111;
        weights1[31562] <= 16'b0000000000100000;
        weights1[31563] <= 16'b1111111111110110;
        weights1[31564] <= 16'b0000000000000101;
        weights1[31565] <= 16'b0000000000000101;
        weights1[31566] <= 16'b0000000000001100;
        weights1[31567] <= 16'b0000000000001001;
        weights1[31568] <= 16'b0000000000000101;
        weights1[31569] <= 16'b0000000000001000;
        weights1[31570] <= 16'b1111111111110101;
        weights1[31571] <= 16'b1111111111101000;
        weights1[31572] <= 16'b1111111111110111;
        weights1[31573] <= 16'b1111111111111101;
        weights1[31574] <= 16'b0000000000010101;
        weights1[31575] <= 16'b0000000000011010;
        weights1[31576] <= 16'b1111111111111001;
        weights1[31577] <= 16'b0000000000010001;
        weights1[31578] <= 16'b0000000000011101;
        weights1[31579] <= 16'b0000000000011110;
        weights1[31580] <= 16'b0000000000010111;
        weights1[31581] <= 16'b0000000000110011;
        weights1[31582] <= 16'b0000000000101010;
        weights1[31583] <= 16'b0000000000100110;
        weights1[31584] <= 16'b0000000000000010;
        weights1[31585] <= 16'b0000000000001110;
        weights1[31586] <= 16'b0000000000001111;
        weights1[31587] <= 16'b0000000000001001;
        weights1[31588] <= 16'b0000000000000100;
        weights1[31589] <= 16'b0000000000010101;
        weights1[31590] <= 16'b0000000000011011;
        weights1[31591] <= 16'b0000000000011010;
        weights1[31592] <= 16'b1111111111110110;
        weights1[31593] <= 16'b0000000000010011;
        weights1[31594] <= 16'b0000000000001100;
        weights1[31595] <= 16'b0000000000000000;
        weights1[31596] <= 16'b0000000000001001;
        weights1[31597] <= 16'b0000000000100001;
        weights1[31598] <= 16'b1111111111111000;
        weights1[31599] <= 16'b1111111111110001;
        weights1[31600] <= 16'b1111111111100111;
        weights1[31601] <= 16'b0000000000001000;
        weights1[31602] <= 16'b0000000000100010;
        weights1[31603] <= 16'b0000000000000001;
        weights1[31604] <= 16'b1111111111111110;
        weights1[31605] <= 16'b0000000000011100;
        weights1[31606] <= 16'b0000000000000001;
        weights1[31607] <= 16'b0000000000000011;
        weights1[31608] <= 16'b0000000000011000;
        weights1[31609] <= 16'b0000000000001000;
        weights1[31610] <= 16'b0000000000100100;
        weights1[31611] <= 16'b0000000000100111;
        weights1[31612] <= 16'b0000000000000111;
        weights1[31613] <= 16'b0000000000001110;
        weights1[31614] <= 16'b0000000000001001;
        weights1[31615] <= 16'b0000000000001101;
        weights1[31616] <= 16'b1111111111111110;
        weights1[31617] <= 16'b0000000000001110;
        weights1[31618] <= 16'b0000000000001101;
        weights1[31619] <= 16'b1111111111111011;
        weights1[31620] <= 16'b1111111111110011;
        weights1[31621] <= 16'b0000000000010000;
        weights1[31622] <= 16'b0000000000001100;
        weights1[31623] <= 16'b1111111111110100;
        weights1[31624] <= 16'b1111111111110000;
        weights1[31625] <= 16'b0000000000101010;
        weights1[31626] <= 16'b0000000000001111;
        weights1[31627] <= 16'b0000000000000001;
        weights1[31628] <= 16'b1111111111100100;
        weights1[31629] <= 16'b0000000000010110;
        weights1[31630] <= 16'b0000000000001111;
        weights1[31631] <= 16'b0000000000000011;
        weights1[31632] <= 16'b0000000000000110;
        weights1[31633] <= 16'b1111111111111111;
        weights1[31634] <= 16'b1111111111110000;
        weights1[31635] <= 16'b0000000000001011;
        weights1[31636] <= 16'b1111111111111011;
        weights1[31637] <= 16'b1111111111111111;
        weights1[31638] <= 16'b0000000000100011;
        weights1[31639] <= 16'b0000000000011011;
        weights1[31640] <= 16'b0000000000001000;
        weights1[31641] <= 16'b0000000000010001;
        weights1[31642] <= 16'b0000000000010010;
        weights1[31643] <= 16'b0000000000011010;
        weights1[31644] <= 16'b0000000000011011;
        weights1[31645] <= 16'b1111111111110101;
        weights1[31646] <= 16'b1111111111111111;
        weights1[31647] <= 16'b0000000000001000;
        weights1[31648] <= 16'b0000000000001001;
        weights1[31649] <= 16'b0000000000011011;
        weights1[31650] <= 16'b0000000000000111;
        weights1[31651] <= 16'b1111111111110001;
        weights1[31652] <= 16'b1111111111111010;
        weights1[31653] <= 16'b0000000000010110;
        weights1[31654] <= 16'b0000000000101011;
        weights1[31655] <= 16'b1111111111101110;
        weights1[31656] <= 16'b1111111111101001;
        weights1[31657] <= 16'b0000000000001011;
        weights1[31658] <= 16'b0000000000000011;
        weights1[31659] <= 16'b1111111111101001;
        weights1[31660] <= 16'b0000000000010010;
        weights1[31661] <= 16'b1111111111111100;
        weights1[31662] <= 16'b1111111111111100;
        weights1[31663] <= 16'b0000000000011001;
        weights1[31664] <= 16'b0000000000000010;
        weights1[31665] <= 16'b0000000000000100;
        weights1[31666] <= 16'b0000000000010010;
        weights1[31667] <= 16'b0000000000100001;
        weights1[31668] <= 16'b0000000000000010;
        weights1[31669] <= 16'b0000000000010001;
        weights1[31670] <= 16'b0000000000010010;
        weights1[31671] <= 16'b0000000000000100;
        weights1[31672] <= 16'b1111111111111101;
        weights1[31673] <= 16'b1111111111110111;
        weights1[31674] <= 16'b0000000000001010;
        weights1[31675] <= 16'b1111111111111110;
        weights1[31676] <= 16'b0000000000010001;
        weights1[31677] <= 16'b0000000000010000;
        weights1[31678] <= 16'b0000000000010101;
        weights1[31679] <= 16'b0000000000000010;
        weights1[31680] <= 16'b1111111111111011;
        weights1[31681] <= 16'b0000000000000010;
        weights1[31682] <= 16'b0000000000010001;
        weights1[31683] <= 16'b1111111111101010;
        weights1[31684] <= 16'b1111111111110111;
        weights1[31685] <= 16'b1111111111111111;
        weights1[31686] <= 16'b1111111111111111;
        weights1[31687] <= 16'b1111111111111000;
        weights1[31688] <= 16'b1111111111110010;
        weights1[31689] <= 16'b1111111111110010;
        weights1[31690] <= 16'b0000000000001110;
        weights1[31691] <= 16'b0000000000010000;
        weights1[31692] <= 16'b0000000000011001;
        weights1[31693] <= 16'b0000000000000010;
        weights1[31694] <= 16'b0000000000100001;
        weights1[31695] <= 16'b0000000000100100;
        weights1[31696] <= 16'b0000000000001010;
        weights1[31697] <= 16'b0000000000010110;
        weights1[31698] <= 16'b0000000000011111;
        weights1[31699] <= 16'b0000000000001011;
        weights1[31700] <= 16'b0000000000000110;
        weights1[31701] <= 16'b0000000000001100;
        weights1[31702] <= 16'b0000000000001000;
        weights1[31703] <= 16'b1111111111111011;
        weights1[31704] <= 16'b0000000000001011;
        weights1[31705] <= 16'b0000000000000011;
        weights1[31706] <= 16'b1111111111111001;
        weights1[31707] <= 16'b0000000000000101;
        weights1[31708] <= 16'b0000000000000010;
        weights1[31709] <= 16'b0000000000000110;
        weights1[31710] <= 16'b0000000000000010;
        weights1[31711] <= 16'b1111111111111010;
        weights1[31712] <= 16'b0000000000001000;
        weights1[31713] <= 16'b0000000000001010;
        weights1[31714] <= 16'b1111111111101111;
        weights1[31715] <= 16'b0000000000010010;
        weights1[31716] <= 16'b1111111111111000;
        weights1[31717] <= 16'b0000000000010000;
        weights1[31718] <= 16'b1111111111111010;
        weights1[31719] <= 16'b1111111111111100;
        weights1[31720] <= 16'b0000000000000110;
        weights1[31721] <= 16'b0000000000001010;
        weights1[31722] <= 16'b0000000000100100;
        weights1[31723] <= 16'b0000000000101111;
        weights1[31724] <= 16'b0000000000010000;
        weights1[31725] <= 16'b0000000000011110;
        weights1[31726] <= 16'b0000000000011011;
        weights1[31727] <= 16'b0000000000100001;
        weights1[31728] <= 16'b0000000000011010;
        weights1[31729] <= 16'b1111111111111111;
        weights1[31730] <= 16'b1111111111111111;
        weights1[31731] <= 16'b1111111111111001;
        weights1[31732] <= 16'b0000000000011011;
        weights1[31733] <= 16'b1111111111111000;
        weights1[31734] <= 16'b0000000000011111;
        weights1[31735] <= 16'b0000000000010010;
        weights1[31736] <= 16'b1111111111101110;
        weights1[31737] <= 16'b1111111111111010;
        weights1[31738] <= 16'b1111111111110001;
        weights1[31739] <= 16'b0000000000100000;
        weights1[31740] <= 16'b1111111111101111;
        weights1[31741] <= 16'b1111111111101010;
        weights1[31742] <= 16'b1111111111111111;
        weights1[31743] <= 16'b0000000000010101;
        weights1[31744] <= 16'b0000000000011110;
        weights1[31745] <= 16'b1111111111111110;
        weights1[31746] <= 16'b0000000000000100;
        weights1[31747] <= 16'b1111111111100101;
        weights1[31748] <= 16'b1111111111111001;
        weights1[31749] <= 16'b0000000000001011;
        weights1[31750] <= 16'b0000000000100111;
        weights1[31751] <= 16'b0000000000101111;
        weights1[31752] <= 16'b0000000000010001;
        weights1[31753] <= 16'b0000000000010101;
        weights1[31754] <= 16'b0000000000011001;
        weights1[31755] <= 16'b0000000000011011;
        weights1[31756] <= 16'b0000000000001000;
        weights1[31757] <= 16'b0000000000001001;
        weights1[31758] <= 16'b0000000000000110;
        weights1[31759] <= 16'b0000000000000111;
        weights1[31760] <= 16'b0000000000001101;
        weights1[31761] <= 16'b1111111111111000;
        weights1[31762] <= 16'b0000000000010000;
        weights1[31763] <= 16'b0000000000001101;
        weights1[31764] <= 16'b1111111111111100;
        weights1[31765] <= 16'b1111111111110011;
        weights1[31766] <= 16'b1111111111111101;
        weights1[31767] <= 16'b0000000000010010;
        weights1[31768] <= 16'b0000000000000110;
        weights1[31769] <= 16'b0000000000000110;
        weights1[31770] <= 16'b0000000000000000;
        weights1[31771] <= 16'b1111111111101110;
        weights1[31772] <= 16'b0000000000000011;
        weights1[31773] <= 16'b0000000000000100;
        weights1[31774] <= 16'b1111111111101001;
        weights1[31775] <= 16'b1111111111100111;
        weights1[31776] <= 16'b1111111111110111;
        weights1[31777] <= 16'b0000000000011001;
        weights1[31778] <= 16'b0000000000011100;
        weights1[31779] <= 16'b0000000000111100;
        weights1[31780] <= 16'b0000000000010100;
        weights1[31781] <= 16'b0000000000011011;
        weights1[31782] <= 16'b0000000000010100;
        weights1[31783] <= 16'b0000000000000100;
        weights1[31784] <= 16'b0000000000011000;
        weights1[31785] <= 16'b0000000000001001;
        weights1[31786] <= 16'b0000000000000010;
        weights1[31787] <= 16'b0000000000100001;
        weights1[31788] <= 16'b0000000000001011;
        weights1[31789] <= 16'b0000000000011010;
        weights1[31790] <= 16'b0000000000001110;
        weights1[31791] <= 16'b1111111111111111;
        weights1[31792] <= 16'b1111111111111011;
        weights1[31793] <= 16'b0000000000011010;
        weights1[31794] <= 16'b1111111111111010;
        weights1[31795] <= 16'b1111111111110100;
        weights1[31796] <= 16'b0000000000011000;
        weights1[31797] <= 16'b0000000000000101;
        weights1[31798] <= 16'b1111111111011101;
        weights1[31799] <= 16'b1111111111111101;
        weights1[31800] <= 16'b1111111111011110;
        weights1[31801] <= 16'b0000000000000010;
        weights1[31802] <= 16'b0000000000001100;
        weights1[31803] <= 16'b1111111111111010;
        weights1[31804] <= 16'b0000000000001000;
        weights1[31805] <= 16'b0000000000100101;
        weights1[31806] <= 16'b0000000000101101;
        weights1[31807] <= 16'b0000000000101001;
        weights1[31808] <= 16'b0000000000010000;
        weights1[31809] <= 16'b0000000000010110;
        weights1[31810] <= 16'b0000000000001011;
        weights1[31811] <= 16'b0000000000000010;
        weights1[31812] <= 16'b1111111111111101;
        weights1[31813] <= 16'b1111111111111111;
        weights1[31814] <= 16'b0000000000000101;
        weights1[31815] <= 16'b0000000000001000;
        weights1[31816] <= 16'b0000000000010100;
        weights1[31817] <= 16'b0000000000000101;
        weights1[31818] <= 16'b0000000000000000;
        weights1[31819] <= 16'b0000000000001101;
        weights1[31820] <= 16'b1111111111111100;
        weights1[31821] <= 16'b0000000000000100;
        weights1[31822] <= 16'b1111111111111100;
        weights1[31823] <= 16'b1111111111101010;
        weights1[31824] <= 16'b1111111111101110;
        weights1[31825] <= 16'b0000000000011010;
        weights1[31826] <= 16'b0000000000001101;
        weights1[31827] <= 16'b1111111111111001;
        weights1[31828] <= 16'b0000000000000000;
        weights1[31829] <= 16'b1111111111110000;
        weights1[31830] <= 16'b0000000000000011;
        weights1[31831] <= 16'b0000000000010010;
        weights1[31832] <= 16'b0000000000001110;
        weights1[31833] <= 16'b0000000000011111;
        weights1[31834] <= 16'b0000000000110100;
        weights1[31835] <= 16'b0000000000100110;
        weights1[31836] <= 16'b0000000000001101;
        weights1[31837] <= 16'b0000000000001001;
        weights1[31838] <= 16'b1111111111111010;
        weights1[31839] <= 16'b1111111111111001;
        weights1[31840] <= 16'b1111111111110111;
        weights1[31841] <= 16'b0000000000010111;
        weights1[31842] <= 16'b0000000000000011;
        weights1[31843] <= 16'b0000000000000010;
        weights1[31844] <= 16'b1111111111111001;
        weights1[31845] <= 16'b0000000000000101;
        weights1[31846] <= 16'b1111111111111110;
        weights1[31847] <= 16'b0000000000000101;
        weights1[31848] <= 16'b0000000000001111;
        weights1[31849] <= 16'b1111111111111100;
        weights1[31850] <= 16'b0000000000000101;
        weights1[31851] <= 16'b1111111111010111;
        weights1[31852] <= 16'b0000000000010101;
        weights1[31853] <= 16'b0000000000010100;
        weights1[31854] <= 16'b0000000000001001;
        weights1[31855] <= 16'b0000000000001011;
        weights1[31856] <= 16'b0000000000001101;
        weights1[31857] <= 16'b0000000000000110;
        weights1[31858] <= 16'b0000000000001101;
        weights1[31859] <= 16'b0000000000010000;
        weights1[31860] <= 16'b0000000000010110;
        weights1[31861] <= 16'b0000000000010110;
        weights1[31862] <= 16'b0000000000100010;
        weights1[31863] <= 16'b0000000000100001;
        weights1[31864] <= 16'b1111111111111110;
        weights1[31865] <= 16'b0000000000000111;
        weights1[31866] <= 16'b0000000000000101;
        weights1[31867] <= 16'b0000000000000101;
        weights1[31868] <= 16'b1111111111111100;
        weights1[31869] <= 16'b0000000000001110;
        weights1[31870] <= 16'b1111111111111110;
        weights1[31871] <= 16'b0000000000010101;
        weights1[31872] <= 16'b0000000000000011;
        weights1[31873] <= 16'b0000000000000010;
        weights1[31874] <= 16'b0000000000001110;
        weights1[31875] <= 16'b0000000000001010;
        weights1[31876] <= 16'b1111111111111000;
        weights1[31877] <= 16'b0000000000100011;
        weights1[31878] <= 16'b0000000000011100;
        weights1[31879] <= 16'b0000000000000110;
        weights1[31880] <= 16'b1111111111111000;
        weights1[31881] <= 16'b0000000000001001;
        weights1[31882] <= 16'b0000000000000110;
        weights1[31883] <= 16'b0000000000001101;
        weights1[31884] <= 16'b0000000000011111;
        weights1[31885] <= 16'b0000000000001001;
        weights1[31886] <= 16'b0000000000100011;
        weights1[31887] <= 16'b0000000000011111;
        weights1[31888] <= 16'b0000000000011111;
        weights1[31889] <= 16'b0000000000011111;
        weights1[31890] <= 16'b0000000000101001;
        weights1[31891] <= 16'b0000000000010110;
        weights1[31892] <= 16'b0000000000000111;
        weights1[31893] <= 16'b0000000000001001;
        weights1[31894] <= 16'b0000000000000110;
        weights1[31895] <= 16'b0000000000000000;
        weights1[31896] <= 16'b0000000000000001;
        weights1[31897] <= 16'b0000000000001110;
        weights1[31898] <= 16'b0000000000010011;
        weights1[31899] <= 16'b0000000000011110;
        weights1[31900] <= 16'b0000000000001001;
        weights1[31901] <= 16'b1111111111110000;
        weights1[31902] <= 16'b0000000000001110;
        weights1[31903] <= 16'b0000000000000011;
        weights1[31904] <= 16'b1111111111111100;
        weights1[31905] <= 16'b1111111111111010;
        weights1[31906] <= 16'b1111111111111011;
        weights1[31907] <= 16'b0000000000010000;
        weights1[31908] <= 16'b0000000000000111;
        weights1[31909] <= 16'b1111111111110100;
        weights1[31910] <= 16'b1111111111111111;
        weights1[31911] <= 16'b0000000000100011;
        weights1[31912] <= 16'b0000000000010100;
        weights1[31913] <= 16'b0000000000011010;
        weights1[31914] <= 16'b0000000000101101;
        weights1[31915] <= 16'b0000000000110001;
        weights1[31916] <= 16'b0000000000010001;
        weights1[31917] <= 16'b0000000000101000;
        weights1[31918] <= 16'b0000000000100101;
        weights1[31919] <= 16'b0000000000100000;
        weights1[31920] <= 16'b0000000000011001;
        weights1[31921] <= 16'b0000000000001111;
        weights1[31922] <= 16'b0000000000010100;
        weights1[31923] <= 16'b0000000000011001;
        weights1[31924] <= 16'b0000000000011110;
        weights1[31925] <= 16'b0000000000010110;
        weights1[31926] <= 16'b0000000000011010;
        weights1[31927] <= 16'b0000000000100000;
        weights1[31928] <= 16'b0000000000001001;
        weights1[31929] <= 16'b1111111111111000;
        weights1[31930] <= 16'b0000000000111100;
        weights1[31931] <= 16'b1111111111101011;
        weights1[31932] <= 16'b0000000000000110;
        weights1[31933] <= 16'b1111111111111000;
        weights1[31934] <= 16'b1111111111101011;
        weights1[31935] <= 16'b0000000000011011;
        weights1[31936] <= 16'b0000000000011010;
        weights1[31937] <= 16'b1111111111101100;
        weights1[31938] <= 16'b0000000000001010;
        weights1[31939] <= 16'b0000000000001111;
        weights1[31940] <= 16'b0000000000000000;
        weights1[31941] <= 16'b0000000000101000;
        weights1[31942] <= 16'b0000000000101001;
        weights1[31943] <= 16'b0000000000101010;
        weights1[31944] <= 16'b0000000000011011;
        weights1[31945] <= 16'b0000000000100100;
        weights1[31946] <= 16'b0000000000011111;
        weights1[31947] <= 16'b0000000000100000;
        weights1[31948] <= 16'b0000000000010010;
        weights1[31949] <= 16'b0000000000010001;
        weights1[31950] <= 16'b0000000000001010;
        weights1[31951] <= 16'b0000000000000111;
        weights1[31952] <= 16'b0000000000000011;
        weights1[31953] <= 16'b0000000000011000;
        weights1[31954] <= 16'b1111111111111100;
        weights1[31955] <= 16'b0000000000011000;
        weights1[31956] <= 16'b0000000000001000;
        weights1[31957] <= 16'b0000000000011111;
        weights1[31958] <= 16'b1111111111110111;
        weights1[31959] <= 16'b0000000000010011;
        weights1[31960] <= 16'b0000000000010101;
        weights1[31961] <= 16'b1111111111101001;
        weights1[31962] <= 16'b1111111111011111;
        weights1[31963] <= 16'b0000000000101001;
        weights1[31964] <= 16'b0000000000010110;
        weights1[31965] <= 16'b1111111111101001;
        weights1[31966] <= 16'b0000000000001010;
        weights1[31967] <= 16'b0000000000101010;
        weights1[31968] <= 16'b0000000000011011;
        weights1[31969] <= 16'b0000000000001110;
        weights1[31970] <= 16'b0000000000011010;
        weights1[31971] <= 16'b0000000000101010;
        weights1[31972] <= 16'b0000000000011010;
        weights1[31973] <= 16'b0000000000101001;
        weights1[31974] <= 16'b0000000000011101;
        weights1[31975] <= 16'b0000000000011110;
        weights1[31976] <= 16'b0000000000011001;
        weights1[31977] <= 16'b0000000000011111;
        weights1[31978] <= 16'b0000000000010100;
        weights1[31979] <= 16'b0000000000001111;
        weights1[31980] <= 16'b1111111111111101;
        weights1[31981] <= 16'b0000000000010101;
        weights1[31982] <= 16'b0000000000001010;
        weights1[31983] <= 16'b0000000000010000;
        weights1[31984] <= 16'b0000000000000101;
        weights1[31985] <= 16'b0000000000010111;
        weights1[31986] <= 16'b1111111111110100;
        weights1[31987] <= 16'b0000000000001111;
        weights1[31988] <= 16'b0000000001000111;
        weights1[31989] <= 16'b0000000000011100;
        weights1[31990] <= 16'b1111111111111000;
        weights1[31991] <= 16'b0000000000110100;
        weights1[31992] <= 16'b0000000000010000;
        weights1[31993] <= 16'b1111111111011110;
        weights1[31994] <= 16'b0000000000010110;
        weights1[31995] <= 16'b0000000000011111;
        weights1[31996] <= 16'b0000000000011011;
        weights1[31997] <= 16'b0000000000011011;
        weights1[31998] <= 16'b0000000000001001;
        weights1[31999] <= 16'b0000000000100101;
        weights1[32000] <= 16'b0000000000101100;
        weights1[32001] <= 16'b0000000000101100;
        weights1[32002] <= 16'b0000000000011010;
        weights1[32003] <= 16'b0000000000010001;
        weights1[32004] <= 16'b0000000000010100;
        weights1[32005] <= 16'b0000000000010110;
        weights1[32006] <= 16'b0000000000011010;
        weights1[32007] <= 16'b0000000000011100;
        weights1[32008] <= 16'b0000000000010100;
        weights1[32009] <= 16'b0000000000010010;
        weights1[32010] <= 16'b0000000000011111;
        weights1[32011] <= 16'b1111111111111100;
        weights1[32012] <= 16'b0000000000011011;
        weights1[32013] <= 16'b0000000000000010;
        weights1[32014] <= 16'b1111111111111111;
        weights1[32015] <= 16'b0000000000010111;
        weights1[32016] <= 16'b0000000000110001;
        weights1[32017] <= 16'b0000000000101100;
        weights1[32018] <= 16'b0000000000001100;
        weights1[32019] <= 16'b0000000000010001;
        weights1[32020] <= 16'b0000000000100111;
        weights1[32021] <= 16'b1111111111111110;
        weights1[32022] <= 16'b0000000000001110;
        weights1[32023] <= 16'b0000000000101010;
        weights1[32024] <= 16'b0000000000001010;
        weights1[32025] <= 16'b1111111111111100;
        weights1[32026] <= 16'b0000000000000101;
        weights1[32027] <= 16'b0000000000100011;
        weights1[32028] <= 16'b0000000000011001;
        weights1[32029] <= 16'b0000000000011111;
        weights1[32030] <= 16'b0000000000001100;
        weights1[32031] <= 16'b0000000000010000;
        weights1[32032] <= 16'b0000000000001100;
        weights1[32033] <= 16'b0000000000001101;
        weights1[32034] <= 16'b0000000000001110;
        weights1[32035] <= 16'b0000000000010011;
        weights1[32036] <= 16'b0000000000010000;
        weights1[32037] <= 16'b0000000000001110;
        weights1[32038] <= 16'b1111111111110101;
        weights1[32039] <= 16'b1111111111111111;
        weights1[32040] <= 16'b0000000000000111;
        weights1[32041] <= 16'b1111111111110011;
        weights1[32042] <= 16'b0000000000000011;
        weights1[32043] <= 16'b0000000000011001;
        weights1[32044] <= 16'b0000000000000000;
        weights1[32045] <= 16'b1111111111111110;
        weights1[32046] <= 16'b0000000000000100;
        weights1[32047] <= 16'b0000000000001000;
        weights1[32048] <= 16'b0000000000001101;
        weights1[32049] <= 16'b1111111111101000;
        weights1[32050] <= 16'b0000000000010000;
        weights1[32051] <= 16'b0000000000010010;
        weights1[32052] <= 16'b0000000000000010;
        weights1[32053] <= 16'b1111111111111011;
        weights1[32054] <= 16'b0000000000000001;
        weights1[32055] <= 16'b0000000000001101;
        weights1[32056] <= 16'b0000000000010101;
        weights1[32057] <= 16'b0000000000100000;
        weights1[32058] <= 16'b0000000000010010;
        weights1[32059] <= 16'b0000000000000101;
        weights1[32060] <= 16'b0000000000000101;
        weights1[32061] <= 16'b0000000000001101;
        weights1[32062] <= 16'b0000000000000100;
        weights1[32063] <= 16'b0000000000010001;
        weights1[32064] <= 16'b0000000000001100;
        weights1[32065] <= 16'b0000000000001111;
        weights1[32066] <= 16'b0000000000001001;
        weights1[32067] <= 16'b0000000000001011;
        weights1[32068] <= 16'b0000000000001101;
        weights1[32069] <= 16'b0000000000010001;
        weights1[32070] <= 16'b0000000000011011;
        weights1[32071] <= 16'b0000000000001010;
        weights1[32072] <= 16'b1111111111101001;
        weights1[32073] <= 16'b1111111111011011;
        weights1[32074] <= 16'b1111111111110111;
        weights1[32075] <= 16'b0000000000000100;
        weights1[32076] <= 16'b1111111111111010;
        weights1[32077] <= 16'b0000000000000001;
        weights1[32078] <= 16'b0000000000001110;
        weights1[32079] <= 16'b0000000000001011;
        weights1[32080] <= 16'b0000000000001111;
        weights1[32081] <= 16'b1111111111110100;
        weights1[32082] <= 16'b0000000000000010;
        weights1[32083] <= 16'b0000000000010010;
        weights1[32084] <= 16'b0000000000010011;
        weights1[32085] <= 16'b0000000000010111;
        weights1[32086] <= 16'b0000000000010001;
        weights1[32087] <= 16'b0000000000000110;
        weights1[32088] <= 16'b0000000000000010;
        weights1[32089] <= 16'b0000000000000110;
        weights1[32090] <= 16'b0000000000000100;
        weights1[32091] <= 16'b1111111111111110;
        weights1[32092] <= 16'b0000000000000111;
        weights1[32093] <= 16'b0000000000001010;
        weights1[32094] <= 16'b0000000000000111;
        weights1[32095] <= 16'b0000000000011000;
        weights1[32096] <= 16'b0000000000011100;
        weights1[32097] <= 16'b0000000000011011;
        weights1[32098] <= 16'b0000000000001011;
        weights1[32099] <= 16'b0000000000011100;
        weights1[32100] <= 16'b0000000000001111;
        weights1[32101] <= 16'b0000000000001001;
        weights1[32102] <= 16'b0000000000100000;
        weights1[32103] <= 16'b0000000000011101;
        weights1[32104] <= 16'b0000000000010101;
        weights1[32105] <= 16'b0000000000011111;
        weights1[32106] <= 16'b0000000000011010;
        weights1[32107] <= 16'b0000000000010111;
        weights1[32108] <= 16'b0000000000000101;
        weights1[32109] <= 16'b0000000000010001;
        weights1[32110] <= 16'b0000000000010010;
        weights1[32111] <= 16'b0000000000010000;
        weights1[32112] <= 16'b0000000000010101;
        weights1[32113] <= 16'b0000000000001111;
        weights1[32114] <= 16'b0000000000000100;
        weights1[32115] <= 16'b1111111111111111;
        weights1[32116] <= 16'b0000000000000010;
        weights1[32117] <= 16'b1111111111111111;
        weights1[32118] <= 16'b0000000000000011;
        weights1[32119] <= 16'b1111111111111110;
        weights1[32120] <= 16'b0000000000000001;
        weights1[32121] <= 16'b0000000000001011;
        weights1[32122] <= 16'b0000000000001010;
        weights1[32123] <= 16'b0000000000010011;
        weights1[32124] <= 16'b0000000000010100;
        weights1[32125] <= 16'b0000000000010001;
        weights1[32126] <= 16'b0000000000001001;
        weights1[32127] <= 16'b0000000000100111;
        weights1[32128] <= 16'b0000000000011110;
        weights1[32129] <= 16'b0000000000011111;
        weights1[32130] <= 16'b0000000000100110;
        weights1[32131] <= 16'b0000000000100010;
        weights1[32132] <= 16'b0000000000000111;
        weights1[32133] <= 16'b0000000000010110;
        weights1[32134] <= 16'b0000000000010000;
        weights1[32135] <= 16'b0000000000001110;
        weights1[32136] <= 16'b0000000000001001;
        weights1[32137] <= 16'b0000000000010000;
        weights1[32138] <= 16'b0000000000001100;
        weights1[32139] <= 16'b0000000000010001;
        weights1[32140] <= 16'b0000000000001100;
        weights1[32141] <= 16'b0000000000000110;
        weights1[32142] <= 16'b0000000000000000;
        weights1[32143] <= 16'b1111111111111100;
        weights1[32144] <= 16'b0000000000000000;
        weights1[32145] <= 16'b0000000000000000;
        weights1[32146] <= 16'b1111111111111111;
        weights1[32147] <= 16'b1111111111111110;
        weights1[32148] <= 16'b1111111111111111;
        weights1[32149] <= 16'b1111111111111110;
        weights1[32150] <= 16'b1111111111111010;
        weights1[32151] <= 16'b1111111111110100;
        weights1[32152] <= 16'b1111111111100011;
        weights1[32153] <= 16'b1111111111100110;
        weights1[32154] <= 16'b1111111111100100;
        weights1[32155] <= 16'b1111111111010001;
        weights1[32156] <= 16'b1111111111001010;
        weights1[32157] <= 16'b1111111111001011;
        weights1[32158] <= 16'b1111111111010101;
        weights1[32159] <= 16'b1111111111001010;
        weights1[32160] <= 16'b1111111111001010;
        weights1[32161] <= 16'b1111111111010100;
        weights1[32162] <= 16'b1111111111011011;
        weights1[32163] <= 16'b1111111111100101;
        weights1[32164] <= 16'b1111111111100100;
        weights1[32165] <= 16'b1111111111110110;
        weights1[32166] <= 16'b1111111111110110;
        weights1[32167] <= 16'b1111111111111011;
        weights1[32168] <= 16'b0000000000000010;
        weights1[32169] <= 16'b0000000000000110;
        weights1[32170] <= 16'b0000000000000000;
        weights1[32171] <= 16'b0000000000000000;
        weights1[32172] <= 16'b0000000000000000;
        weights1[32173] <= 16'b0000000000000000;
        weights1[32174] <= 16'b1111111111111100;
        weights1[32175] <= 16'b1111111111111110;
        weights1[32176] <= 16'b1111111111111100;
        weights1[32177] <= 16'b1111111111111000;
        weights1[32178] <= 16'b1111111111111010;
        weights1[32179] <= 16'b1111111111110000;
        weights1[32180] <= 16'b1111111111011011;
        weights1[32181] <= 16'b1111111111010111;
        weights1[32182] <= 16'b1111111111011011;
        weights1[32183] <= 16'b1111111111100100;
        weights1[32184] <= 16'b1111111111100100;
        weights1[32185] <= 16'b1111111111100100;
        weights1[32186] <= 16'b1111111111100100;
        weights1[32187] <= 16'b1111111111010101;
        weights1[32188] <= 16'b1111111111100010;
        weights1[32189] <= 16'b1111111111100000;
        weights1[32190] <= 16'b1111111111100111;
        weights1[32191] <= 16'b1111111111111000;
        weights1[32192] <= 16'b1111111111110100;
        weights1[32193] <= 16'b0000000000000010;
        weights1[32194] <= 16'b0000000000000011;
        weights1[32195] <= 16'b0000000000000110;
        weights1[32196] <= 16'b0000000000000001;
        weights1[32197] <= 16'b0000000000000101;
        weights1[32198] <= 16'b0000000000000010;
        weights1[32199] <= 16'b0000000000000000;
        weights1[32200] <= 16'b0000000000000010;
        weights1[32201] <= 16'b0000000000000001;
        weights1[32202] <= 16'b1111111111111001;
        weights1[32203] <= 16'b1111111111111011;
        weights1[32204] <= 16'b0000000000000011;
        weights1[32205] <= 16'b0000000000000010;
        weights1[32206] <= 16'b1111111111111001;
        weights1[32207] <= 16'b1111111111111000;
        weights1[32208] <= 16'b1111111111101001;
        weights1[32209] <= 16'b1111111111101011;
        weights1[32210] <= 16'b1111111111101111;
        weights1[32211] <= 16'b0000000000000010;
        weights1[32212] <= 16'b1111111111100101;
        weights1[32213] <= 16'b1111111111110010;
        weights1[32214] <= 16'b1111111111110010;
        weights1[32215] <= 16'b1111111111111111;
        weights1[32216] <= 16'b0000000000000011;
        weights1[32217] <= 16'b0000000000000000;
        weights1[32218] <= 16'b0000000000000110;
        weights1[32219] <= 16'b1111111111110110;
        weights1[32220] <= 16'b0000000000000111;
        weights1[32221] <= 16'b0000000000000011;
        weights1[32222] <= 16'b1111111111111101;
        weights1[32223] <= 16'b1111111111111010;
        weights1[32224] <= 16'b0000000000000110;
        weights1[32225] <= 16'b1111111111111101;
        weights1[32226] <= 16'b1111111111111001;
        weights1[32227] <= 16'b1111111111111010;
        weights1[32228] <= 16'b0000000000000010;
        weights1[32229] <= 16'b1111111111111101;
        weights1[32230] <= 16'b1111111111111000;
        weights1[32231] <= 16'b0000000000000000;
        weights1[32232] <= 16'b0000000000001010;
        weights1[32233] <= 16'b0000000000001101;
        weights1[32234] <= 16'b0000000000001011;
        weights1[32235] <= 16'b0000000000000110;
        weights1[32236] <= 16'b0000000000000001;
        weights1[32237] <= 16'b0000000000000111;
        weights1[32238] <= 16'b0000000000000111;
        weights1[32239] <= 16'b1111111111111110;
        weights1[32240] <= 16'b1111111111110110;
        weights1[32241] <= 16'b0000000000010010;
        weights1[32242] <= 16'b0000000000001111;
        weights1[32243] <= 16'b1111111111110100;
        weights1[32244] <= 16'b0000000000000000;
        weights1[32245] <= 16'b0000000000000000;
        weights1[32246] <= 16'b1111111111110011;
        weights1[32247] <= 16'b1111111111101001;
        weights1[32248] <= 16'b1111111111111001;
        weights1[32249] <= 16'b0000000000000111;
        weights1[32250] <= 16'b1111111111100010;
        weights1[32251] <= 16'b1111111111101101;
        weights1[32252] <= 16'b0000000000000011;
        weights1[32253] <= 16'b1111111111111011;
        weights1[32254] <= 16'b1111111111111010;
        weights1[32255] <= 16'b1111111111111100;
        weights1[32256] <= 16'b0000000000000001;
        weights1[32257] <= 16'b0000000000000000;
        weights1[32258] <= 16'b1111111111111101;
        weights1[32259] <= 16'b0000000000000011;
        weights1[32260] <= 16'b0000000000010000;
        weights1[32261] <= 16'b0000000000010100;
        weights1[32262] <= 16'b0000000000010101;
        weights1[32263] <= 16'b0000000000001110;
        weights1[32264] <= 16'b0000000000001011;
        weights1[32265] <= 16'b0000000000010011;
        weights1[32266] <= 16'b0000000000000111;
        weights1[32267] <= 16'b0000000000011000;
        weights1[32268] <= 16'b0000000000010100;
        weights1[32269] <= 16'b0000000000001101;
        weights1[32270] <= 16'b0000000000011011;
        weights1[32271] <= 16'b0000000000011011;
        weights1[32272] <= 16'b0000000000001011;
        weights1[32273] <= 16'b0000000000000100;
        weights1[32274] <= 16'b0000000000001100;
        weights1[32275] <= 16'b0000000000001111;
        weights1[32276] <= 16'b1111111111100100;
        weights1[32277] <= 16'b1111111111110110;
        weights1[32278] <= 16'b1111111111101011;
        weights1[32279] <= 16'b1111111111101010;
        weights1[32280] <= 16'b0000000000001011;
        weights1[32281] <= 16'b1111111111111000;
        weights1[32282] <= 16'b1111111111111001;
        weights1[32283] <= 16'b0000000000000000;
        weights1[32284] <= 16'b0000000000000010;
        weights1[32285] <= 16'b0000000000001000;
        weights1[32286] <= 16'b0000000000001011;
        weights1[32287] <= 16'b1111111111111111;
        weights1[32288] <= 16'b0000000000000101;
        weights1[32289] <= 16'b0000000000101101;
        weights1[32290] <= 16'b0000000000011010;
        weights1[32291] <= 16'b0000000000010011;
        weights1[32292] <= 16'b1111111111110000;
        weights1[32293] <= 16'b0000000000010011;
        weights1[32294] <= 16'b1111111111101111;
        weights1[32295] <= 16'b0000000000010111;
        weights1[32296] <= 16'b0000000000100011;
        weights1[32297] <= 16'b0000000000010011;
        weights1[32298] <= 16'b0000000000000001;
        weights1[32299] <= 16'b1111111111111011;
        weights1[32300] <= 16'b0000000000001100;
        weights1[32301] <= 16'b0000000000000100;
        weights1[32302] <= 16'b1111111111111000;
        weights1[32303] <= 16'b1111111111110110;
        weights1[32304] <= 16'b0000000000011010;
        weights1[32305] <= 16'b0000000000001001;
        weights1[32306] <= 16'b0000000000010000;
        weights1[32307] <= 16'b0000000000101100;
        weights1[32308] <= 16'b0000000000010111;
        weights1[32309] <= 16'b0000000000000010;
        weights1[32310] <= 16'b1111111111111110;
        weights1[32311] <= 16'b1111111111111010;
        weights1[32312] <= 16'b0000000000000000;
        weights1[32313] <= 16'b1111111111111001;
        weights1[32314] <= 16'b0000000000000011;
        weights1[32315] <= 16'b0000000000000010;
        weights1[32316] <= 16'b1111111111111010;
        weights1[32317] <= 16'b0000000000011101;
        weights1[32318] <= 16'b0000000000010001;
        weights1[32319] <= 16'b0000000000011110;
        weights1[32320] <= 16'b0000000000001111;
        weights1[32321] <= 16'b1111111111111000;
        weights1[32322] <= 16'b0000000000100011;
        weights1[32323] <= 16'b0000000000100001;
        weights1[32324] <= 16'b0000000000010110;
        weights1[32325] <= 16'b0000000000001100;
        weights1[32326] <= 16'b0000000000001000;
        weights1[32327] <= 16'b0000000000001011;
        weights1[32328] <= 16'b0000000000000111;
        weights1[32329] <= 16'b0000000000100011;
        weights1[32330] <= 16'b0000000000011100;
        weights1[32331] <= 16'b0000000000011100;
        weights1[32332] <= 16'b0000000000011000;
        weights1[32333] <= 16'b0000000000011100;
        weights1[32334] <= 16'b0000000000010110;
        weights1[32335] <= 16'b0000000000010001;
        weights1[32336] <= 16'b0000000000000001;
        weights1[32337] <= 16'b0000000000000101;
        weights1[32338] <= 16'b0000000000000111;
        weights1[32339] <= 16'b0000000000000100;
        weights1[32340] <= 16'b1111111111111111;
        weights1[32341] <= 16'b1111111111110011;
        weights1[32342] <= 16'b1111111111110000;
        weights1[32343] <= 16'b1111111111111110;
        weights1[32344] <= 16'b0000000000010100;
        weights1[32345] <= 16'b0000000000011111;
        weights1[32346] <= 16'b0000000000010100;
        weights1[32347] <= 16'b1111111111111100;
        weights1[32348] <= 16'b1111111111111111;
        weights1[32349] <= 16'b1111111111111010;
        weights1[32350] <= 16'b0000000000000010;
        weights1[32351] <= 16'b0000000000010100;
        weights1[32352] <= 16'b1111111111101011;
        weights1[32353] <= 16'b0000000000001110;
        weights1[32354] <= 16'b0000000000001010;
        weights1[32355] <= 16'b0000000000100110;
        weights1[32356] <= 16'b0000000000101101;
        weights1[32357] <= 16'b0000000000101000;
        weights1[32358] <= 16'b0000000000010110;
        weights1[32359] <= 16'b0000000000110011;
        weights1[32360] <= 16'b0000000000001100;
        weights1[32361] <= 16'b0000000000010000;
        weights1[32362] <= 16'b1111111111111000;
        weights1[32363] <= 16'b0000000000010111;
        weights1[32364] <= 16'b0000000000100011;
        weights1[32365] <= 16'b0000000000101000;
        weights1[32366] <= 16'b0000000000010111;
        weights1[32367] <= 16'b0000000000001011;
        weights1[32368] <= 16'b1111111111110110;
        weights1[32369] <= 16'b1111111111110000;
        weights1[32370] <= 16'b1111111111110010;
        weights1[32371] <= 16'b0000000000000001;
        weights1[32372] <= 16'b0000000000000100;
        weights1[32373] <= 16'b0000000000101001;
        weights1[32374] <= 16'b0000000000110100;
        weights1[32375] <= 16'b1111111111111000;
        weights1[32376] <= 16'b1111111111110001;
        weights1[32377] <= 16'b0000000000000010;
        weights1[32378] <= 16'b1111111111110000;
        weights1[32379] <= 16'b1111111111111101;
        weights1[32380] <= 16'b0000000000010101;
        weights1[32381] <= 16'b0000000000100010;
        weights1[32382] <= 16'b0000000000011010;
        weights1[32383] <= 16'b0000000000101100;
        weights1[32384] <= 16'b0000000000011001;
        weights1[32385] <= 16'b0000000000000001;
        weights1[32386] <= 16'b0000000000100110;
        weights1[32387] <= 16'b0000000000001110;
        weights1[32388] <= 16'b0000000000001011;
        weights1[32389] <= 16'b0000000000000000;
        weights1[32390] <= 16'b0000000000010011;
        weights1[32391] <= 16'b0000000000110001;
        weights1[32392] <= 16'b0000000000111101;
        weights1[32393] <= 16'b0000000000110001;
        weights1[32394] <= 16'b0000000000011000;
        weights1[32395] <= 16'b0000000000000101;
        weights1[32396] <= 16'b1111111111110101;
        weights1[32397] <= 16'b1111111111101011;
        weights1[32398] <= 16'b1111111111110000;
        weights1[32399] <= 16'b0000000000000101;
        weights1[32400] <= 16'b0000000000011100;
        weights1[32401] <= 16'b0000000000111001;
        weights1[32402] <= 16'b0000000000111011;
        weights1[32403] <= 16'b0000000000011101;
        weights1[32404] <= 16'b0000000000100011;
        weights1[32405] <= 16'b0000000000010011;
        weights1[32406] <= 16'b0000000000000011;
        weights1[32407] <= 16'b1111111111110011;
        weights1[32408] <= 16'b1111111111011010;
        weights1[32409] <= 16'b1111111111110000;
        weights1[32410] <= 16'b1111111111100101;
        weights1[32411] <= 16'b1111111111101011;
        weights1[32412] <= 16'b1111111111101000;
        weights1[32413] <= 16'b1111111111111010;
        weights1[32414] <= 16'b1111111111111001;
        weights1[32415] <= 16'b1111111111110100;
        weights1[32416] <= 16'b0000000000010100;
        weights1[32417] <= 16'b0000000000100001;
        weights1[32418] <= 16'b0000000000100101;
        weights1[32419] <= 16'b0000000000111110;
        weights1[32420] <= 16'b0000000000110111;
        weights1[32421] <= 16'b0000000000001100;
        weights1[32422] <= 16'b0000000000001010;
        weights1[32423] <= 16'b1111111111111010;
        weights1[32424] <= 16'b1111111111110110;
        weights1[32425] <= 16'b1111111111110011;
        weights1[32426] <= 16'b1111111111100011;
        weights1[32427] <= 16'b0000000000000010;
        weights1[32428] <= 16'b0000000000011000;
        weights1[32429] <= 16'b0000000000101000;
        weights1[32430] <= 16'b0000000000101011;
        weights1[32431] <= 16'b0000000000100010;
        weights1[32432] <= 16'b0000000000100100;
        weights1[32433] <= 16'b0000000000101101;
        weights1[32434] <= 16'b0000000000010011;
        weights1[32435] <= 16'b1111111111100010;
        weights1[32436] <= 16'b1111111111110010;
        weights1[32437] <= 16'b1111111111001101;
        weights1[32438] <= 16'b1111111111011011;
        weights1[32439] <= 16'b1111111111001001;
        weights1[32440] <= 16'b1111111111011110;
        weights1[32441] <= 16'b1111111111011100;
        weights1[32442] <= 16'b1111111111101000;
        weights1[32443] <= 16'b1111111111110110;
        weights1[32444] <= 16'b0000000000001000;
        weights1[32445] <= 16'b1111111111111101;
        weights1[32446] <= 16'b0000000000100101;
        weights1[32447] <= 16'b0000000000001110;
        weights1[32448] <= 16'b0000000000010010;
        weights1[32449] <= 16'b1111111111101010;
        weights1[32450] <= 16'b1111111111100000;
        weights1[32451] <= 16'b1111111111100001;
        weights1[32452] <= 16'b1111111111110111;
        weights1[32453] <= 16'b1111111111100000;
        weights1[32454] <= 16'b1111111111010011;
        weights1[32455] <= 16'b1111111111110101;
        weights1[32456] <= 16'b0000000000000100;
        weights1[32457] <= 16'b0000000000010010;
        weights1[32458] <= 16'b0000000000100010;
        weights1[32459] <= 16'b0000000000110000;
        weights1[32460] <= 16'b0000000000010111;
        weights1[32461] <= 16'b0000000000100100;
        weights1[32462] <= 16'b0000000000101111;
        weights1[32463] <= 16'b0000000000010100;
        weights1[32464] <= 16'b0000000000011100;
        weights1[32465] <= 16'b0000000000000101;
        weights1[32466] <= 16'b0000000000101000;
        weights1[32467] <= 16'b1111111111110100;
        weights1[32468] <= 16'b0000000000001101;
        weights1[32469] <= 16'b0000000000011111;
        weights1[32470] <= 16'b0000000000010101;
        weights1[32471] <= 16'b0000000000010000;
        weights1[32472] <= 16'b1111111111110100;
        weights1[32473] <= 16'b0000000000001101;
        weights1[32474] <= 16'b1111111111011111;
        weights1[32475] <= 16'b1111111111011101;
        weights1[32476] <= 16'b1111111111010101;
        weights1[32477] <= 16'b1111111110111101;
        weights1[32478] <= 16'b1111111111000111;
        weights1[32479] <= 16'b1111111111011100;
        weights1[32480] <= 16'b1111111111101101;
        weights1[32481] <= 16'b1111111111011111;
        weights1[32482] <= 16'b1111111111001100;
        weights1[32483] <= 16'b1111111111010000;
        weights1[32484] <= 16'b1111111111111011;
        weights1[32485] <= 16'b0000000000011010;
        weights1[32486] <= 16'b0000000000010111;
        weights1[32487] <= 16'b0000000000110001;
        weights1[32488] <= 16'b0000000000110011;
        weights1[32489] <= 16'b0000000000110010;
        weights1[32490] <= 16'b0000000000001001;
        weights1[32491] <= 16'b0000000000100011;
        weights1[32492] <= 16'b0000000000011111;
        weights1[32493] <= 16'b0000000000010101;
        weights1[32494] <= 16'b0000000000110100;
        weights1[32495] <= 16'b0000000000010010;
        weights1[32496] <= 16'b0000000000001011;
        weights1[32497] <= 16'b0000000000011011;
        weights1[32498] <= 16'b0000000000010101;
        weights1[32499] <= 16'b0000000000100001;
        weights1[32500] <= 16'b0000000000101110;
        weights1[32501] <= 16'b0000000000001000;
        weights1[32502] <= 16'b1111111111110000;
        weights1[32503] <= 16'b1111111111010000;
        weights1[32504] <= 16'b1111111110101011;
        weights1[32505] <= 16'b1111111110110010;
        weights1[32506] <= 16'b1111111111000011;
        weights1[32507] <= 16'b1111111111010011;
        weights1[32508] <= 16'b1111111111101001;
        weights1[32509] <= 16'b1111111111011011;
        weights1[32510] <= 16'b1111111111000010;
        weights1[32511] <= 16'b1111111110111101;
        weights1[32512] <= 16'b1111111111011101;
        weights1[32513] <= 16'b1111111111100111;
        weights1[32514] <= 16'b0000000000010100;
        weights1[32515] <= 16'b0000000000110100;
        weights1[32516] <= 16'b0000000000110010;
        weights1[32517] <= 16'b0000000000011110;
        weights1[32518] <= 16'b0000000000100101;
        weights1[32519] <= 16'b0000000001001100;
        weights1[32520] <= 16'b0000000000101000;
        weights1[32521] <= 16'b0000000000100011;
        weights1[32522] <= 16'b0000000000001001;
        weights1[32523] <= 16'b0000000000010110;
        weights1[32524] <= 16'b0000000000011110;
        weights1[32525] <= 16'b0000000000010100;
        weights1[32526] <= 16'b0000000000011100;
        weights1[32527] <= 16'b0000000000001100;
        weights1[32528] <= 16'b0000000000011000;
        weights1[32529] <= 16'b0000000000000111;
        weights1[32530] <= 16'b1111111111010111;
        weights1[32531] <= 16'b1111111111010101;
        weights1[32532] <= 16'b1111111111000011;
        weights1[32533] <= 16'b1111111111001110;
        weights1[32534] <= 16'b1111111111010100;
        weights1[32535] <= 16'b1111111111011000;
        weights1[32536] <= 16'b1111111111100101;
        weights1[32537] <= 16'b1111111111010110;
        weights1[32538] <= 16'b1111111110111001;
        weights1[32539] <= 16'b1111111110100100;
        weights1[32540] <= 16'b1111111110100011;
        weights1[32541] <= 16'b1111111110111001;
        weights1[32542] <= 16'b1111111111110001;
        weights1[32543] <= 16'b1111111111111110;
        weights1[32544] <= 16'b0000000000101110;
        weights1[32545] <= 16'b0000000000100101;
        weights1[32546] <= 16'b0000000001001101;
        weights1[32547] <= 16'b0000000000010100;
        weights1[32548] <= 16'b0000000000100100;
        weights1[32549] <= 16'b0000000000101101;
        weights1[32550] <= 16'b0000000000011100;
        weights1[32551] <= 16'b0000000000100001;
        weights1[32552] <= 16'b0000000000011101;
        weights1[32553] <= 16'b0000000000010110;
        weights1[32554] <= 16'b0000000000010011;
        weights1[32555] <= 16'b1111111111011111;
        weights1[32556] <= 16'b1111111111100101;
        weights1[32557] <= 16'b1111111111100111;
        weights1[32558] <= 16'b1111111111001101;
        weights1[32559] <= 16'b1111111111100100;
        weights1[32560] <= 16'b1111111111101000;
        weights1[32561] <= 16'b1111111111101000;
        weights1[32562] <= 16'b1111111111011110;
        weights1[32563] <= 16'b1111111111011111;
        weights1[32564] <= 16'b1111111111101111;
        weights1[32565] <= 16'b1111111111100001;
        weights1[32566] <= 16'b1111111110111101;
        weights1[32567] <= 16'b1111111110110110;
        weights1[32568] <= 16'b1111111110001001;
        weights1[32569] <= 16'b1111111101100111;
        weights1[32570] <= 16'b1111111110000101;
        weights1[32571] <= 16'b1111111110101001;
        weights1[32572] <= 16'b1111111111010010;
        weights1[32573] <= 16'b1111111111111100;
        weights1[32574] <= 16'b0000000000101111;
        weights1[32575] <= 16'b0000000000100111;
        weights1[32576] <= 16'b0000000000010101;
        weights1[32577] <= 16'b0000000001000100;
        weights1[32578] <= 16'b0000000000100110;
        weights1[32579] <= 16'b0000000000100100;
        weights1[32580] <= 16'b0000000000010010;
        weights1[32581] <= 16'b0000000000001100;
        weights1[32582] <= 16'b1111111111101011;
        weights1[32583] <= 16'b1111111111110100;
        weights1[32584] <= 16'b1111111111101010;
        weights1[32585] <= 16'b1111111111011011;
        weights1[32586] <= 16'b1111111111110110;
        weights1[32587] <= 16'b1111111111111001;
        weights1[32588] <= 16'b1111111111111000;
        weights1[32589] <= 16'b1111111111101110;
        weights1[32590] <= 16'b1111111111011101;
        weights1[32591] <= 16'b1111111111100011;
        weights1[32592] <= 16'b1111111111110011;
        weights1[32593] <= 16'b1111111111101100;
        weights1[32594] <= 16'b1111111111010110;
        weights1[32595] <= 16'b1111111111000010;
        weights1[32596] <= 16'b1111111110001101;
        weights1[32597] <= 16'b1111111110001000;
        weights1[32598] <= 16'b1111111101010011;
        weights1[32599] <= 16'b1111111101010101;
        weights1[32600] <= 16'b1111111101111001;
        weights1[32601] <= 16'b1111111110010111;
        weights1[32602] <= 16'b1111111110111100;
        weights1[32603] <= 16'b1111111111110001;
        weights1[32604] <= 16'b0000000000010111;
        weights1[32605] <= 16'b0000000000010011;
        weights1[32606] <= 16'b0000000000001110;
        weights1[32607] <= 16'b0000000000010010;
        weights1[32608] <= 16'b0000000000001000;
        weights1[32609] <= 16'b1111111111101010;
        weights1[32610] <= 16'b1111111111101010;
        weights1[32611] <= 16'b1111111111101101;
        weights1[32612] <= 16'b1111111111010101;
        weights1[32613] <= 16'b1111111111110111;
        weights1[32614] <= 16'b1111111111111001;
        weights1[32615] <= 16'b0000000000010000;
        weights1[32616] <= 16'b0000000000010000;
        weights1[32617] <= 16'b1111111111111011;
        weights1[32618] <= 16'b1111111111101010;
        weights1[32619] <= 16'b1111111111100110;
        weights1[32620] <= 16'b1111111111111100;
        weights1[32621] <= 16'b1111111111111011;
        weights1[32622] <= 16'b1111111111110111;
        weights1[32623] <= 16'b1111111111110010;
        weights1[32624] <= 16'b1111111111100100;
        weights1[32625] <= 16'b1111111111010111;
        weights1[32626] <= 16'b1111111110100111;
        weights1[32627] <= 16'b1111111110001111;
        weights1[32628] <= 16'b1111111101111010;
        weights1[32629] <= 16'b1111111101101010;
        weights1[32630] <= 16'b1111111110000010;
        weights1[32631] <= 16'b1111111110011001;
        weights1[32632] <= 16'b1111111110100010;
        weights1[32633] <= 16'b1111111110100011;
        weights1[32634] <= 16'b1111111110111010;
        weights1[32635] <= 16'b1111111111001111;
        weights1[32636] <= 16'b1111111111110000;
        weights1[32637] <= 16'b1111111111101010;
        weights1[32638] <= 16'b1111111111110010;
        weights1[32639] <= 16'b1111111111011111;
        weights1[32640] <= 16'b0000000000000101;
        weights1[32641] <= 16'b0000000000011100;
        weights1[32642] <= 16'b1111111111111101;
        weights1[32643] <= 16'b0000000000100111;
        weights1[32644] <= 16'b0000000000000100;
        weights1[32645] <= 16'b1111111111111011;
        weights1[32646] <= 16'b0000000000000000;
        weights1[32647] <= 16'b1111111111100110;
        weights1[32648] <= 16'b1111111111111100;
        weights1[32649] <= 16'b1111111111111100;
        weights1[32650] <= 16'b0000000000000010;
        weights1[32651] <= 16'b0000000000001101;
        weights1[32652] <= 16'b0000000000001001;
        weights1[32653] <= 16'b0000000000010111;
        weights1[32654] <= 16'b0000000000011001;
        weights1[32655] <= 16'b1111111111101110;
        weights1[32656] <= 16'b1111111111001100;
        weights1[32657] <= 16'b1111111110110100;
        weights1[32658] <= 16'b1111111110111110;
        weights1[32659] <= 16'b1111111110111101;
        weights1[32660] <= 16'b1111111110100101;
        weights1[32661] <= 16'b1111111110111001;
        weights1[32662] <= 16'b1111111110101110;
        weights1[32663] <= 16'b1111111111011000;
        weights1[32664] <= 16'b1111111111100000;
        weights1[32665] <= 16'b1111111111100001;
        weights1[32666] <= 16'b1111111111100101;
        weights1[32667] <= 16'b1111111111111111;
        weights1[32668] <= 16'b0000000000001001;
        weights1[32669] <= 16'b0000000000000010;
        weights1[32670] <= 16'b0000000000001001;
        weights1[32671] <= 16'b0000000000010110;
        weights1[32672] <= 16'b0000000000000110;
        weights1[32673] <= 16'b0000000000000111;
        weights1[32674] <= 16'b1111111111110010;
        weights1[32675] <= 16'b1111111111101011;
        weights1[32676] <= 16'b0000000000000011;
        weights1[32677] <= 16'b0000000000001110;
        weights1[32678] <= 16'b0000000000001001;
        weights1[32679] <= 16'b0000000000001111;
        weights1[32680] <= 16'b0000000000100000;
        weights1[32681] <= 16'b0000000001000000;
        weights1[32682] <= 16'b0000000000111010;
        weights1[32683] <= 16'b0000000000101101;
        weights1[32684] <= 16'b0000000000100011;
        weights1[32685] <= 16'b0000000000001101;
        weights1[32686] <= 16'b0000000000000101;
        weights1[32687] <= 16'b1111111111100101;
        weights1[32688] <= 16'b1111111111110111;
        weights1[32689] <= 16'b1111111111110110;
        weights1[32690] <= 16'b1111111111101100;
        weights1[32691] <= 16'b1111111111100010;
        weights1[32692] <= 16'b1111111111101011;
        weights1[32693] <= 16'b0000000000001001;
        weights1[32694] <= 16'b1111111111110010;
        weights1[32695] <= 16'b1111111111101011;
        weights1[32696] <= 16'b1111111111101100;
        weights1[32697] <= 16'b1111111111101111;
        weights1[32698] <= 16'b1111111111110100;
        weights1[32699] <= 16'b1111111111110100;
        weights1[32700] <= 16'b0000000000001100;
        weights1[32701] <= 16'b0000000000010001;
        weights1[32702] <= 16'b1111111111111011;
        weights1[32703] <= 16'b1111111111110011;
        weights1[32704] <= 16'b0000000000000101;
        weights1[32705] <= 16'b0000000000001000;
        weights1[32706] <= 16'b0000000000001101;
        weights1[32707] <= 16'b0000000000010001;
        weights1[32708] <= 16'b0000000000001011;
        weights1[32709] <= 16'b0000000000001101;
        weights1[32710] <= 16'b0000000000010011;
        weights1[32711] <= 16'b0000000000010100;
        weights1[32712] <= 16'b0000000000011010;
        weights1[32713] <= 16'b0000000000000101;
        weights1[32714] <= 16'b0000000000001001;
        weights1[32715] <= 16'b0000000000010101;
        weights1[32716] <= 16'b1111111111111001;
        weights1[32717] <= 16'b1111111111111111;
        weights1[32718] <= 16'b0000000000001010;
        weights1[32719] <= 16'b0000000000000001;
        weights1[32720] <= 16'b1111111111110010;
        weights1[32721] <= 16'b0000000000000111;
        weights1[32722] <= 16'b1111111111101011;
        weights1[32723] <= 16'b1111111111110011;
        weights1[32724] <= 16'b1111111111110000;
        weights1[32725] <= 16'b0000000000001101;
        weights1[32726] <= 16'b1111111111110100;
        weights1[32727] <= 16'b1111111111111111;
        weights1[32728] <= 16'b0000000000000101;
        weights1[32729] <= 16'b0000000000001110;
        weights1[32730] <= 16'b1111111111111101;
        weights1[32731] <= 16'b1111111111101101;
        weights1[32732] <= 16'b1111111111111110;
        weights1[32733] <= 16'b0000000000000111;
        weights1[32734] <= 16'b1111111111111110;
        weights1[32735] <= 16'b1111111111111010;
        weights1[32736] <= 16'b1111111111110110;
        weights1[32737] <= 16'b0000000000100011;
        weights1[32738] <= 16'b0000000000010101;
        weights1[32739] <= 16'b1111111111110011;
        weights1[32740] <= 16'b0000000000000000;
        weights1[32741] <= 16'b0000000000011000;
        weights1[32742] <= 16'b0000000000001101;
        weights1[32743] <= 16'b1111111111110010;
        weights1[32744] <= 16'b0000000000010001;
        weights1[32745] <= 16'b1111111111101010;
        weights1[32746] <= 16'b1111111111110001;
        weights1[32747] <= 16'b1111111111101001;
        weights1[32748] <= 16'b1111111111101011;
        weights1[32749] <= 16'b1111111111111110;
        weights1[32750] <= 16'b1111111111110101;
        weights1[32751] <= 16'b1111111111111011;
        weights1[32752] <= 16'b0000000000010000;
        weights1[32753] <= 16'b0000000000010000;
        weights1[32754] <= 16'b0000000000001010;
        weights1[32755] <= 16'b1111111111011011;
        weights1[32756] <= 16'b0000000000001011;
        weights1[32757] <= 16'b0000000000010000;
        weights1[32758] <= 16'b1111111111111011;
        weights1[32759] <= 16'b1111111111111001;
        weights1[32760] <= 16'b1111111111110100;
        weights1[32761] <= 16'b1111111111111000;
        weights1[32762] <= 16'b1111111111101011;
        weights1[32763] <= 16'b1111111111110111;
        weights1[32764] <= 16'b0000000000001001;
        weights1[32765] <= 16'b0000000000010000;
        weights1[32766] <= 16'b1111111111101100;
        weights1[32767] <= 16'b0000000000001110;
        weights1[32768] <= 16'b1111111111110001;
        weights1[32769] <= 16'b0000000000001111;
        weights1[32770] <= 16'b1111111111101100;
        weights1[32771] <= 16'b1111111111101011;
        weights1[32772] <= 16'b1111111111111101;
        weights1[32773] <= 16'b0000000000000010;
        weights1[32774] <= 16'b0000000000001010;
        weights1[32775] <= 16'b0000000000000110;
        weights1[32776] <= 16'b0000000000001101;
        weights1[32777] <= 16'b0000000000000101;
        weights1[32778] <= 16'b1111111111101001;
        weights1[32779] <= 16'b1111111111110001;
        weights1[32780] <= 16'b1111111111110100;
        weights1[32781] <= 16'b0000000000011010;
        weights1[32782] <= 16'b1111111111101110;
        weights1[32783] <= 16'b1111111111111111;
        weights1[32784] <= 16'b1111111111111000;
        weights1[32785] <= 16'b1111111111111001;
        weights1[32786] <= 16'b1111111111110001;
        weights1[32787] <= 16'b1111111111111011;
        weights1[32788] <= 16'b1111111111111000;
        weights1[32789] <= 16'b1111111111110011;
        weights1[32790] <= 16'b1111111111101101;
        weights1[32791] <= 16'b1111111111110100;
        weights1[32792] <= 16'b1111111111101110;
        weights1[32793] <= 16'b1111111111101111;
        weights1[32794] <= 16'b0000000000001000;
        weights1[32795] <= 16'b1111111111110000;
        weights1[32796] <= 16'b0000000000010000;
        weights1[32797] <= 16'b0000000000000100;
        weights1[32798] <= 16'b1111111111111101;
        weights1[32799] <= 16'b0000000000100111;
        weights1[32800] <= 16'b0000000000001110;
        weights1[32801] <= 16'b0000000000000000;
        weights1[32802] <= 16'b0000000000010010;
        weights1[32803] <= 16'b1111111111110001;
        weights1[32804] <= 16'b1111111111111000;
        weights1[32805] <= 16'b1111111111110111;
        weights1[32806] <= 16'b1111111111110011;
        weights1[32807] <= 16'b1111111111111101;
        weights1[32808] <= 16'b1111111111101110;
        weights1[32809] <= 16'b0000000000010011;
        weights1[32810] <= 16'b1111111111101100;
        weights1[32811] <= 16'b1111111111111100;
        weights1[32812] <= 16'b1111111111101110;
        weights1[32813] <= 16'b1111111111111001;
        weights1[32814] <= 16'b1111111111111101;
        weights1[32815] <= 16'b1111111111111110;
        weights1[32816] <= 16'b1111111111110111;
        weights1[32817] <= 16'b1111111111111011;
        weights1[32818] <= 16'b1111111111110001;
        weights1[32819] <= 16'b1111111111101110;
        weights1[32820] <= 16'b1111111111111001;
        weights1[32821] <= 16'b1111111111110000;
        weights1[32822] <= 16'b1111111111110011;
        weights1[32823] <= 16'b0000000000000111;
        weights1[32824] <= 16'b0000000000000110;
        weights1[32825] <= 16'b1111111111100011;
        weights1[32826] <= 16'b0000000000000110;
        weights1[32827] <= 16'b0000000000010100;
        weights1[32828] <= 16'b1111111111101010;
        weights1[32829] <= 16'b0000000000001101;
        weights1[32830] <= 16'b0000000000000010;
        weights1[32831] <= 16'b1111111111110100;
        weights1[32832] <= 16'b1111111111101010;
        weights1[32833] <= 16'b1111111111101010;
        weights1[32834] <= 16'b1111111111100101;
        weights1[32835] <= 16'b1111111111111100;
        weights1[32836] <= 16'b0000000000001010;
        weights1[32837] <= 16'b0000000000000110;
        weights1[32838] <= 16'b1111111111101110;
        weights1[32839] <= 16'b1111111111110010;
        weights1[32840] <= 16'b1111111111110011;
        weights1[32841] <= 16'b1111111111110000;
        weights1[32842] <= 16'b0000000000000001;
        weights1[32843] <= 16'b1111111111111110;
        weights1[32844] <= 16'b1111111111111011;
        weights1[32845] <= 16'b1111111111110111;
        weights1[32846] <= 16'b1111111111110110;
        weights1[32847] <= 16'b1111111111110100;
        weights1[32848] <= 16'b1111111111100111;
        weights1[32849] <= 16'b1111111111100111;
        weights1[32850] <= 16'b1111111111011010;
        weights1[32851] <= 16'b1111111111110101;
        weights1[32852] <= 16'b1111111111110001;
        weights1[32853] <= 16'b1111111111101011;
        weights1[32854] <= 16'b1111111111110111;
        weights1[32855] <= 16'b0000000000000010;
        weights1[32856] <= 16'b1111111111100110;
        weights1[32857] <= 16'b0000000000010000;
        weights1[32858] <= 16'b1111111111100110;
        weights1[32859] <= 16'b1111111111110000;
        weights1[32860] <= 16'b0000000000000001;
        weights1[32861] <= 16'b0000000000000100;
        weights1[32862] <= 16'b1111111111110110;
        weights1[32863] <= 16'b0000000000010000;
        weights1[32864] <= 16'b0000000000010000;
        weights1[32865] <= 16'b0000000000000000;
        weights1[32866] <= 16'b0000000000000110;
        weights1[32867] <= 16'b1111111111111101;
        weights1[32868] <= 16'b1111111111111001;
        weights1[32869] <= 16'b1111111111111000;
        weights1[32870] <= 16'b1111111111111011;
        weights1[32871] <= 16'b1111111111111110;
        weights1[32872] <= 16'b1111111111111110;
        weights1[32873] <= 16'b1111111111110111;
        weights1[32874] <= 16'b1111111111110101;
        weights1[32875] <= 16'b1111111111111010;
        weights1[32876] <= 16'b1111111111110111;
        weights1[32877] <= 16'b1111111111111010;
        weights1[32878] <= 16'b1111111111101001;
        weights1[32879] <= 16'b1111111111101001;
        weights1[32880] <= 16'b1111111111101001;
        weights1[32881] <= 16'b1111111111100010;
        weights1[32882] <= 16'b1111111111110110;
        weights1[32883] <= 16'b1111111111101110;
        weights1[32884] <= 16'b1111111111110010;
        weights1[32885] <= 16'b1111111111111101;
        weights1[32886] <= 16'b0000000000001001;
        weights1[32887] <= 16'b1111111111101110;
        weights1[32888] <= 16'b0000000000010110;
        weights1[32889] <= 16'b0000000000001001;
        weights1[32890] <= 16'b1111111111101110;
        weights1[32891] <= 16'b1111111111110111;
        weights1[32892] <= 16'b1111111111111010;
        weights1[32893] <= 16'b1111111111111010;
        weights1[32894] <= 16'b0000000000000111;
        weights1[32895] <= 16'b0000000000000010;
        weights1[32896] <= 16'b1111111111111011;
        weights1[32897] <= 16'b1111111111111011;
        weights1[32898] <= 16'b1111111111111101;
        weights1[32899] <= 16'b0000000000000000;
        weights1[32900] <= 16'b0000000000000000;
        weights1[32901] <= 16'b1111111111111100;
        weights1[32902] <= 16'b1111111111111100;
        weights1[32903] <= 16'b1111111111110110;
        weights1[32904] <= 16'b1111111111110110;
        weights1[32905] <= 16'b1111111111110101;
        weights1[32906] <= 16'b1111111111110110;
        weights1[32907] <= 16'b1111111111101011;
        weights1[32908] <= 16'b1111111111011110;
        weights1[32909] <= 16'b1111111111011111;
        weights1[32910] <= 16'b1111111111100100;
        weights1[32911] <= 16'b1111111111100000;
        weights1[32912] <= 16'b1111111111011110;
        weights1[32913] <= 16'b1111111111110000;
        weights1[32914] <= 16'b1111111111111110;
        weights1[32915] <= 16'b1111111111110001;
        weights1[32916] <= 16'b1111111111110000;
        weights1[32917] <= 16'b1111111111110100;
        weights1[32918] <= 16'b1111111111111011;
        weights1[32919] <= 16'b1111111111111100;
        weights1[32920] <= 16'b1111111111111101;
        weights1[32921] <= 16'b1111111111111001;
        weights1[32922] <= 16'b1111111111111010;
        weights1[32923] <= 16'b1111111111111010;
        weights1[32924] <= 16'b1111111111111011;
        weights1[32925] <= 16'b1111111111111101;
        weights1[32926] <= 16'b1111111111111110;
        weights1[32927] <= 16'b0000000000000000;
        weights1[32928] <= 16'b0000000000000000;
        weights1[32929] <= 16'b0000000000000000;
        weights1[32930] <= 16'b1111111111111111;
        weights1[32931] <= 16'b1111111111111111;
        weights1[32932] <= 16'b1111111111111111;
        weights1[32933] <= 16'b1111111111111110;
        weights1[32934] <= 16'b1111111111111110;
        weights1[32935] <= 16'b1111111111111010;
        weights1[32936] <= 16'b1111111111110110;
        weights1[32937] <= 16'b1111111111101110;
        weights1[32938] <= 16'b1111111111110000;
        weights1[32939] <= 16'b1111111111110111;
        weights1[32940] <= 16'b1111111111110110;
        weights1[32941] <= 16'b1111111111110000;
        weights1[32942] <= 16'b1111111111101111;
        weights1[32943] <= 16'b1111111111101111;
        weights1[32944] <= 16'b1111111111111011;
        weights1[32945] <= 16'b1111111111111000;
        weights1[32946] <= 16'b1111111111110110;
        weights1[32947] <= 16'b1111111111110110;
        weights1[32948] <= 16'b1111111111111000;
        weights1[32949] <= 16'b1111111111110111;
        weights1[32950] <= 16'b1111111111111101;
        weights1[32951] <= 16'b1111111111111110;
        weights1[32952] <= 16'b1111111111111110;
        weights1[32953] <= 16'b1111111111111111;
        weights1[32954] <= 16'b0000000000000000;
        weights1[32955] <= 16'b0000000000000000;
        weights1[32956] <= 16'b0000000000000000;
        weights1[32957] <= 16'b0000000000000000;
        weights1[32958] <= 16'b0000000000000000;
        weights1[32959] <= 16'b1111111111111111;
        weights1[32960] <= 16'b0000000000000000;
        weights1[32961] <= 16'b1111111111111111;
        weights1[32962] <= 16'b1111111111111001;
        weights1[32963] <= 16'b1111111111110100;
        weights1[32964] <= 16'b1111111111101100;
        weights1[32965] <= 16'b1111111111100011;
        weights1[32966] <= 16'b1111111111011111;
        weights1[32967] <= 16'b1111111111110001;
        weights1[32968] <= 16'b1111111111110010;
        weights1[32969] <= 16'b1111111111100111;
        weights1[32970] <= 16'b1111111111011100;
        weights1[32971] <= 16'b1111111111100011;
        weights1[32972] <= 16'b1111111111101010;
        weights1[32973] <= 16'b1111111111101110;
        weights1[32974] <= 16'b1111111111101100;
        weights1[32975] <= 16'b1111111111110010;
        weights1[32976] <= 16'b1111111111110101;
        weights1[32977] <= 16'b1111111111110111;
        weights1[32978] <= 16'b1111111111111100;
        weights1[32979] <= 16'b1111111111111100;
        weights1[32980] <= 16'b1111111111111011;
        weights1[32981] <= 16'b1111111111111111;
        weights1[32982] <= 16'b1111111111111110;
        weights1[32983] <= 16'b1111111111111110;
        weights1[32984] <= 16'b0000000000000000;
        weights1[32985] <= 16'b0000000000000000;
        weights1[32986] <= 16'b0000000000000000;
        weights1[32987] <= 16'b1111111111111111;
        weights1[32988] <= 16'b1111111111111111;
        weights1[32989] <= 16'b1111111111111011;
        weights1[32990] <= 16'b1111111111110100;
        weights1[32991] <= 16'b1111111111101111;
        weights1[32992] <= 16'b1111111111101000;
        weights1[32993] <= 16'b1111111111100010;
        weights1[32994] <= 16'b1111111111011011;
        weights1[32995] <= 16'b1111111111010100;
        weights1[32996] <= 16'b1111111111101100;
        weights1[32997] <= 16'b1111111111011111;
        weights1[32998] <= 16'b1111111111001110;
        weights1[32999] <= 16'b1111111111010111;
        weights1[33000] <= 16'b1111111111100001;
        weights1[33001] <= 16'b1111111111101111;
        weights1[33002] <= 16'b1111111111101101;
        weights1[33003] <= 16'b1111111111101010;
        weights1[33004] <= 16'b1111111111101011;
        weights1[33005] <= 16'b1111111111101000;
        weights1[33006] <= 16'b1111111111101100;
        weights1[33007] <= 16'b1111111111110101;
        weights1[33008] <= 16'b1111111111111010;
        weights1[33009] <= 16'b1111111111111110;
        weights1[33010] <= 16'b0000000000000010;
        weights1[33011] <= 16'b1111111111111101;
        weights1[33012] <= 16'b0000000000000000;
        weights1[33013] <= 16'b1111111111111111;
        weights1[33014] <= 16'b1111111111111101;
        weights1[33015] <= 16'b1111111111111111;
        weights1[33016] <= 16'b1111111111111011;
        weights1[33017] <= 16'b1111111111111100;
        weights1[33018] <= 16'b1111111111101110;
        weights1[33019] <= 16'b1111111111100111;
        weights1[33020] <= 16'b1111111111101011;
        weights1[33021] <= 16'b1111111111001111;
        weights1[33022] <= 16'b1111111111001011;
        weights1[33023] <= 16'b1111111111001111;
        weights1[33024] <= 16'b1111111111101101;
        weights1[33025] <= 16'b1111111111001100;
        weights1[33026] <= 16'b1111111111001001;
        weights1[33027] <= 16'b1111111110110011;
        weights1[33028] <= 16'b1111111111010101;
        weights1[33029] <= 16'b1111111111001011;
        weights1[33030] <= 16'b1111111111001001;
        weights1[33031] <= 16'b1111111111010001;
        weights1[33032] <= 16'b1111111111011111;
        weights1[33033] <= 16'b1111111111100000;
        weights1[33034] <= 16'b1111111111101001;
        weights1[33035] <= 16'b1111111111101111;
        weights1[33036] <= 16'b1111111111110110;
        weights1[33037] <= 16'b0000000000000000;
        weights1[33038] <= 16'b0000000000000011;
        weights1[33039] <= 16'b1111111111111110;
        weights1[33040] <= 16'b1111111111111111;
        weights1[33041] <= 16'b1111111111111011;
        weights1[33042] <= 16'b1111111111111100;
        weights1[33043] <= 16'b1111111111111011;
        weights1[33044] <= 16'b1111111111111110;
        weights1[33045] <= 16'b1111111111110101;
        weights1[33046] <= 16'b1111111111101110;
        weights1[33047] <= 16'b1111111111010010;
        weights1[33048] <= 16'b1111111111010110;
        weights1[33049] <= 16'b1111111110110111;
        weights1[33050] <= 16'b1111111110111110;
        weights1[33051] <= 16'b1111111111000001;
        weights1[33052] <= 16'b1111111111010001;
        weights1[33053] <= 16'b1111111111010111;
        weights1[33054] <= 16'b1111111111010100;
        weights1[33055] <= 16'b1111111111001101;
        weights1[33056] <= 16'b1111111111111101;
        weights1[33057] <= 16'b1111111111101101;
        weights1[33058] <= 16'b1111111111011110;
        weights1[33059] <= 16'b1111111111011000;
        weights1[33060] <= 16'b1111111111011000;
        weights1[33061] <= 16'b1111111111101100;
        weights1[33062] <= 16'b1111111111111001;
        weights1[33063] <= 16'b1111111111111100;
        weights1[33064] <= 16'b0000000000000001;
        weights1[33065] <= 16'b0000000000000101;
        weights1[33066] <= 16'b0000000000000011;
        weights1[33067] <= 16'b1111111111111101;
        weights1[33068] <= 16'b1111111111111101;
        weights1[33069] <= 16'b1111111111111010;
        weights1[33070] <= 16'b1111111111111011;
        weights1[33071] <= 16'b1111111111111001;
        weights1[33072] <= 16'b1111111111110111;
        weights1[33073] <= 16'b1111111111101111;
        weights1[33074] <= 16'b1111111111111010;
        weights1[33075] <= 16'b1111111111101010;
        weights1[33076] <= 16'b1111111111101000;
        weights1[33077] <= 16'b1111111111011001;
        weights1[33078] <= 16'b1111111111101110;
        weights1[33079] <= 16'b1111111111000101;
        weights1[33080] <= 16'b1111111111011010;
        weights1[33081] <= 16'b1111111111011011;
        weights1[33082] <= 16'b1111111111110001;
        weights1[33083] <= 16'b1111111111101001;
        weights1[33084] <= 16'b1111111111101000;
        weights1[33085] <= 16'b1111111111101011;
        weights1[33086] <= 16'b1111111111110100;
        weights1[33087] <= 16'b1111111111100110;
        weights1[33088] <= 16'b1111111111110001;
        weights1[33089] <= 16'b1111111111101100;
        weights1[33090] <= 16'b1111111111111000;
        weights1[33091] <= 16'b1111111111111100;
        weights1[33092] <= 16'b0000000000001100;
        weights1[33093] <= 16'b0000000000000110;
        weights1[33094] <= 16'b1111111111111010;
        weights1[33095] <= 16'b1111111111111011;
        weights1[33096] <= 16'b1111111111111100;
        weights1[33097] <= 16'b1111111111110111;
        weights1[33098] <= 16'b1111111111110000;
        weights1[33099] <= 16'b1111111111101110;
        weights1[33100] <= 16'b1111111111110110;
        weights1[33101] <= 16'b1111111111111101;
        weights1[33102] <= 16'b1111111111111000;
        weights1[33103] <= 16'b0000000000000010;
        weights1[33104] <= 16'b0000000000010100;
        weights1[33105] <= 16'b1111111111011110;
        weights1[33106] <= 16'b0000000000010100;
        weights1[33107] <= 16'b1111111111110001;
        weights1[33108] <= 16'b0000000000010010;
        weights1[33109] <= 16'b0000000000010001;
        weights1[33110] <= 16'b1111111111100110;
        weights1[33111] <= 16'b1111111111111001;
        weights1[33112] <= 16'b1111111111101110;
        weights1[33113] <= 16'b1111111111110000;
        weights1[33114] <= 16'b0000000000010100;
        weights1[33115] <= 16'b0000000000001000;
        weights1[33116] <= 16'b1111111111111010;
        weights1[33117] <= 16'b0000000000001010;
        weights1[33118] <= 16'b0000000000001001;
        weights1[33119] <= 16'b0000000000010011;
        weights1[33120] <= 16'b0000000000010110;
        weights1[33121] <= 16'b1111111111111100;
        weights1[33122] <= 16'b1111111111111011;
        weights1[33123] <= 16'b1111111111111101;
        weights1[33124] <= 16'b1111111111111011;
        weights1[33125] <= 16'b1111111111110111;
        weights1[33126] <= 16'b1111111111101101;
        weights1[33127] <= 16'b1111111111101100;
        weights1[33128] <= 16'b1111111111101011;
        weights1[33129] <= 16'b1111111111101000;
        weights1[33130] <= 16'b1111111111111000;
        weights1[33131] <= 16'b0000000000010000;
        weights1[33132] <= 16'b0000000000001111;
        weights1[33133] <= 16'b0000000000010000;
        weights1[33134] <= 16'b0000000000010110;
        weights1[33135] <= 16'b0000000000011101;
        weights1[33136] <= 16'b0000000000100000;
        weights1[33137] <= 16'b1111111111111000;
        weights1[33138] <= 16'b1111111111111000;
        weights1[33139] <= 16'b1111111111111000;
        weights1[33140] <= 16'b0000000000000110;
        weights1[33141] <= 16'b1111111111111000;
        weights1[33142] <= 16'b0000000000010010;
        weights1[33143] <= 16'b0000000000010100;
        weights1[33144] <= 16'b0000000000000000;
        weights1[33145] <= 16'b0000000000010001;
        weights1[33146] <= 16'b0000000000010001;
        weights1[33147] <= 16'b0000000000010101;
        weights1[33148] <= 16'b0000000000001101;
        weights1[33149] <= 16'b0000000000001001;
        weights1[33150] <= 16'b1111111111111110;
        weights1[33151] <= 16'b0000000000000001;
        weights1[33152] <= 16'b1111111111111010;
        weights1[33153] <= 16'b1111111111110010;
        weights1[33154] <= 16'b1111111111101101;
        weights1[33155] <= 16'b1111111111011110;
        weights1[33156] <= 16'b1111111111001001;
        weights1[33157] <= 16'b1111111111110011;
        weights1[33158] <= 16'b1111111111010100;
        weights1[33159] <= 16'b0000000000000010;
        weights1[33160] <= 16'b0000000000011101;
        weights1[33161] <= 16'b1111111111111101;
        weights1[33162] <= 16'b0000000000011010;
        weights1[33163] <= 16'b0000000000110001;
        weights1[33164] <= 16'b0000000000110000;
        weights1[33165] <= 16'b0000000000010000;
        weights1[33166] <= 16'b0000000000010011;
        weights1[33167] <= 16'b0000000000001101;
        weights1[33168] <= 16'b0000000000010010;
        weights1[33169] <= 16'b0000000000010010;
        weights1[33170] <= 16'b0000000000010000;
        weights1[33171] <= 16'b0000000000000010;
        weights1[33172] <= 16'b0000000000100000;
        weights1[33173] <= 16'b0000000000000011;
        weights1[33174] <= 16'b1111111111110111;
        weights1[33175] <= 16'b0000000000001110;
        weights1[33176] <= 16'b0000000000000110;
        weights1[33177] <= 16'b0000000000000110;
        weights1[33178] <= 16'b0000000000000011;
        weights1[33179] <= 16'b1111111111111010;
        weights1[33180] <= 16'b1111111111111000;
        weights1[33181] <= 16'b1111111111110110;
        weights1[33182] <= 16'b1111111111101011;
        weights1[33183] <= 16'b1111111111101011;
        weights1[33184] <= 16'b1111111111101111;
        weights1[33185] <= 16'b0000000000000000;
        weights1[33186] <= 16'b0000000000001101;
        weights1[33187] <= 16'b1111111111110100;
        weights1[33188] <= 16'b0000000000100011;
        weights1[33189] <= 16'b0000000000011111;
        weights1[33190] <= 16'b0000000000111110;
        weights1[33191] <= 16'b0000000000101010;
        weights1[33192] <= 16'b0000000000011001;
        weights1[33193] <= 16'b0000000000110001;
        weights1[33194] <= 16'b0000000000101100;
        weights1[33195] <= 16'b0000000000011010;
        weights1[33196] <= 16'b1111111111110010;
        weights1[33197] <= 16'b0000000000010110;
        weights1[33198] <= 16'b0000000000011100;
        weights1[33199] <= 16'b0000000000010100;
        weights1[33200] <= 16'b0000000000101110;
        weights1[33201] <= 16'b0000000000011001;
        weights1[33202] <= 16'b0000000000010011;
        weights1[33203] <= 16'b0000000000000000;
        weights1[33204] <= 16'b0000000000000100;
        weights1[33205] <= 16'b0000000000000000;
        weights1[33206] <= 16'b1111111111101110;
        weights1[33207] <= 16'b0000000000010001;
        weights1[33208] <= 16'b1111111111111010;
        weights1[33209] <= 16'b1111111111101111;
        weights1[33210] <= 16'b1111111111110010;
        weights1[33211] <= 16'b1111111111110001;
        weights1[33212] <= 16'b0000000000000001;
        weights1[33213] <= 16'b1111111111111011;
        weights1[33214] <= 16'b0000000000000011;
        weights1[33215] <= 16'b0000000000000110;
        weights1[33216] <= 16'b0000000000001101;
        weights1[33217] <= 16'b0000000000010111;
        weights1[33218] <= 16'b0000000000000001;
        weights1[33219] <= 16'b0000000000110100;
        weights1[33220] <= 16'b0000000000101010;
        weights1[33221] <= 16'b0000000000111100;
        weights1[33222] <= 16'b0000000000110000;
        weights1[33223] <= 16'b0000000000101110;
        weights1[33224] <= 16'b0000000000001011;
        weights1[33225] <= 16'b0000000000101110;
        weights1[33226] <= 16'b0000000000000001;
        weights1[33227] <= 16'b0000000000001101;
        weights1[33228] <= 16'b0000000000001001;
        weights1[33229] <= 16'b0000000000011011;
        weights1[33230] <= 16'b0000000000011101;
        weights1[33231] <= 16'b0000000000000001;
        weights1[33232] <= 16'b0000000000000100;
        weights1[33233] <= 16'b0000000000000001;
        weights1[33234] <= 16'b0000000000000110;
        weights1[33235] <= 16'b0000000000010001;
        weights1[33236] <= 16'b1111111111111001;
        weights1[33237] <= 16'b1111111111110111;
        weights1[33238] <= 16'b1111111111110111;
        weights1[33239] <= 16'b1111111111111000;
        weights1[33240] <= 16'b1111111111101101;
        weights1[33241] <= 16'b1111111111101111;
        weights1[33242] <= 16'b1111111111111101;
        weights1[33243] <= 16'b1111111111111000;
        weights1[33244] <= 16'b1111111111101000;
        weights1[33245] <= 16'b0000000000001100;
        weights1[33246] <= 16'b0000000000100010;
        weights1[33247] <= 16'b0000000000011100;
        weights1[33248] <= 16'b0000000000010100;
        weights1[33249] <= 16'b1111111111110001;
        weights1[33250] <= 16'b1111111111101010;
        weights1[33251] <= 16'b0000000000001110;
        weights1[33252] <= 16'b1111111111111000;
        weights1[33253] <= 16'b0000000000010001;
        weights1[33254] <= 16'b0000000000100010;
        weights1[33255] <= 16'b0000000000001111;
        weights1[33256] <= 16'b0000000000100101;
        weights1[33257] <= 16'b0000000000000010;
        weights1[33258] <= 16'b0000000000011111;
        weights1[33259] <= 16'b0000000000000111;
        weights1[33260] <= 16'b1111111111111011;
        weights1[33261] <= 16'b1111111111101000;
        weights1[33262] <= 16'b0000000000000101;
        weights1[33263] <= 16'b0000000000010111;
        weights1[33264] <= 16'b1111111111111100;
        weights1[33265] <= 16'b0000000000000010;
        weights1[33266] <= 16'b0000000000000011;
        weights1[33267] <= 16'b1111111111101111;
        weights1[33268] <= 16'b1111111111110111;
        weights1[33269] <= 16'b1111111111101001;
        weights1[33270] <= 16'b0000000000001001;
        weights1[33271] <= 16'b1111111111110100;
        weights1[33272] <= 16'b1111111111111011;
        weights1[33273] <= 16'b0000000000000101;
        weights1[33274] <= 16'b0000000000001001;
        weights1[33275] <= 16'b0000000000001111;
        weights1[33276] <= 16'b0000000000000010;
        weights1[33277] <= 16'b1111111110110111;
        weights1[33278] <= 16'b1111111110111100;
        weights1[33279] <= 16'b1111111111010110;
        weights1[33280] <= 16'b1111111111110010;
        weights1[33281] <= 16'b1111111111111111;
        weights1[33282] <= 16'b1111111111110100;
        weights1[33283] <= 16'b1111111111110000;
        weights1[33284] <= 16'b0000000000001011;
        weights1[33285] <= 16'b1111111111110101;
        weights1[33286] <= 16'b0000000000001110;
        weights1[33287] <= 16'b0000000000000101;
        weights1[33288] <= 16'b0000000000000010;
        weights1[33289] <= 16'b1111111111101010;
        weights1[33290] <= 16'b1111111111111100;
        weights1[33291] <= 16'b0000000000001111;
        weights1[33292] <= 16'b1111111111111101;
        weights1[33293] <= 16'b0000000000001000;
        weights1[33294] <= 16'b1111111111111001;
        weights1[33295] <= 16'b1111111111110010;
        weights1[33296] <= 16'b1111111111111101;
        weights1[33297] <= 16'b1111111111111100;
        weights1[33298] <= 16'b1111111111111001;
        weights1[33299] <= 16'b0000000000000011;
        weights1[33300] <= 16'b0000000000010011;
        weights1[33301] <= 16'b0000000000001000;
        weights1[33302] <= 16'b0000000000001110;
        weights1[33303] <= 16'b0000000000000100;
        weights1[33304] <= 16'b1111111111001111;
        weights1[33305] <= 16'b1111111110000001;
        weights1[33306] <= 16'b1111111110001010;
        weights1[33307] <= 16'b1111111111010011;
        weights1[33308] <= 16'b1111111111101101;
        weights1[33309] <= 16'b0000000000000100;
        weights1[33310] <= 16'b1111111111010110;
        weights1[33311] <= 16'b0000000000000111;
        weights1[33312] <= 16'b1111111111111001;
        weights1[33313] <= 16'b1111111111111100;
        weights1[33314] <= 16'b0000000000000001;
        weights1[33315] <= 16'b1111111111111010;
        weights1[33316] <= 16'b1111111111111100;
        weights1[33317] <= 16'b1111111111101111;
        weights1[33318] <= 16'b0000000000000000;
        weights1[33319] <= 16'b0000000000000111;
        weights1[33320] <= 16'b0000000000000110;
        weights1[33321] <= 16'b0000000000001011;
        weights1[33322] <= 16'b1111111111110101;
        weights1[33323] <= 16'b1111111111111011;
        weights1[33324] <= 16'b1111111111110010;
        weights1[33325] <= 16'b0000000000100110;
        weights1[33326] <= 16'b0000000000000100;
        weights1[33327] <= 16'b0000000000010101;
        weights1[33328] <= 16'b0000000000000001;
        weights1[33329] <= 16'b1111111111111100;
        weights1[33330] <= 16'b0000000000011100;
        weights1[33331] <= 16'b0000000000000110;
        weights1[33332] <= 16'b1111111110100011;
        weights1[33333] <= 16'b1111111101011011;
        weights1[33334] <= 16'b1111111111010010;
        weights1[33335] <= 16'b1111111111101111;
        weights1[33336] <= 16'b1111111111110000;
        weights1[33337] <= 16'b1111111111010110;
        weights1[33338] <= 16'b1111111111011101;
        weights1[33339] <= 16'b1111111111011111;
        weights1[33340] <= 16'b1111111111110110;
        weights1[33341] <= 16'b1111111111101101;
        weights1[33342] <= 16'b1111111111111111;
        weights1[33343] <= 16'b0000000000000111;
        weights1[33344] <= 16'b0000000000001000;
        weights1[33345] <= 16'b1111111111100001;
        weights1[33346] <= 16'b1111111111111011;
        weights1[33347] <= 16'b0000000000000000;
        weights1[33348] <= 16'b0000000000001000;
        weights1[33349] <= 16'b0000000000001100;
        weights1[33350] <= 16'b1111111111111000;
        weights1[33351] <= 16'b0000000000000011;
        weights1[33352] <= 16'b0000000000000000;
        weights1[33353] <= 16'b0000000000010010;
        weights1[33354] <= 16'b0000000000100001;
        weights1[33355] <= 16'b0000000000011101;
        weights1[33356] <= 16'b0000000000000100;
        weights1[33357] <= 16'b0000000000010000;
        weights1[33358] <= 16'b0000000000101100;
        weights1[33359] <= 16'b1111111111011100;
        weights1[33360] <= 16'b1111111101101111;
        weights1[33361] <= 16'b1111111100111110;
        weights1[33362] <= 16'b1111111111011011;
        weights1[33363] <= 16'b1111111111111011;
        weights1[33364] <= 16'b1111111111101010;
        weights1[33365] <= 16'b1111111111010101;
        weights1[33366] <= 16'b1111111111101001;
        weights1[33367] <= 16'b1111111111011101;
        weights1[33368] <= 16'b1111111111100011;
        weights1[33369] <= 16'b1111111111111110;
        weights1[33370] <= 16'b1111111111101010;
        weights1[33371] <= 16'b1111111111110011;
        weights1[33372] <= 16'b1111111111111100;
        weights1[33373] <= 16'b1111111111110000;
        weights1[33374] <= 16'b1111111111110000;
        weights1[33375] <= 16'b1111111111111111;
        weights1[33376] <= 16'b0000000000001100;
        weights1[33377] <= 16'b0000000000001100;
        weights1[33378] <= 16'b0000000000000111;
        weights1[33379] <= 16'b0000000000010001;
        weights1[33380] <= 16'b1111111111110101;
        weights1[33381] <= 16'b0000000000001110;
        weights1[33382] <= 16'b0000000000010010;
        weights1[33383] <= 16'b1111111111111100;
        weights1[33384] <= 16'b0000000000100000;
        weights1[33385] <= 16'b0000000000000111;
        weights1[33386] <= 16'b0000000000010100;
        weights1[33387] <= 16'b1111111110101000;
        weights1[33388] <= 16'b1111111101001100;
        weights1[33389] <= 16'b1111111110011101;
        weights1[33390] <= 16'b1111111111101010;
        weights1[33391] <= 16'b1111111111101101;
        weights1[33392] <= 16'b1111111111010101;
        weights1[33393] <= 16'b1111111111011111;
        weights1[33394] <= 16'b1111111111101100;
        weights1[33395] <= 16'b1111111111111101;
        weights1[33396] <= 16'b1111111111101111;
        weights1[33397] <= 16'b0000000000001001;
        weights1[33398] <= 16'b1111111111101101;
        weights1[33399] <= 16'b1111111111101011;
        weights1[33400] <= 16'b0000000000000001;
        weights1[33401] <= 16'b1111111111101101;
        weights1[33402] <= 16'b1111111111110111;
        weights1[33403] <= 16'b1111111111111101;
        weights1[33404] <= 16'b0000000000001010;
        weights1[33405] <= 16'b0000000000001100;
        weights1[33406] <= 16'b0000000000001110;
        weights1[33407] <= 16'b1111111111111101;
        weights1[33408] <= 16'b0000000000001000;
        weights1[33409] <= 16'b0000000000000111;
        weights1[33410] <= 16'b0000000000001010;
        weights1[33411] <= 16'b0000000000001100;
        weights1[33412] <= 16'b0000000000000000;
        weights1[33413] <= 16'b1111111111111111;
        weights1[33414] <= 16'b1111111111001010;
        weights1[33415] <= 16'b1111111101110000;
        weights1[33416] <= 16'b1111111101000101;
        weights1[33417] <= 16'b1111111111101111;
        weights1[33418] <= 16'b0000000000000011;
        weights1[33419] <= 16'b1111111111011100;
        weights1[33420] <= 16'b1111111111011101;
        weights1[33421] <= 16'b0000000000000010;
        weights1[33422] <= 16'b1111111111110110;
        weights1[33423] <= 16'b1111111111101100;
        weights1[33424] <= 16'b0000000000000000;
        weights1[33425] <= 16'b1111111111110000;
        weights1[33426] <= 16'b0000000000000011;
        weights1[33427] <= 16'b1111111111111011;
        weights1[33428] <= 16'b1111111111111000;
        weights1[33429] <= 16'b1111111111101010;
        weights1[33430] <= 16'b1111111111110110;
        weights1[33431] <= 16'b1111111111111011;
        weights1[33432] <= 16'b0000000000001110;
        weights1[33433] <= 16'b0000000000011100;
        weights1[33434] <= 16'b0000000000010100;
        weights1[33435] <= 16'b0000000000001110;
        weights1[33436] <= 16'b0000000000000111;
        weights1[33437] <= 16'b0000000000001110;
        weights1[33438] <= 16'b0000000000000111;
        weights1[33439] <= 16'b0000000000000010;
        weights1[33440] <= 16'b1111111111110011;
        weights1[33441] <= 16'b0000000000000010;
        weights1[33442] <= 16'b1111111111010100;
        weights1[33443] <= 16'b1111111101101101;
        weights1[33444] <= 16'b1111111110110000;
        weights1[33445] <= 16'b1111111111101111;
        weights1[33446] <= 16'b0000000000000111;
        weights1[33447] <= 16'b1111111111101111;
        weights1[33448] <= 16'b0000000000001011;
        weights1[33449] <= 16'b0000000000010000;
        weights1[33450] <= 16'b0000000000000011;
        weights1[33451] <= 16'b1111111111111111;
        weights1[33452] <= 16'b1111111111111001;
        weights1[33453] <= 16'b0000000000011110;
        weights1[33454] <= 16'b1111111111111110;
        weights1[33455] <= 16'b1111111111101111;
        weights1[33456] <= 16'b1111111111101110;
        weights1[33457] <= 16'b1111111111100011;
        weights1[33458] <= 16'b1111111111111000;
        weights1[33459] <= 16'b1111111111111111;
        weights1[33460] <= 16'b0000000000010011;
        weights1[33461] <= 16'b0000000000001010;
        weights1[33462] <= 16'b0000000000010000;
        weights1[33463] <= 16'b0000000000000001;
        weights1[33464] <= 16'b1111111111110100;
        weights1[33465] <= 16'b0000000000000100;
        weights1[33466] <= 16'b0000000000000100;
        weights1[33467] <= 16'b1111111111111001;
        weights1[33468] <= 16'b1111111111110110;
        weights1[33469] <= 16'b1111111111110011;
        weights1[33470] <= 16'b1111111111011110;
        weights1[33471] <= 16'b1111111110101100;
        weights1[33472] <= 16'b1111111111001111;
        weights1[33473] <= 16'b1111111111100111;
        weights1[33474] <= 16'b0000000000001101;
        weights1[33475] <= 16'b0000000000001010;
        weights1[33476] <= 16'b0000000000000011;
        weights1[33477] <= 16'b1111111111111101;
        weights1[33478] <= 16'b0000000000010010;
        weights1[33479] <= 16'b1111111111101101;
        weights1[33480] <= 16'b0000000000000010;
        weights1[33481] <= 16'b0000000000001111;
        weights1[33482] <= 16'b1111111111101101;
        weights1[33483] <= 16'b1111111111100110;
        weights1[33484] <= 16'b1111111111100010;
        weights1[33485] <= 16'b1111111111101001;
        weights1[33486] <= 16'b1111111111111001;
        weights1[33487] <= 16'b0000000000000100;
        weights1[33488] <= 16'b0000000000010100;
        weights1[33489] <= 16'b0000000000001111;
        weights1[33490] <= 16'b0000000000000111;
        weights1[33491] <= 16'b0000000000000011;
        weights1[33492] <= 16'b0000000000010100;
        weights1[33493] <= 16'b0000000000000111;
        weights1[33494] <= 16'b0000000000011010;
        weights1[33495] <= 16'b0000000000000000;
        weights1[33496] <= 16'b1111111111111010;
        weights1[33497] <= 16'b1111111111101111;
        weights1[33498] <= 16'b1111111111110011;
        weights1[33499] <= 16'b0000000000000001;
        weights1[33500] <= 16'b1111111111110111;
        weights1[33501] <= 16'b1111111111101010;
        weights1[33502] <= 16'b0000000000000010;
        weights1[33503] <= 16'b1111111111111100;
        weights1[33504] <= 16'b1111111111101101;
        weights1[33505] <= 16'b1111111111111000;
        weights1[33506] <= 16'b1111111111100011;
        weights1[33507] <= 16'b0000000000001111;
        weights1[33508] <= 16'b1111111111101001;
        weights1[33509] <= 16'b1111111111101111;
        weights1[33510] <= 16'b1111111111110001;
        weights1[33511] <= 16'b1111111111101101;
        weights1[33512] <= 16'b1111111111101101;
        weights1[33513] <= 16'b1111111111101100;
        weights1[33514] <= 16'b1111111111110011;
        weights1[33515] <= 16'b1111111111111101;
        weights1[33516] <= 16'b0000000000001101;
        weights1[33517] <= 16'b0000000000000111;
        weights1[33518] <= 16'b0000000000000011;
        weights1[33519] <= 16'b0000000000001011;
        weights1[33520] <= 16'b0000000000010001;
        weights1[33521] <= 16'b0000000000010100;
        weights1[33522] <= 16'b1111111111111110;
        weights1[33523] <= 16'b0000000000000110;
        weights1[33524] <= 16'b1111111111101101;
        weights1[33525] <= 16'b0000000000001011;
        weights1[33526] <= 16'b0000000000010101;
        weights1[33527] <= 16'b0000000000010100;
        weights1[33528] <= 16'b0000000000000010;
        weights1[33529] <= 16'b0000000000000100;
        weights1[33530] <= 16'b1111111111101101;
        weights1[33531] <= 16'b0000000000001101;
        weights1[33532] <= 16'b0000000000000001;
        weights1[33533] <= 16'b1111111111111001;
        weights1[33534] <= 16'b1111111111101100;
        weights1[33535] <= 16'b1111111111010010;
        weights1[33536] <= 16'b1111111111110010;
        weights1[33537] <= 16'b1111111111110100;
        weights1[33538] <= 16'b1111111111010101;
        weights1[33539] <= 16'b1111111111100010;
        weights1[33540] <= 16'b1111111111101010;
        weights1[33541] <= 16'b1111111111101110;
        weights1[33542] <= 16'b1111111111110110;
        weights1[33543] <= 16'b1111111111111100;
        weights1[33544] <= 16'b0000000000000111;
        weights1[33545] <= 16'b0000000000001001;
        weights1[33546] <= 16'b0000000000000010;
        weights1[33547] <= 16'b0000000000000111;
        weights1[33548] <= 16'b1111111111101101;
        weights1[33549] <= 16'b0000000000000010;
        weights1[33550] <= 16'b0000000000011101;
        weights1[33551] <= 16'b1111111111110100;
        weights1[33552] <= 16'b0000000000100100;
        weights1[33553] <= 16'b0000000000110001;
        weights1[33554] <= 16'b0000000000001011;
        weights1[33555] <= 16'b1111111111111111;
        weights1[33556] <= 16'b0000000000001010;
        weights1[33557] <= 16'b0000000000011101;
        weights1[33558] <= 16'b0000000000010111;
        weights1[33559] <= 16'b0000000000000101;
        weights1[33560] <= 16'b1111111111111010;
        weights1[33561] <= 16'b0000000000000101;
        weights1[33562] <= 16'b0000000000010011;
        weights1[33563] <= 16'b1111111111111000;
        weights1[33564] <= 16'b1111111111101000;
        weights1[33565] <= 16'b1111111111101100;
        weights1[33566] <= 16'b1111111111101011;
        weights1[33567] <= 16'b1111111111101101;
        weights1[33568] <= 16'b1111111111100101;
        weights1[33569] <= 16'b1111111111101100;
        weights1[33570] <= 16'b1111111111111010;
        weights1[33571] <= 16'b1111111111111100;
        weights1[33572] <= 16'b0000000000000101;
        weights1[33573] <= 16'b0000000000000010;
        weights1[33574] <= 16'b1111111111111100;
        weights1[33575] <= 16'b0000000000000100;
        weights1[33576] <= 16'b0000000000001111;
        weights1[33577] <= 16'b0000000000000100;
        weights1[33578] <= 16'b0000000000100010;
        weights1[33579] <= 16'b0000000000100111;
        weights1[33580] <= 16'b0000000000000001;
        weights1[33581] <= 16'b1111111111111111;
        weights1[33582] <= 16'b0000000000100001;
        weights1[33583] <= 16'b0000000000000000;
        weights1[33584] <= 16'b0000000000000101;
        weights1[33585] <= 16'b0000000000010000;
        weights1[33586] <= 16'b0000000000001101;
        weights1[33587] <= 16'b0000000000011001;
        weights1[33588] <= 16'b0000000000000001;
        weights1[33589] <= 16'b0000000000101010;
        weights1[33590] <= 16'b0000000000000001;
        weights1[33591] <= 16'b0000000000000001;
        weights1[33592] <= 16'b1111111111101110;
        weights1[33593] <= 16'b0000000000000101;
        weights1[33594] <= 16'b1111111111110010;
        weights1[33595] <= 16'b1111111111110111;
        weights1[33596] <= 16'b1111111111110010;
        weights1[33597] <= 16'b1111111111111000;
        weights1[33598] <= 16'b1111111111111111;
        weights1[33599] <= 16'b1111111111111111;
        weights1[33600] <= 16'b1111111111111011;
        weights1[33601] <= 16'b0000000000000111;
        weights1[33602] <= 16'b1111111111110011;
        weights1[33603] <= 16'b0000000000000011;
        weights1[33604] <= 16'b0000000000001111;
        weights1[33605] <= 16'b0000000000011101;
        weights1[33606] <= 16'b0000000000100011;
        weights1[33607] <= 16'b0000000000001101;
        weights1[33608] <= 16'b0000000000011011;
        weights1[33609] <= 16'b0000000000100010;
        weights1[33610] <= 16'b0000000000011111;
        weights1[33611] <= 16'b0000000000010010;
        weights1[33612] <= 16'b0000000000000100;
        weights1[33613] <= 16'b1111111111101010;
        weights1[33614] <= 16'b0000000000001010;
        weights1[33615] <= 16'b1111111111100010;
        weights1[33616] <= 16'b1111111111100001;
        weights1[33617] <= 16'b0000000000001000;
        weights1[33618] <= 16'b1111111111100000;
        weights1[33619] <= 16'b1111111111101000;
        weights1[33620] <= 16'b1111111111110001;
        weights1[33621] <= 16'b0000000000000100;
        weights1[33622] <= 16'b1111111111110101;
        weights1[33623] <= 16'b1111111111110111;
        weights1[33624] <= 16'b1111111111111000;
        weights1[33625] <= 16'b1111111111111001;
        weights1[33626] <= 16'b1111111111111101;
        weights1[33627] <= 16'b0000000000000001;
        weights1[33628] <= 16'b1111111111111111;
        weights1[33629] <= 16'b0000000000000000;
        weights1[33630] <= 16'b0000000000000011;
        weights1[33631] <= 16'b0000000000001010;
        weights1[33632] <= 16'b0000000000001101;
        weights1[33633] <= 16'b0000000000000111;
        weights1[33634] <= 16'b0000000000100011;
        weights1[33635] <= 16'b0000000000011000;
        weights1[33636] <= 16'b0000000000001101;
        weights1[33637] <= 16'b0000000000000010;
        weights1[33638] <= 16'b0000000000001010;
        weights1[33639] <= 16'b0000000000000101;
        weights1[33640] <= 16'b0000000000001011;
        weights1[33641] <= 16'b1111111111111101;
        weights1[33642] <= 16'b0000000000001011;
        weights1[33643] <= 16'b1111111111110010;
        weights1[33644] <= 16'b1111111111110000;
        weights1[33645] <= 16'b1111111111010110;
        weights1[33646] <= 16'b1111111111110100;
        weights1[33647] <= 16'b1111111111110010;
        weights1[33648] <= 16'b1111111111101011;
        weights1[33649] <= 16'b0000000000000110;
        weights1[33650] <= 16'b1111111111110000;
        weights1[33651] <= 16'b1111111111111000;
        weights1[33652] <= 16'b1111111111110011;
        weights1[33653] <= 16'b1111111111110110;
        weights1[33654] <= 16'b1111111111111000;
        weights1[33655] <= 16'b1111111111111011;
        weights1[33656] <= 16'b0000000000000000;
        weights1[33657] <= 16'b1111111111111001;
        weights1[33658] <= 16'b1111111111111111;
        weights1[33659] <= 16'b0000000000000000;
        weights1[33660] <= 16'b0000000000000001;
        weights1[33661] <= 16'b0000000000001011;
        weights1[33662] <= 16'b1111111111111111;
        weights1[33663] <= 16'b0000000000001101;
        weights1[33664] <= 16'b0000000000011011;
        weights1[33665] <= 16'b0000000000001000;
        weights1[33666] <= 16'b0000000000000100;
        weights1[33667] <= 16'b0000000000011101;
        weights1[33668] <= 16'b1111111111110110;
        weights1[33669] <= 16'b0000000000000010;
        weights1[33670] <= 16'b0000000000000111;
        weights1[33671] <= 16'b0000000000001001;
        weights1[33672] <= 16'b0000000000000011;
        weights1[33673] <= 16'b0000000000000001;
        weights1[33674] <= 16'b1111111111101111;
        weights1[33675] <= 16'b0000000000010000;
        weights1[33676] <= 16'b1111111111101010;
        weights1[33677] <= 16'b1111111111110001;
        weights1[33678] <= 16'b1111111111100110;
        weights1[33679] <= 16'b1111111111101011;
        weights1[33680] <= 16'b1111111111110001;
        weights1[33681] <= 16'b1111111111110111;
        weights1[33682] <= 16'b1111111111111101;
        weights1[33683] <= 16'b1111111111111101;
        weights1[33684] <= 16'b1111111111111110;
        weights1[33685] <= 16'b1111111111111110;
        weights1[33686] <= 16'b1111111111111110;
        weights1[33687] <= 16'b1111111111111101;
        weights1[33688] <= 16'b1111111111110011;
        weights1[33689] <= 16'b1111111111110011;
        weights1[33690] <= 16'b1111111111110000;
        weights1[33691] <= 16'b1111111111110100;
        weights1[33692] <= 16'b0000000000000111;
        weights1[33693] <= 16'b1111111111111010;
        weights1[33694] <= 16'b1111111111111100;
        weights1[33695] <= 16'b0000000000000010;
        weights1[33696] <= 16'b0000000000011000;
        weights1[33697] <= 16'b1111111111111111;
        weights1[33698] <= 16'b1111111111101001;
        weights1[33699] <= 16'b1111111111010101;
        weights1[33700] <= 16'b1111111111011100;
        weights1[33701] <= 16'b1111111111011001;
        weights1[33702] <= 16'b1111111111011010;
        weights1[33703] <= 16'b1111111111001101;
        weights1[33704] <= 16'b1111111111100010;
        weights1[33705] <= 16'b1111111111011011;
        weights1[33706] <= 16'b1111111111011111;
        weights1[33707] <= 16'b1111111111101101;
        weights1[33708] <= 16'b1111111111110000;
        weights1[33709] <= 16'b1111111111110110;
        weights1[33710] <= 16'b0000000000000110;
        weights1[33711] <= 16'b0000000000000010;
        weights1[33712] <= 16'b0000000000000001;
        weights1[33713] <= 16'b0000000000000001;
        weights1[33714] <= 16'b0000000000000001;
        weights1[33715] <= 16'b0000000000001000;
        weights1[33716] <= 16'b0000000000000000;
        weights1[33717] <= 16'b1111111111110001;
        weights1[33718] <= 16'b1111111111100100;
        weights1[33719] <= 16'b1111111111010110;
        weights1[33720] <= 16'b1111111111001101;
        weights1[33721] <= 16'b1111111111001101;
        weights1[33722] <= 16'b1111111111011110;
        weights1[33723] <= 16'b0000000000001000;
        weights1[33724] <= 16'b0000000000101100;
        weights1[33725] <= 16'b0000000000101100;
        weights1[33726] <= 16'b0000000000011100;
        weights1[33727] <= 16'b0000000000001011;
        weights1[33728] <= 16'b1111111111100010;
        weights1[33729] <= 16'b1111111110110001;
        weights1[33730] <= 16'b1111111110010101;
        weights1[33731] <= 16'b1111111110110111;
        weights1[33732] <= 16'b1111111111011011;
        weights1[33733] <= 16'b1111111111101101;
        weights1[33734] <= 16'b0000000000000001;
        weights1[33735] <= 16'b0000000000001000;
        weights1[33736] <= 16'b0000000000000101;
        weights1[33737] <= 16'b0000000000000100;
        weights1[33738] <= 16'b0000000000000101;
        weights1[33739] <= 16'b0000000000000101;
        weights1[33740] <= 16'b0000000000000001;
        weights1[33741] <= 16'b0000000000000001;
        weights1[33742] <= 16'b0000000000000011;
        weights1[33743] <= 16'b0000000000001110;
        weights1[33744] <= 16'b0000000000000010;
        weights1[33745] <= 16'b1111111111101000;
        weights1[33746] <= 16'b1111111111011000;
        weights1[33747] <= 16'b1111111111000111;
        weights1[33748] <= 16'b1111111110111000;
        weights1[33749] <= 16'b1111111111001101;
        weights1[33750] <= 16'b1111111111101101;
        weights1[33751] <= 16'b0000000000101101;
        weights1[33752] <= 16'b0000000000110001;
        weights1[33753] <= 16'b0000000000101111;
        weights1[33754] <= 16'b0000000000010000;
        weights1[33755] <= 16'b1111111111110101;
        weights1[33756] <= 16'b1111111110100110;
        weights1[33757] <= 16'b1111111110000011;
        weights1[33758] <= 16'b1111111110000000;
        weights1[33759] <= 16'b1111111110111001;
        weights1[33760] <= 16'b1111111111100010;
        weights1[33761] <= 16'b0000000000000111;
        weights1[33762] <= 16'b0000000000001000;
        weights1[33763] <= 16'b0000000000001101;
        weights1[33764] <= 16'b0000000000011001;
        weights1[33765] <= 16'b0000000000001001;
        weights1[33766] <= 16'b0000000000000011;
        weights1[33767] <= 16'b0000000000000001;
        weights1[33768] <= 16'b0000000000000010;
        weights1[33769] <= 16'b0000000000000100;
        weights1[33770] <= 16'b0000000000001001;
        weights1[33771] <= 16'b0000000000001100;
        weights1[33772] <= 16'b0000000000000011;
        weights1[33773] <= 16'b1111111111101010;
        weights1[33774] <= 16'b1111111111001010;
        weights1[33775] <= 16'b1111111110110000;
        weights1[33776] <= 16'b1111111110100101;
        weights1[33777] <= 16'b1111111111001011;
        weights1[33778] <= 16'b1111111111111011;
        weights1[33779] <= 16'b0000000000110100;
        weights1[33780] <= 16'b0000000000100110;
        weights1[33781] <= 16'b0000000000110100;
        weights1[33782] <= 16'b0000000000011010;
        weights1[33783] <= 16'b1111111111011011;
        weights1[33784] <= 16'b1111111101100101;
        weights1[33785] <= 16'b1111111101001100;
        weights1[33786] <= 16'b1111111110010001;
        weights1[33787] <= 16'b1111111111011011;
        weights1[33788] <= 16'b1111111111101111;
        weights1[33789] <= 16'b0000000000000110;
        weights1[33790] <= 16'b0000000000010110;
        weights1[33791] <= 16'b0000000000100000;
        weights1[33792] <= 16'b0000000000001111;
        weights1[33793] <= 16'b0000000000000111;
        weights1[33794] <= 16'b0000000000000000;
        weights1[33795] <= 16'b1111111111111100;
        weights1[33796] <= 16'b0000000000000000;
        weights1[33797] <= 16'b0000000000000011;
        weights1[33798] <= 16'b0000000000010000;
        weights1[33799] <= 16'b0000000000010100;
        weights1[33800] <= 16'b0000000000000100;
        weights1[33801] <= 16'b1111111111101100;
        weights1[33802] <= 16'b1111111111001010;
        weights1[33803] <= 16'b1111111110011000;
        weights1[33804] <= 16'b1111111110011000;
        weights1[33805] <= 16'b1111111111010111;
        weights1[33806] <= 16'b0000000000000111;
        weights1[33807] <= 16'b0000000000110110;
        weights1[33808] <= 16'b0000000000101011;
        weights1[33809] <= 16'b0000000000111000;
        weights1[33810] <= 16'b0000000000010011;
        weights1[33811] <= 16'b1111111110111001;
        weights1[33812] <= 16'b1111111100011101;
        weights1[33813] <= 16'b1111111101011001;
        weights1[33814] <= 16'b1111111111000000;
        weights1[33815] <= 16'b0000000000000000;
        weights1[33816] <= 16'b0000000000100100;
        weights1[33817] <= 16'b0000000000011100;
        weights1[33818] <= 16'b0000000000110110;
        weights1[33819] <= 16'b0000000000011111;
        weights1[33820] <= 16'b0000000000001101;
        weights1[33821] <= 16'b1111111111111101;
        weights1[33822] <= 16'b1111111111101101;
        weights1[33823] <= 16'b1111111111110001;
        weights1[33824] <= 16'b0000000000000010;
        weights1[33825] <= 16'b0000000000001010;
        weights1[33826] <= 16'b0000000000010100;
        weights1[33827] <= 16'b0000000000011010;
        weights1[33828] <= 16'b0000000000000101;
        weights1[33829] <= 16'b1111111111101010;
        weights1[33830] <= 16'b1111111110111011;
        weights1[33831] <= 16'b1111111110001111;
        weights1[33832] <= 16'b1111111110001100;
        weights1[33833] <= 16'b1111111111000111;
        weights1[33834] <= 16'b0000000000010101;
        weights1[33835] <= 16'b0000000000111101;
        weights1[33836] <= 16'b0000000000111011;
        weights1[33837] <= 16'b0000000000111100;
        weights1[33838] <= 16'b1111111111101011;
        weights1[33839] <= 16'b1111111101111010;
        weights1[33840] <= 16'b1111111100011001;
        weights1[33841] <= 16'b1111111101101111;
        weights1[33842] <= 16'b1111111111100000;
        weights1[33843] <= 16'b0000000000101111;
        weights1[33844] <= 16'b0000000000101011;
        weights1[33845] <= 16'b0000000000010110;
        weights1[33846] <= 16'b0000000000011100;
        weights1[33847] <= 16'b0000000000000110;
        weights1[33848] <= 16'b0000000000001110;
        weights1[33849] <= 16'b1111111111110010;
        weights1[33850] <= 16'b1111111111101000;
        weights1[33851] <= 16'b1111111111101110;
        weights1[33852] <= 16'b0000000000000110;
        weights1[33853] <= 16'b0000000000001000;
        weights1[33854] <= 16'b0000000000011111;
        weights1[33855] <= 16'b0000000000010111;
        weights1[33856] <= 16'b0000000000010100;
        weights1[33857] <= 16'b1111111111110110;
        weights1[33858] <= 16'b1111111111001000;
        weights1[33859] <= 16'b1111111110001100;
        weights1[33860] <= 16'b1111111101110101;
        weights1[33861] <= 16'b0000000000000000;
        weights1[33862] <= 16'b0000000000111100;
        weights1[33863] <= 16'b0000000000100010;
        weights1[33864] <= 16'b0000000001000011;
        weights1[33865] <= 16'b0000000000110101;
        weights1[33866] <= 16'b1111111111100101;
        weights1[33867] <= 16'b1111111101011110;
        weights1[33868] <= 16'b1111111100001110;
        weights1[33869] <= 16'b1111111111011010;
        weights1[33870] <= 16'b0000000001000011;
        weights1[33871] <= 16'b0000000000101000;
        weights1[33872] <= 16'b0000000000111011;
        weights1[33873] <= 16'b0000000000010110;
        weights1[33874] <= 16'b0000000000001010;
        weights1[33875] <= 16'b0000000000100111;
        weights1[33876] <= 16'b0000000000000110;
        weights1[33877] <= 16'b1111111111011101;
        weights1[33878] <= 16'b1111111111100100;
        weights1[33879] <= 16'b1111111111100011;
        weights1[33880] <= 16'b0000000000000001;
        weights1[33881] <= 16'b0000000000001101;
        weights1[33882] <= 16'b0000000000011110;
        weights1[33883] <= 16'b0000000000011000;
        weights1[33884] <= 16'b0000000000010000;
        weights1[33885] <= 16'b0000000000000110;
        weights1[33886] <= 16'b1111111111000011;
        weights1[33887] <= 16'b1111111101111110;
        weights1[33888] <= 16'b1111111101110000;
        weights1[33889] <= 16'b0000000000000000;
        weights1[33890] <= 16'b0000000000010100;
        weights1[33891] <= 16'b0000000000100101;
        weights1[33892] <= 16'b0000000000100111;
        weights1[33893] <= 16'b0000000000011100;
        weights1[33894] <= 16'b1111111111111101;
        weights1[33895] <= 16'b1111111100111111;
        weights1[33896] <= 16'b1111111101100011;
        weights1[33897] <= 16'b0000000000100011;
        weights1[33898] <= 16'b0000000000111000;
        weights1[33899] <= 16'b0000000000010001;
        weights1[33900] <= 16'b0000000000010010;
        weights1[33901] <= 16'b0000000000011011;
        weights1[33902] <= 16'b0000000000011000;
        weights1[33903] <= 16'b1111111111111100;
        weights1[33904] <= 16'b1111111111010000;
        weights1[33905] <= 16'b1111111111010011;
        weights1[33906] <= 16'b1111111111010100;
        weights1[33907] <= 16'b1111111111011001;
        weights1[33908] <= 16'b0000000000000101;
        weights1[33909] <= 16'b0000000000001011;
        weights1[33910] <= 16'b0000000000011111;
        weights1[33911] <= 16'b0000000000011000;
        weights1[33912] <= 16'b0000000000001110;
        weights1[33913] <= 16'b0000000000010011;
        weights1[33914] <= 16'b1111111111011110;
        weights1[33915] <= 16'b1111111110101001;
        weights1[33916] <= 16'b1111111110110010;
        weights1[33917] <= 16'b1111111111100010;
        weights1[33918] <= 16'b0000000000011011;
        weights1[33919] <= 16'b0000000000011000;
        weights1[33920] <= 16'b0000000000101010;
        weights1[33921] <= 16'b0000000000000001;
        weights1[33922] <= 16'b1111111111100001;
        weights1[33923] <= 16'b1111111101001000;
        weights1[33924] <= 16'b1111111111000101;
        weights1[33925] <= 16'b0000000000010100;
        weights1[33926] <= 16'b0000000000101100;
        weights1[33927] <= 16'b0000000000001111;
        weights1[33928] <= 16'b0000000000010001;
        weights1[33929] <= 16'b0000000000010110;
        weights1[33930] <= 16'b0000000000000100;
        weights1[33931] <= 16'b1111111111101010;
        weights1[33932] <= 16'b1111111110111101;
        weights1[33933] <= 16'b1111111111000110;
        weights1[33934] <= 16'b1111111111001001;
        weights1[33935] <= 16'b1111111111100010;
        weights1[33936] <= 16'b0000000000000100;
        weights1[33937] <= 16'b0000000000001011;
        weights1[33938] <= 16'b0000000000010000;
        weights1[33939] <= 16'b0000000000011110;
        weights1[33940] <= 16'b0000000000011010;
        weights1[33941] <= 16'b0000000000001100;
        weights1[33942] <= 16'b1111111111110110;
        weights1[33943] <= 16'b1111111111010011;
        weights1[33944] <= 16'b1111111110110100;
        weights1[33945] <= 16'b1111111111111011;
        weights1[33946] <= 16'b0000000000001000;
        weights1[33947] <= 16'b0000000000011101;
        weights1[33948] <= 16'b0000000000100010;
        weights1[33949] <= 16'b0000000000010100;
        weights1[33950] <= 16'b1111111111010111;
        weights1[33951] <= 16'b1111111110010000;
        weights1[33952] <= 16'b1111111111101111;
        weights1[33953] <= 16'b0000000000011011;
        weights1[33954] <= 16'b0000000000100111;
        weights1[33955] <= 16'b0000000000010100;
        weights1[33956] <= 16'b0000000000001001;
        weights1[33957] <= 16'b0000000000011110;
        weights1[33958] <= 16'b1111111111110010;
        weights1[33959] <= 16'b1111111111010011;
        weights1[33960] <= 16'b1111111110111100;
        weights1[33961] <= 16'b1111111111010110;
        weights1[33962] <= 16'b1111111111100011;
        weights1[33963] <= 16'b1111111111101100;
        weights1[33964] <= 16'b0000000000000110;
        weights1[33965] <= 16'b0000000000010110;
        weights1[33966] <= 16'b0000000000011110;
        weights1[33967] <= 16'b0000000000001000;
        weights1[33968] <= 16'b0000000000011000;
        weights1[33969] <= 16'b0000000000010101;
        weights1[33970] <= 16'b1111111111111010;
        weights1[33971] <= 16'b1111111111010010;
        weights1[33972] <= 16'b1111111111011011;
        weights1[33973] <= 16'b1111111111011111;
        weights1[33974] <= 16'b1111111111100001;
        weights1[33975] <= 16'b0000000000010010;
        weights1[33976] <= 16'b0000000000011100;
        weights1[33977] <= 16'b0000000000000110;
        weights1[33978] <= 16'b1111111111001100;
        weights1[33979] <= 16'b1111111111000110;
        weights1[33980] <= 16'b1111111111111001;
        weights1[33981] <= 16'b0000000000100001;
        weights1[33982] <= 16'b0000000000001101;
        weights1[33983] <= 16'b0000000000001111;
        weights1[33984] <= 16'b1111111111111110;
        weights1[33985] <= 16'b1111111111110100;
        weights1[33986] <= 16'b1111111111011101;
        weights1[33987] <= 16'b1111111110110111;
        weights1[33988] <= 16'b1111111111010101;
        weights1[33989] <= 16'b1111111111111011;
        weights1[33990] <= 16'b1111111111111111;
        weights1[33991] <= 16'b0000000000001010;
        weights1[33992] <= 16'b0000000000000001;
        weights1[33993] <= 16'b0000000000000000;
        weights1[33994] <= 16'b0000000000010111;
        weights1[33995] <= 16'b0000000000000101;
        weights1[33996] <= 16'b0000000000010011;
        weights1[33997] <= 16'b0000000000011110;
        weights1[33998] <= 16'b1111111111110010;
        weights1[33999] <= 16'b1111111111011100;
        weights1[34000] <= 16'b1111111111010001;
        weights1[34001] <= 16'b0000000000001001;
        weights1[34002] <= 16'b1111111111101110;
        weights1[34003] <= 16'b0000000000101011;
        weights1[34004] <= 16'b0000000000010000;
        weights1[34005] <= 16'b1111111111110010;
        weights1[34006] <= 16'b1111111111101000;
        weights1[34007] <= 16'b1111111111011110;
        weights1[34008] <= 16'b0000000000001110;
        weights1[34009] <= 16'b0000000000001111;
        weights1[34010] <= 16'b0000000000001100;
        weights1[34011] <= 16'b0000000000001011;
        weights1[34012] <= 16'b1111111111110000;
        weights1[34013] <= 16'b1111111111111110;
        weights1[34014] <= 16'b1111111111011000;
        weights1[34015] <= 16'b1111111111011000;
        weights1[34016] <= 16'b1111111111111011;
        weights1[34017] <= 16'b0000000000001110;
        weights1[34018] <= 16'b0000000000010010;
        weights1[34019] <= 16'b0000000000010111;
        weights1[34020] <= 16'b0000000000000101;
        weights1[34021] <= 16'b1111111111111111;
        weights1[34022] <= 16'b0000000000001001;
        weights1[34023] <= 16'b1111111111110010;
        weights1[34024] <= 16'b1111111111111001;
        weights1[34025] <= 16'b0000000000100011;
        weights1[34026] <= 16'b0000000000000101;
        weights1[34027] <= 16'b1111111111111110;
        weights1[34028] <= 16'b1111111111111011;
        weights1[34029] <= 16'b1111111111101111;
        weights1[34030] <= 16'b1111111111110110;
        weights1[34031] <= 16'b0000000000000000;
        weights1[34032] <= 16'b0000000000001001;
        weights1[34033] <= 16'b1111111111111100;
        weights1[34034] <= 16'b1111111111111011;
        weights1[34035] <= 16'b1111111111100101;
        weights1[34036] <= 16'b0000000000011000;
        weights1[34037] <= 16'b0000000000000110;
        weights1[34038] <= 16'b1111111111111010;
        weights1[34039] <= 16'b0000000000010000;
        weights1[34040] <= 16'b1111111111101110;
        weights1[34041] <= 16'b1111111111110011;
        weights1[34042] <= 16'b1111111111001000;
        weights1[34043] <= 16'b0000000000000001;
        weights1[34044] <= 16'b0000000000001011;
        weights1[34045] <= 16'b0000000000010001;
        weights1[34046] <= 16'b0000000000100010;
        weights1[34047] <= 16'b0000000000100110;
        weights1[34048] <= 16'b1111111111111011;
        weights1[34049] <= 16'b1111111111111100;
        weights1[34050] <= 16'b0000000000010000;
        weights1[34051] <= 16'b0000000000010101;
        weights1[34052] <= 16'b0000000000011001;
        weights1[34053] <= 16'b1111111111111011;
        weights1[34054] <= 16'b0000000000001100;
        weights1[34055] <= 16'b0000000000001101;
        weights1[34056] <= 16'b1111111111101111;
        weights1[34057] <= 16'b1111111111101001;
        weights1[34058] <= 16'b1111111111111110;
        weights1[34059] <= 16'b0000000000000111;
        weights1[34060] <= 16'b0000000000000011;
        weights1[34061] <= 16'b0000000000000011;
        weights1[34062] <= 16'b1111111111110110;
        weights1[34063] <= 16'b0000000000001000;
        weights1[34064] <= 16'b0000000000001010;
        weights1[34065] <= 16'b0000000000000001;
        weights1[34066] <= 16'b1111111111111110;
        weights1[34067] <= 16'b1111111111110110;
        weights1[34068] <= 16'b1111111111101100;
        weights1[34069] <= 16'b1111111111101110;
        weights1[34070] <= 16'b1111111111101110;
        weights1[34071] <= 16'b0000000000001001;
        weights1[34072] <= 16'b0000000000011111;
        weights1[34073] <= 16'b0000000000001000;
        weights1[34074] <= 16'b0000000000001001;
        weights1[34075] <= 16'b0000000000011011;
        weights1[34076] <= 16'b1111111111111001;
        weights1[34077] <= 16'b0000000000000110;
        weights1[34078] <= 16'b0000000000000110;
        weights1[34079] <= 16'b1111111111111111;
        weights1[34080] <= 16'b0000000000001111;
        weights1[34081] <= 16'b1111111111110100;
        weights1[34082] <= 16'b1111111111111100;
        weights1[34083] <= 16'b0000000000001101;
        weights1[34084] <= 16'b0000000000001100;
        weights1[34085] <= 16'b0000000000011001;
        weights1[34086] <= 16'b1111111111111111;
        weights1[34087] <= 16'b0000000000000100;
        weights1[34088] <= 16'b0000000000000110;
        weights1[34089] <= 16'b0000000000000100;
        weights1[34090] <= 16'b1111111111101111;
        weights1[34091] <= 16'b1111111111110011;
        weights1[34092] <= 16'b1111111111111000;
        weights1[34093] <= 16'b0000000000000100;
        weights1[34094] <= 16'b1111111111110111;
        weights1[34095] <= 16'b1111111111111001;
        weights1[34096] <= 16'b0000000000000111;
        weights1[34097] <= 16'b1111111111101101;
        weights1[34098] <= 16'b0000000000010000;
        weights1[34099] <= 16'b0000000000001000;
        weights1[34100] <= 16'b0000000000001111;
        weights1[34101] <= 16'b0000000000000011;
        weights1[34102] <= 16'b0000000000010111;
        weights1[34103] <= 16'b0000000000010110;
        weights1[34104] <= 16'b1111111111110001;
        weights1[34105] <= 16'b1111111111111111;
        weights1[34106] <= 16'b1111111111111100;
        weights1[34107] <= 16'b1111111111110011;
        weights1[34108] <= 16'b1111111111111111;
        weights1[34109] <= 16'b0000000000011001;
        weights1[34110] <= 16'b0000000000000001;
        weights1[34111] <= 16'b0000000000001001;
        weights1[34112] <= 16'b0000000000000100;
        weights1[34113] <= 16'b1111111111111100;
        weights1[34114] <= 16'b1111111111111011;
        weights1[34115] <= 16'b0000000000001111;
        weights1[34116] <= 16'b0000000000001100;
        weights1[34117] <= 16'b1111111111110110;
        weights1[34118] <= 16'b0000000000001111;
        weights1[34119] <= 16'b0000000000010111;
        weights1[34120] <= 16'b0000000000001100;
        weights1[34121] <= 16'b1111111111111011;
        weights1[34122] <= 16'b1111111111110011;
        weights1[34123] <= 16'b0000000000011000;
        weights1[34124] <= 16'b0000000000000010;
        weights1[34125] <= 16'b0000000000010010;
        weights1[34126] <= 16'b0000000000000000;
        weights1[34127] <= 16'b0000000000001111;
        weights1[34128] <= 16'b0000000000001110;
        weights1[34129] <= 16'b0000000000001110;
        weights1[34130] <= 16'b0000000000010100;
        weights1[34131] <= 16'b0000000000000000;
        weights1[34132] <= 16'b0000000000000100;
        weights1[34133] <= 16'b1111111111111000;
        weights1[34134] <= 16'b0000000000000100;
        weights1[34135] <= 16'b0000000000001000;
        weights1[34136] <= 16'b0000000000000101;
        weights1[34137] <= 16'b0000000000000100;
        weights1[34138] <= 16'b1111111111111110;
        weights1[34139] <= 16'b0000000000000011;
        weights1[34140] <= 16'b0000000000000010;
        weights1[34141] <= 16'b0000000000000111;
        weights1[34142] <= 16'b0000000000100011;
        weights1[34143] <= 16'b1111111111111111;
        weights1[34144] <= 16'b0000000000000110;
        weights1[34145] <= 16'b0000000000001111;
        weights1[34146] <= 16'b0000000000001011;
        weights1[34147] <= 16'b0000000000000100;
        weights1[34148] <= 16'b1111111111111010;
        weights1[34149] <= 16'b0000000000000001;
        weights1[34150] <= 16'b1111111111111001;
        weights1[34151] <= 16'b0000000000000100;
        weights1[34152] <= 16'b0000000000001110;
        weights1[34153] <= 16'b0000000000000111;
        weights1[34154] <= 16'b0000000000010111;
        weights1[34155] <= 16'b0000000000001010;
        weights1[34156] <= 16'b1111111111110011;
        weights1[34157] <= 16'b1111111111111111;
        weights1[34158] <= 16'b1111111111111010;
        weights1[34159] <= 16'b1111111111111111;
        weights1[34160] <= 16'b1111111111111010;
        weights1[34161] <= 16'b1111111111111010;
        weights1[34162] <= 16'b0000000000001011;
        weights1[34163] <= 16'b0000000000000010;
        weights1[34164] <= 16'b0000000000000100;
        weights1[34165] <= 16'b0000000000001001;
        weights1[34166] <= 16'b0000000000011101;
        weights1[34167] <= 16'b1111111111111010;
        weights1[34168] <= 16'b0000000000000111;
        weights1[34169] <= 16'b1111111111110111;
        weights1[34170] <= 16'b1111111111110111;
        weights1[34171] <= 16'b1111111111111000;
        weights1[34172] <= 16'b1111111111111011;
        weights1[34173] <= 16'b1111111111111111;
        weights1[34174] <= 16'b0000000000001001;
        weights1[34175] <= 16'b0000000000001111;
        weights1[34176] <= 16'b1111111111111110;
        weights1[34177] <= 16'b1111111111101011;
        weights1[34178] <= 16'b1111111111110111;
        weights1[34179] <= 16'b0000000000000100;
        weights1[34180] <= 16'b1111111111111010;
        weights1[34181] <= 16'b0000000000000111;
        weights1[34182] <= 16'b0000000000010011;
        weights1[34183] <= 16'b0000000000000111;
        weights1[34184] <= 16'b0000000000100111;
        weights1[34185] <= 16'b1111111111111010;
        weights1[34186] <= 16'b1111111111110011;
        weights1[34187] <= 16'b1111111111111011;
        weights1[34188] <= 16'b1111111111111011;
        weights1[34189] <= 16'b0000000000001000;
        weights1[34190] <= 16'b0000000000010100;
        weights1[34191] <= 16'b1111111111111110;
        weights1[34192] <= 16'b0000000000001100;
        weights1[34193] <= 16'b1111111111101010;
        weights1[34194] <= 16'b1111111111111101;
        weights1[34195] <= 16'b0000000000000010;
        weights1[34196] <= 16'b1111111111111101;
        weights1[34197] <= 16'b1111111111111001;
        weights1[34198] <= 16'b0000000000010010;
        weights1[34199] <= 16'b1111111111110111;
        weights1[34200] <= 16'b0000000000000001;
        weights1[34201] <= 16'b1111111111110011;
        weights1[34202] <= 16'b0000000000001111;
        weights1[34203] <= 16'b1111111111111001;
        weights1[34204] <= 16'b0000000000000110;
        weights1[34205] <= 16'b1111111111111101;
        weights1[34206] <= 16'b0000000000001010;
        weights1[34207] <= 16'b1111111111111110;
        weights1[34208] <= 16'b0000000000000110;
        weights1[34209] <= 16'b0000000000001011;
        weights1[34210] <= 16'b0000000000000011;
        weights1[34211] <= 16'b0000000000000001;
        weights1[34212] <= 16'b0000000000011110;
        weights1[34213] <= 16'b1111111111111010;
        weights1[34214] <= 16'b1111111111111001;
        weights1[34215] <= 16'b1111111111110111;
        weights1[34216] <= 16'b1111111111111110;
        weights1[34217] <= 16'b0000000000001011;
        weights1[34218] <= 16'b0000000000000011;
        weights1[34219] <= 16'b0000000000000001;
        weights1[34220] <= 16'b1111111111111111;
        weights1[34221] <= 16'b1111111111111101;
        weights1[34222] <= 16'b0000000000010001;
        weights1[34223] <= 16'b1111111111111101;
        weights1[34224] <= 16'b0000000000010110;
        weights1[34225] <= 16'b0000000000000000;
        weights1[34226] <= 16'b0000000000000001;
        weights1[34227] <= 16'b0000000000000011;
        weights1[34228] <= 16'b0000000000001110;
        weights1[34229] <= 16'b0000000000001010;
        weights1[34230] <= 16'b0000000000010001;
        weights1[34231] <= 16'b1111111111111111;
        weights1[34232] <= 16'b1111111111111100;
        weights1[34233] <= 16'b0000000000000111;
        weights1[34234] <= 16'b0000000000000111;
        weights1[34235] <= 16'b1111111111111011;
        weights1[34236] <= 16'b1111111111111001;
        weights1[34237] <= 16'b0000000000000110;
        weights1[34238] <= 16'b0000000000000000;
        weights1[34239] <= 16'b0000000000000100;
        weights1[34240] <= 16'b0000000000000111;
        weights1[34241] <= 16'b0000000000001100;
        weights1[34242] <= 16'b0000000000001100;
        weights1[34243] <= 16'b1111111111111001;
        weights1[34244] <= 16'b0000000000000001;
        weights1[34245] <= 16'b1111111111111110;
        weights1[34246] <= 16'b0000000000000111;
        weights1[34247] <= 16'b0000000000011000;
        weights1[34248] <= 16'b0000000000001010;
        weights1[34249] <= 16'b1111111111111100;
        weights1[34250] <= 16'b1111111111111100;
        weights1[34251] <= 16'b1111111111111111;
        weights1[34252] <= 16'b0000000000000111;
        weights1[34253] <= 16'b1111111111110100;
        weights1[34254] <= 16'b0000000000000011;
        weights1[34255] <= 16'b0000000000000001;
        weights1[34256] <= 16'b1111111111110100;
        weights1[34257] <= 16'b1111111111111000;
        weights1[34258] <= 16'b0000000000010110;
        weights1[34259] <= 16'b0000000000001100;
        weights1[34260] <= 16'b0000000000000101;
        weights1[34261] <= 16'b1111111111111100;
        weights1[34262] <= 16'b1111111111111011;
        weights1[34263] <= 16'b1111111111111000;
        weights1[34264] <= 16'b0000000000000111;
        weights1[34265] <= 16'b0000000000000001;
        weights1[34266] <= 16'b0000000000001101;
        weights1[34267] <= 16'b0000000000000010;
        weights1[34268] <= 16'b1111111111101110;
        weights1[34269] <= 16'b1111111111111110;
        weights1[34270] <= 16'b0000000000001111;
        weights1[34271] <= 16'b1111111111110110;
        weights1[34272] <= 16'b0000000000000111;
        weights1[34273] <= 16'b0000000000000011;
        weights1[34274] <= 16'b0000000000001000;
        weights1[34275] <= 16'b1111111111111110;
        weights1[34276] <= 16'b1111111111110100;
        weights1[34277] <= 16'b1111111111111100;
        weights1[34278] <= 16'b1111111111111010;
        weights1[34279] <= 16'b0000000000001101;
        weights1[34280] <= 16'b1111111111110110;
        weights1[34281] <= 16'b0000000000000001;
        weights1[34282] <= 16'b1111111111111110;
        weights1[34283] <= 16'b1111111111110011;
        weights1[34284] <= 16'b1111111111101110;
        weights1[34285] <= 16'b0000000000000000;
        weights1[34286] <= 16'b0000000000000011;
        weights1[34287] <= 16'b0000000000001010;
        weights1[34288] <= 16'b1111111111111100;
        weights1[34289] <= 16'b1111111111111101;
        weights1[34290] <= 16'b0000000000000000;
        weights1[34291] <= 16'b0000000000010011;
        weights1[34292] <= 16'b1111111111110010;
        weights1[34293] <= 16'b1111111111111111;
        weights1[34294] <= 16'b1111111111111000;
        weights1[34295] <= 16'b0000000000000100;
        weights1[34296] <= 16'b1111111111111111;
        weights1[34297] <= 16'b1111111111111111;
        weights1[34298] <= 16'b0000000000000001;
        weights1[34299] <= 16'b1111111111111001;
        weights1[34300] <= 16'b0000000000000011;
        weights1[34301] <= 16'b1111111111111011;
        weights1[34302] <= 16'b1111111111111110;
        weights1[34303] <= 16'b0000000000000111;
        weights1[34304] <= 16'b0000000000000111;
        weights1[34305] <= 16'b0000000000000010;
        weights1[34306] <= 16'b0000000000001011;
        weights1[34307] <= 16'b1111111111110110;
        weights1[34308] <= 16'b0000000000001101;
        weights1[34309] <= 16'b1111111111111001;
        weights1[34310] <= 16'b1111111111110100;
        weights1[34311] <= 16'b0000000000000010;
        weights1[34312] <= 16'b1111111111101111;
        weights1[34313] <= 16'b0000000000000111;
        weights1[34314] <= 16'b1111111111111101;
        weights1[34315] <= 16'b0000000000000011;
        weights1[34316] <= 16'b0000000000011000;
        weights1[34317] <= 16'b0000000000000100;
        weights1[34318] <= 16'b1111111111111100;
        weights1[34319] <= 16'b1111111111111100;
        weights1[34320] <= 16'b0000000000000000;
        weights1[34321] <= 16'b0000000000000010;
        weights1[34322] <= 16'b1111111111111010;
        weights1[34323] <= 16'b1111111111111100;
        weights1[34324] <= 16'b1111111111111010;
        weights1[34325] <= 16'b1111111111110101;
        weights1[34326] <= 16'b1111111111111110;
        weights1[34327] <= 16'b1111111111101111;
        weights1[34328] <= 16'b0000000000000001;
        weights1[34329] <= 16'b0000000000000000;
        weights1[34330] <= 16'b0000000000000110;
        weights1[34331] <= 16'b1111111111111011;
        weights1[34332] <= 16'b1111111111101111;
        weights1[34333] <= 16'b0000000000010000;
        weights1[34334] <= 16'b0000000000010010;
        weights1[34335] <= 16'b1111111111111011;
        weights1[34336] <= 16'b1111111111111001;
        weights1[34337] <= 16'b1111111111111011;
        weights1[34338] <= 16'b0000000000000110;
        weights1[34339] <= 16'b1111111111110100;
        weights1[34340] <= 16'b1111111111110101;
        weights1[34341] <= 16'b1111111111111011;
        weights1[34342] <= 16'b1111111111100010;
        weights1[34343] <= 16'b1111111111110000;
        weights1[34344] <= 16'b1111111111111100;
        weights1[34345] <= 16'b1111111111110000;
        weights1[34346] <= 16'b0000000000001101;
        weights1[34347] <= 16'b1111111111111100;
        weights1[34348] <= 16'b0000000000010001;
        weights1[34349] <= 16'b0000000000001101;
        weights1[34350] <= 16'b1111111111111001;
        weights1[34351] <= 16'b1111111111110100;
        weights1[34352] <= 16'b1111111111111111;
        weights1[34353] <= 16'b1111111111101011;
        weights1[34354] <= 16'b1111111111110101;
        weights1[34355] <= 16'b1111111111110101;
        weights1[34356] <= 16'b0000000000000010;
        weights1[34357] <= 16'b0000000000000101;
        weights1[34358] <= 16'b0000000000000100;
        weights1[34359] <= 16'b1111111111111001;
        weights1[34360] <= 16'b1111111111101101;
        weights1[34361] <= 16'b1111111111110111;
        weights1[34362] <= 16'b1111111111110111;
        weights1[34363] <= 16'b1111111111111100;
        weights1[34364] <= 16'b1111111111111100;
        weights1[34365] <= 16'b0000000000001001;
        weights1[34366] <= 16'b1111111111101000;
        weights1[34367] <= 16'b0000000000000000;
        weights1[34368] <= 16'b1111111111101111;
        weights1[34369] <= 16'b1111111111111001;
        weights1[34370] <= 16'b0000000000001000;
        weights1[34371] <= 16'b1111111111100010;
        weights1[34372] <= 16'b0000000000010110;
        weights1[34373] <= 16'b0000000000001000;
        weights1[34374] <= 16'b1111111111111001;
        weights1[34375] <= 16'b1111111111111010;
        weights1[34376] <= 16'b0000000000001011;
        weights1[34377] <= 16'b1111111111101000;
        weights1[34378] <= 16'b0000000000001000;
        weights1[34379] <= 16'b0000000000001011;
        weights1[34380] <= 16'b1111111111101110;
        weights1[34381] <= 16'b1111111111110110;
        weights1[34382] <= 16'b1111111111111000;
        weights1[34383] <= 16'b1111111111110010;
        weights1[34384] <= 16'b0000000000000001;
        weights1[34385] <= 16'b0000000000000000;
        weights1[34386] <= 16'b1111111111111001;
        weights1[34387] <= 16'b1111111111101101;
        weights1[34388] <= 16'b1111111111111010;
        weights1[34389] <= 16'b0000000000000101;
        weights1[34390] <= 16'b0000000000000001;
        weights1[34391] <= 16'b0000000000000011;
        weights1[34392] <= 16'b1111111111110000;
        weights1[34393] <= 16'b0000000000001011;
        weights1[34394] <= 16'b0000000000000111;
        weights1[34395] <= 16'b1111111111110101;
        weights1[34396] <= 16'b1111111111111000;
        weights1[34397] <= 16'b0000000000010101;
        weights1[34398] <= 16'b0000000000010101;
        weights1[34399] <= 16'b1111111111101110;
        weights1[34400] <= 16'b1111111111101010;
        weights1[34401] <= 16'b1111111111100101;
        weights1[34402] <= 16'b1111111111101101;
        weights1[34403] <= 16'b0000000000000011;
        weights1[34404] <= 16'b1111111111100111;
        weights1[34405] <= 16'b1111111111101111;
        weights1[34406] <= 16'b1111111111111011;
        weights1[34407] <= 16'b0000000000000100;
        weights1[34408] <= 16'b1111111111110110;
        weights1[34409] <= 16'b1111111111111100;
        weights1[34410] <= 16'b1111111111110111;
        weights1[34411] <= 16'b1111111111111010;
        weights1[34412] <= 16'b1111111111111111;
        weights1[34413] <= 16'b1111111111111010;
        weights1[34414] <= 16'b1111111111111111;
        weights1[34415] <= 16'b1111111111111100;
        weights1[34416] <= 16'b0000000000000110;
        weights1[34417] <= 16'b1111111111111001;
        weights1[34418] <= 16'b1111111111111101;
        weights1[34419] <= 16'b1111111111111110;
        weights1[34420] <= 16'b0000000000000111;
        weights1[34421] <= 16'b1111111111111111;
        weights1[34422] <= 16'b1111111111111111;
        weights1[34423] <= 16'b1111111111111000;
        weights1[34424] <= 16'b1111111111100110;
        weights1[34425] <= 16'b1111111111101110;
        weights1[34426] <= 16'b1111111111111010;
        weights1[34427] <= 16'b1111111111110101;
        weights1[34428] <= 16'b1111111111110011;
        weights1[34429] <= 16'b1111111111111110;
        weights1[34430] <= 16'b1111111111101001;
        weights1[34431] <= 16'b1111111111101010;
        weights1[34432] <= 16'b1111111111101100;
        weights1[34433] <= 16'b1111111111101111;
        weights1[34434] <= 16'b1111111111100000;
        weights1[34435] <= 16'b1111111111110001;
        weights1[34436] <= 16'b1111111111110010;
        weights1[34437] <= 16'b1111111111110100;
        weights1[34438] <= 16'b1111111111111111;
        weights1[34439] <= 16'b0000000000000000;
        weights1[34440] <= 16'b0000000000000000;
        weights1[34441] <= 16'b1111111111111110;
        weights1[34442] <= 16'b0000000000000010;
        weights1[34443] <= 16'b1111111111111111;
        weights1[34444] <= 16'b1111111111111011;
        weights1[34445] <= 16'b1111111111110011;
        weights1[34446] <= 16'b1111111111110001;
        weights1[34447] <= 16'b1111111111111010;
        weights1[34448] <= 16'b0000000000000000;
        weights1[34449] <= 16'b0000000000000100;
        weights1[34450] <= 16'b1111111111111010;
        weights1[34451] <= 16'b1111111111110110;
        weights1[34452] <= 16'b0000000000000100;
        weights1[34453] <= 16'b1111111111100100;
        weights1[34454] <= 16'b1111111111111001;
        weights1[34455] <= 16'b1111111111100110;
        weights1[34456] <= 16'b1111111111111001;
        weights1[34457] <= 16'b1111111111101110;
        weights1[34458] <= 16'b1111111111111111;
        weights1[34459] <= 16'b1111111111101101;
        weights1[34460] <= 16'b0000000000000000;
        weights1[34461] <= 16'b1111111111111000;
        weights1[34462] <= 16'b1111111111101101;
        weights1[34463] <= 16'b1111111111111001;
        weights1[34464] <= 16'b1111111111101110;
        weights1[34465] <= 16'b1111111111111011;
        weights1[34466] <= 16'b1111111111111111;
        weights1[34467] <= 16'b0000000000000001;
        weights1[34468] <= 16'b0000000000000000;
        weights1[34469] <= 16'b0000000000000001;
        weights1[34470] <= 16'b0000000000000100;
        weights1[34471] <= 16'b0000000000001000;
        weights1[34472] <= 16'b0000000000000100;
        weights1[34473] <= 16'b1111111111110001;
        weights1[34474] <= 16'b1111111111100110;
        weights1[34475] <= 16'b1111111111110001;
        weights1[34476] <= 16'b1111111111111000;
        weights1[34477] <= 16'b0000000000000010;
        weights1[34478] <= 16'b1111111111111101;
        weights1[34479] <= 16'b1111111111110000;
        weights1[34480] <= 16'b0000000000000011;
        weights1[34481] <= 16'b1111111111111001;
        weights1[34482] <= 16'b1111111111100011;
        weights1[34483] <= 16'b1111111111110001;
        weights1[34484] <= 16'b1111111111101111;
        weights1[34485] <= 16'b1111111111101111;
        weights1[34486] <= 16'b1111111111101010;
        weights1[34487] <= 16'b1111111111100100;
        weights1[34488] <= 16'b1111111111111010;
        weights1[34489] <= 16'b1111111111110000;
        weights1[34490] <= 16'b1111111111110101;
        weights1[34491] <= 16'b1111111111110111;
        weights1[34492] <= 16'b1111111111110011;
        weights1[34493] <= 16'b1111111111111100;
        weights1[34494] <= 16'b0000000000000001;
        weights1[34495] <= 16'b0000000000000001;
        weights1[34496] <= 16'b1111111111111111;
        weights1[34497] <= 16'b1111111111111111;
        weights1[34498] <= 16'b1111111111111101;
        weights1[34499] <= 16'b1111111111111101;
        weights1[34500] <= 16'b1111111111111011;
        weights1[34501] <= 16'b1111111111110111;
        weights1[34502] <= 16'b1111111111111000;
        weights1[34503] <= 16'b1111111111111001;
        weights1[34504] <= 16'b1111111111101111;
        weights1[34505] <= 16'b1111111111101110;
        weights1[34506] <= 16'b1111111111100111;
        weights1[34507] <= 16'b1111111111010011;
        weights1[34508] <= 16'b1111111111001010;
        weights1[34509] <= 16'b1111111110111000;
        weights1[34510] <= 16'b1111111110110000;
        weights1[34511] <= 16'b1111111110101001;
        weights1[34512] <= 16'b1111111110010011;
        weights1[34513] <= 16'b1111111110100110;
        weights1[34514] <= 16'b1111111111000000;
        weights1[34515] <= 16'b1111111111001110;
        weights1[34516] <= 16'b1111111111011001;
        weights1[34517] <= 16'b1111111111100011;
        weights1[34518] <= 16'b1111111111110000;
        weights1[34519] <= 16'b1111111111111100;
        weights1[34520] <= 16'b1111111111111111;
        weights1[34521] <= 16'b0000000000000000;
        weights1[34522] <= 16'b0000000000000000;
        weights1[34523] <= 16'b0000000000000000;
        weights1[34524] <= 16'b1111111111111111;
        weights1[34525] <= 16'b0000000000000000;
        weights1[34526] <= 16'b1111111111111010;
        weights1[34527] <= 16'b1111111111111110;
        weights1[34528] <= 16'b1111111111111010;
        weights1[34529] <= 16'b1111111111110011;
        weights1[34530] <= 16'b1111111111111100;
        weights1[34531] <= 16'b1111111111111011;
        weights1[34532] <= 16'b0000000000010011;
        weights1[34533] <= 16'b1111111111111110;
        weights1[34534] <= 16'b0000000000000011;
        weights1[34535] <= 16'b0000000000000110;
        weights1[34536] <= 16'b1111111111110110;
        weights1[34537] <= 16'b1111111111100000;
        weights1[34538] <= 16'b1111111111011010;
        weights1[34539] <= 16'b1111111111001000;
        weights1[34540] <= 16'b1111111110101010;
        weights1[34541] <= 16'b1111111110010111;
        weights1[34542] <= 16'b1111111110101000;
        weights1[34543] <= 16'b1111111110111000;
        weights1[34544] <= 16'b1111111111001001;
        weights1[34545] <= 16'b1111111111011011;
        weights1[34546] <= 16'b1111111111101100;
        weights1[34547] <= 16'b1111111111110100;
        weights1[34548] <= 16'b1111111111111100;
        weights1[34549] <= 16'b1111111111111100;
        weights1[34550] <= 16'b1111111111111110;
        weights1[34551] <= 16'b1111111111111111;
        weights1[34552] <= 16'b1111111111111110;
        weights1[34553] <= 16'b1111111111111011;
        weights1[34554] <= 16'b1111111111111101;
        weights1[34555] <= 16'b0000000000000001;
        weights1[34556] <= 16'b1111111111111000;
        weights1[34557] <= 16'b1111111111111000;
        weights1[34558] <= 16'b1111111111111111;
        weights1[34559] <= 16'b0000000000000001;
        weights1[34560] <= 16'b0000000000010100;
        weights1[34561] <= 16'b0000000000100000;
        weights1[34562] <= 16'b0000000000100100;
        weights1[34563] <= 16'b0000000000010000;
        weights1[34564] <= 16'b0000000000110001;
        weights1[34565] <= 16'b0000000000101001;
        weights1[34566] <= 16'b1111111111111100;
        weights1[34567] <= 16'b1111111111101100;
        weights1[34568] <= 16'b1111111111100011;
        weights1[34569] <= 16'b1111111110111100;
        weights1[34570] <= 16'b1111111110010100;
        weights1[34571] <= 16'b1111111110011010;
        weights1[34572] <= 16'b1111111110101001;
        weights1[34573] <= 16'b1111111111000101;
        weights1[34574] <= 16'b1111111111010111;
        weights1[34575] <= 16'b1111111111101101;
        weights1[34576] <= 16'b1111111111110001;
        weights1[34577] <= 16'b1111111111110111;
        weights1[34578] <= 16'b1111111111111010;
        weights1[34579] <= 16'b1111111111111111;
        weights1[34580] <= 16'b1111111111111110;
        weights1[34581] <= 16'b1111111111111111;
        weights1[34582] <= 16'b0000000000000010;
        weights1[34583] <= 16'b1111111111111100;
        weights1[34584] <= 16'b0000000000000101;
        weights1[34585] <= 16'b1111111111110011;
        weights1[34586] <= 16'b0000000000000010;
        weights1[34587] <= 16'b1111111111111111;
        weights1[34588] <= 16'b0000000000010000;
        weights1[34589] <= 16'b0000000000001011;
        weights1[34590] <= 16'b0000000000010011;
        weights1[34591] <= 16'b0000000000110011;
        weights1[34592] <= 16'b0000000000100110;
        weights1[34593] <= 16'b0000000000101110;
        weights1[34594] <= 16'b0000000000101001;
        weights1[34595] <= 16'b0000000000010001;
        weights1[34596] <= 16'b1111111111110100;
        weights1[34597] <= 16'b1111111111111100;
        weights1[34598] <= 16'b1111111111001011;
        weights1[34599] <= 16'b1111111110011010;
        weights1[34600] <= 16'b1111111110000110;
        weights1[34601] <= 16'b1111111110001111;
        weights1[34602] <= 16'b1111111110111100;
        weights1[34603] <= 16'b1111111111011100;
        weights1[34604] <= 16'b1111111111101010;
        weights1[34605] <= 16'b1111111111101110;
        weights1[34606] <= 16'b1111111111111000;
        weights1[34607] <= 16'b1111111111111110;
        weights1[34608] <= 16'b1111111111111110;
        weights1[34609] <= 16'b0000000000000101;
        weights1[34610] <= 16'b0000000000000010;
        weights1[34611] <= 16'b1111111111111001;
        weights1[34612] <= 16'b0000000000000011;
        weights1[34613] <= 16'b0000000000000000;
        weights1[34614] <= 16'b0000000000010001;
        weights1[34615] <= 16'b0000000000010000;
        weights1[34616] <= 16'b0000000000000001;
        weights1[34617] <= 16'b0000000000101010;
        weights1[34618] <= 16'b0000000000011010;
        weights1[34619] <= 16'b0000000000110111;
        weights1[34620] <= 16'b0000000001000110;
        weights1[34621] <= 16'b0000000001000100;
        weights1[34622] <= 16'b0000000000101001;
        weights1[34623] <= 16'b0000000000011001;
        weights1[34624] <= 16'b0000000000001111;
        weights1[34625] <= 16'b1111111111111110;
        weights1[34626] <= 16'b1111111111101010;
        weights1[34627] <= 16'b1111111111011110;
        weights1[34628] <= 16'b1111111110110011;
        weights1[34629] <= 16'b1111111101110100;
        weights1[34630] <= 16'b1111111110011101;
        weights1[34631] <= 16'b1111111111001101;
        weights1[34632] <= 16'b1111111111100001;
        weights1[34633] <= 16'b1111111111101000;
        weights1[34634] <= 16'b1111111111111010;
        weights1[34635] <= 16'b1111111111111110;
        weights1[34636] <= 16'b1111111111111010;
        weights1[34637] <= 16'b1111111111111011;
        weights1[34638] <= 16'b1111111111111010;
        weights1[34639] <= 16'b1111111111110010;
        weights1[34640] <= 16'b1111111111111010;
        weights1[34641] <= 16'b0000000000000100;
        weights1[34642] <= 16'b0000000000001010;
        weights1[34643] <= 16'b0000000000001110;
        weights1[34644] <= 16'b0000000000010011;
        weights1[34645] <= 16'b0000000000001100;
        weights1[34646] <= 16'b0000000000011001;
        weights1[34647] <= 16'b0000000000011100;
        weights1[34648] <= 16'b0000000000100011;
        weights1[34649] <= 16'b0000000000110000;
        weights1[34650] <= 16'b1111111111111110;
        weights1[34651] <= 16'b0000000000101000;
        weights1[34652] <= 16'b0000000000001001;
        weights1[34653] <= 16'b1111111111110111;
        weights1[34654] <= 16'b0000000000000001;
        weights1[34655] <= 16'b1111111111111111;
        weights1[34656] <= 16'b1111111111100100;
        weights1[34657] <= 16'b1111111110101100;
        weights1[34658] <= 16'b1111111110010110;
        weights1[34659] <= 16'b1111111111000001;
        weights1[34660] <= 16'b1111111111010100;
        weights1[34661] <= 16'b1111111111101000;
        weights1[34662] <= 16'b1111111111110111;
        weights1[34663] <= 16'b1111111111111011;
        weights1[34664] <= 16'b1111111111110100;
        weights1[34665] <= 16'b1111111111110100;
        weights1[34666] <= 16'b1111111111110000;
        weights1[34667] <= 16'b1111111111101011;
        weights1[34668] <= 16'b1111111111011001;
        weights1[34669] <= 16'b1111111111110110;
        weights1[34670] <= 16'b1111111111111100;
        weights1[34671] <= 16'b1111111111101001;
        weights1[34672] <= 16'b1111111111111111;
        weights1[34673] <= 16'b1111111111110111;
        weights1[34674] <= 16'b1111111111110010;
        weights1[34675] <= 16'b0000000000000011;
        weights1[34676] <= 16'b1111111111111001;
        weights1[34677] <= 16'b0000000000101010;
        weights1[34678] <= 16'b0000000001001000;
        weights1[34679] <= 16'b0000000000010110;
        weights1[34680] <= 16'b0000000000100101;
        weights1[34681] <= 16'b0000000000010111;
        weights1[34682] <= 16'b0000000000010111;
        weights1[34683] <= 16'b1111111111110110;
        weights1[34684] <= 16'b1111111111100111;
        weights1[34685] <= 16'b1111111110111010;
        weights1[34686] <= 16'b1111111110010110;
        weights1[34687] <= 16'b1111111110010010;
        weights1[34688] <= 16'b1111111110111110;
        weights1[34689] <= 16'b1111111111011101;
        weights1[34690] <= 16'b1111111111110001;
        weights1[34691] <= 16'b1111111111111100;
        weights1[34692] <= 16'b1111111111110101;
        weights1[34693] <= 16'b1111111111110101;
        weights1[34694] <= 16'b1111111111100101;
        weights1[34695] <= 16'b1111111111010001;
        weights1[34696] <= 16'b1111111111010010;
        weights1[34697] <= 16'b1111111111001100;
        weights1[34698] <= 16'b1111111111110010;
        weights1[34699] <= 16'b1111111111010011;
        weights1[34700] <= 16'b1111111111011110;
        weights1[34701] <= 16'b1111111110111011;
        weights1[34702] <= 16'b1111111111101000;
        weights1[34703] <= 16'b1111111111110000;
        weights1[34704] <= 16'b1111111111110110;
        weights1[34705] <= 16'b0000000000110011;
        weights1[34706] <= 16'b0000000001011101;
        weights1[34707] <= 16'b0000000000110011;
        weights1[34708] <= 16'b0000000000100100;
        weights1[34709] <= 16'b0000000000100000;
        weights1[34710] <= 16'b0000000000000110;
        weights1[34711] <= 16'b0000000000000010;
        weights1[34712] <= 16'b1111111111111011;
        weights1[34713] <= 16'b1111111111110110;
        weights1[34714] <= 16'b1111111111001011;
        weights1[34715] <= 16'b1111111110001011;
        weights1[34716] <= 16'b1111111110110111;
        weights1[34717] <= 16'b1111111111011110;
        weights1[34718] <= 16'b1111111111101011;
        weights1[34719] <= 16'b1111111111111011;
        weights1[34720] <= 16'b1111111111111010;
        weights1[34721] <= 16'b1111111111101110;
        weights1[34722] <= 16'b1111111111011110;
        weights1[34723] <= 16'b1111111111100100;
        weights1[34724] <= 16'b1111111111001010;
        weights1[34725] <= 16'b1111111111001111;
        weights1[34726] <= 16'b1111111111011001;
        weights1[34727] <= 16'b1111111111000101;
        weights1[34728] <= 16'b1111111111001101;
        weights1[34729] <= 16'b1111111111110000;
        weights1[34730] <= 16'b1111111111110100;
        weights1[34731] <= 16'b1111111111100101;
        weights1[34732] <= 16'b1111111111101001;
        weights1[34733] <= 16'b1111111111111101;
        weights1[34734] <= 16'b0000000000101001;
        weights1[34735] <= 16'b0000000001010100;
        weights1[34736] <= 16'b0000000001001000;
        weights1[34737] <= 16'b0000000000100010;
        weights1[34738] <= 16'b0000000000100000;
        weights1[34739] <= 16'b0000000000001111;
        weights1[34740] <= 16'b0000000000000001;
        weights1[34741] <= 16'b1111111111111010;
        weights1[34742] <= 16'b1111111111011000;
        weights1[34743] <= 16'b1111111110010110;
        weights1[34744] <= 16'b1111111110101010;
        weights1[34745] <= 16'b1111111111001100;
        weights1[34746] <= 16'b1111111111101100;
        weights1[34747] <= 16'b1111111111110100;
        weights1[34748] <= 16'b1111111111111011;
        weights1[34749] <= 16'b1111111111101100;
        weights1[34750] <= 16'b1111111111010111;
        weights1[34751] <= 16'b1111111111100000;
        weights1[34752] <= 16'b1111111111011001;
        weights1[34753] <= 16'b1111111111001001;
        weights1[34754] <= 16'b1111111111100100;
        weights1[34755] <= 16'b1111111111101011;
        weights1[34756] <= 16'b1111111111110101;
        weights1[34757] <= 16'b1111111111101011;
        weights1[34758] <= 16'b1111111111111001;
        weights1[34759] <= 16'b1111111111100101;
        weights1[34760] <= 16'b1111111111011011;
        weights1[34761] <= 16'b1111111111101111;
        weights1[34762] <= 16'b0000000000001011;
        weights1[34763] <= 16'b0000000000110001;
        weights1[34764] <= 16'b0000000001000101;
        weights1[34765] <= 16'b0000000000100000;
        weights1[34766] <= 16'b0000000000100010;
        weights1[34767] <= 16'b0000000000010001;
        weights1[34768] <= 16'b0000000000000101;
        weights1[34769] <= 16'b0000000000000101;
        weights1[34770] <= 16'b1111111111001111;
        weights1[34771] <= 16'b1111111110101110;
        weights1[34772] <= 16'b1111111110111001;
        weights1[34773] <= 16'b1111111111011010;
        weights1[34774] <= 16'b1111111111101110;
        weights1[34775] <= 16'b1111111111110101;
        weights1[34776] <= 16'b1111111111111101;
        weights1[34777] <= 16'b1111111111101110;
        weights1[34778] <= 16'b1111111111100000;
        weights1[34779] <= 16'b1111111111101011;
        weights1[34780] <= 16'b1111111111110100;
        weights1[34781] <= 16'b0000000000000000;
        weights1[34782] <= 16'b0000000000001100;
        weights1[34783] <= 16'b1111111111110010;
        weights1[34784] <= 16'b0000000000000100;
        weights1[34785] <= 16'b1111111111101100;
        weights1[34786] <= 16'b1111111111110100;
        weights1[34787] <= 16'b1111111111110101;
        weights1[34788] <= 16'b1111111111110110;
        weights1[34789] <= 16'b1111111111001111;
        weights1[34790] <= 16'b1111111111110101;
        weights1[34791] <= 16'b0000000000010100;
        weights1[34792] <= 16'b0000000000110111;
        weights1[34793] <= 16'b0000000000110110;
        weights1[34794] <= 16'b0000000000100010;
        weights1[34795] <= 16'b0000000000101000;
        weights1[34796] <= 16'b1111111111110011;
        weights1[34797] <= 16'b0000000000000011;
        weights1[34798] <= 16'b1111111111110100;
        weights1[34799] <= 16'b1111111110100100;
        weights1[34800] <= 16'b1111111110110110;
        weights1[34801] <= 16'b1111111111011010;
        weights1[34802] <= 16'b1111111111100101;
        weights1[34803] <= 16'b1111111111110110;
        weights1[34804] <= 16'b1111111111111100;
        weights1[34805] <= 16'b1111111111110111;
        weights1[34806] <= 16'b1111111111101101;
        weights1[34807] <= 16'b0000000000000100;
        weights1[34808] <= 16'b1111111111111110;
        weights1[34809] <= 16'b0000000000011010;
        weights1[34810] <= 16'b0000000000010000;
        weights1[34811] <= 16'b0000000000010111;
        weights1[34812] <= 16'b1111111111111111;
        weights1[34813] <= 16'b0000000000001010;
        weights1[34814] <= 16'b1111111111110111;
        weights1[34815] <= 16'b1111111111110010;
        weights1[34816] <= 16'b1111111111001011;
        weights1[34817] <= 16'b1111111111101111;
        weights1[34818] <= 16'b1111111111100111;
        weights1[34819] <= 16'b0000000000011100;
        weights1[34820] <= 16'b0000000000000111;
        weights1[34821] <= 16'b0000000000101111;
        weights1[34822] <= 16'b0000000000100010;
        weights1[34823] <= 16'b0000000000101100;
        weights1[34824] <= 16'b0000000000101100;
        weights1[34825] <= 16'b0000000000000111;
        weights1[34826] <= 16'b1111111111011101;
        weights1[34827] <= 16'b1111111111001001;
        weights1[34828] <= 16'b1111111110101011;
        weights1[34829] <= 16'b1111111111100010;
        weights1[34830] <= 16'b1111111111110101;
        weights1[34831] <= 16'b1111111111111000;
        weights1[34832] <= 16'b0000000000001001;
        weights1[34833] <= 16'b0000000000000000;
        weights1[34834] <= 16'b1111111111111010;
        weights1[34835] <= 16'b0000000000000110;
        weights1[34836] <= 16'b0000000000000111;
        weights1[34837] <= 16'b1111111111110111;
        weights1[34838] <= 16'b0000000000001100;
        weights1[34839] <= 16'b1111111111111000;
        weights1[34840] <= 16'b1111111111111011;
        weights1[34841] <= 16'b1111111111111101;
        weights1[34842] <= 16'b1111111111101000;
        weights1[34843] <= 16'b1111111111011101;
        weights1[34844] <= 16'b1111111111010111;
        weights1[34845] <= 16'b1111111111011111;
        weights1[34846] <= 16'b1111111111110001;
        weights1[34847] <= 16'b0000000000000111;
        weights1[34848] <= 16'b1111111111111111;
        weights1[34849] <= 16'b0000000000011110;
        weights1[34850] <= 16'b0000000000001101;
        weights1[34851] <= 16'b0000000000010011;
        weights1[34852] <= 16'b0000000000011110;
        weights1[34853] <= 16'b0000000000010010;
        weights1[34854] <= 16'b1111111111100110;
        weights1[34855] <= 16'b1111111110111110;
        weights1[34856] <= 16'b1111111111010111;
        weights1[34857] <= 16'b1111111111101101;
        weights1[34858] <= 16'b1111111111111110;
        weights1[34859] <= 16'b0000000000000100;
        weights1[34860] <= 16'b0000000000010101;
        weights1[34861] <= 16'b0000000000000110;
        weights1[34862] <= 16'b1111111111111011;
        weights1[34863] <= 16'b0000000000000000;
        weights1[34864] <= 16'b1111111111110111;
        weights1[34865] <= 16'b1111111111110001;
        weights1[34866] <= 16'b0000000000000011;
        weights1[34867] <= 16'b1111111111101001;
        weights1[34868] <= 16'b1111111111111001;
        weights1[34869] <= 16'b1111111111110001;
        weights1[34870] <= 16'b1111111111100011;
        weights1[34871] <= 16'b1111111111110001;
        weights1[34872] <= 16'b1111111111101111;
        weights1[34873] <= 16'b1111111111010011;
        weights1[34874] <= 16'b1111111111101011;
        weights1[34875] <= 16'b1111111111110111;
        weights1[34876] <= 16'b0000000000010110;
        weights1[34877] <= 16'b0000000000011000;
        weights1[34878] <= 16'b0000000000001111;
        weights1[34879] <= 16'b0000000000010111;
        weights1[34880] <= 16'b0000000000000010;
        weights1[34881] <= 16'b1111111111111011;
        weights1[34882] <= 16'b1111111111111010;
        weights1[34883] <= 16'b1111111111011110;
        weights1[34884] <= 16'b1111111111100000;
        weights1[34885] <= 16'b1111111111110001;
        weights1[34886] <= 16'b1111111111111000;
        weights1[34887] <= 16'b1111111111111100;
        weights1[34888] <= 16'b0000000000010000;
        weights1[34889] <= 16'b0000000000001111;
        weights1[34890] <= 16'b1111111111111111;
        weights1[34891] <= 16'b0000000000001010;
        weights1[34892] <= 16'b0000000000001000;
        weights1[34893] <= 16'b1111111111111011;
        weights1[34894] <= 16'b1111111111011110;
        weights1[34895] <= 16'b1111111111111010;
        weights1[34896] <= 16'b1111111111111000;
        weights1[34897] <= 16'b1111111111110111;
        weights1[34898] <= 16'b1111111111101100;
        weights1[34899] <= 16'b1111111111111101;
        weights1[34900] <= 16'b1111111111110001;
        weights1[34901] <= 16'b1111111111110100;
        weights1[34902] <= 16'b1111111111101111;
        weights1[34903] <= 16'b0000000000000001;
        weights1[34904] <= 16'b0000000000000010;
        weights1[34905] <= 16'b0000000000011111;
        weights1[34906] <= 16'b0000000000010100;
        weights1[34907] <= 16'b0000000000001010;
        weights1[34908] <= 16'b1111111111111001;
        weights1[34909] <= 16'b1111111111110010;
        weights1[34910] <= 16'b1111111111110111;
        weights1[34911] <= 16'b1111111111110010;
        weights1[34912] <= 16'b1111111111111101;
        weights1[34913] <= 16'b1111111111101011;
        weights1[34914] <= 16'b0000000000001010;
        weights1[34915] <= 16'b1111111111111101;
        weights1[34916] <= 16'b0000000000001011;
        weights1[34917] <= 16'b0000000000001111;
        weights1[34918] <= 16'b0000000000001010;
        weights1[34919] <= 16'b1111111111111101;
        weights1[34920] <= 16'b1111111111110110;
        weights1[34921] <= 16'b1111111111111111;
        weights1[34922] <= 16'b1111111111111011;
        weights1[34923] <= 16'b1111111111111001;
        weights1[34924] <= 16'b1111111111111100;
        weights1[34925] <= 16'b1111111111111100;
        weights1[34926] <= 16'b1111111111110100;
        weights1[34927] <= 16'b0000000000001011;
        weights1[34928] <= 16'b1111111111110110;
        weights1[34929] <= 16'b1111111111111100;
        weights1[34930] <= 16'b1111111111111001;
        weights1[34931] <= 16'b0000000000000001;
        weights1[34932] <= 16'b0000000000000011;
        weights1[34933] <= 16'b0000000000010100;
        weights1[34934] <= 16'b1111111111111111;
        weights1[34935] <= 16'b1111111111111010;
        weights1[34936] <= 16'b0000000000000101;
        weights1[34937] <= 16'b1111111111011101;
        weights1[34938] <= 16'b1111111111100110;
        weights1[34939] <= 16'b1111111111111001;
        weights1[34940] <= 16'b1111111111101001;
        weights1[34941] <= 16'b0000000000000101;
        weights1[34942] <= 16'b0000000000000111;
        weights1[34943] <= 16'b0000000000000001;
        weights1[34944] <= 16'b0000000000001110;
        weights1[34945] <= 16'b0000000000011000;
        weights1[34946] <= 16'b0000000000010001;
        weights1[34947] <= 16'b0000000000001001;
        weights1[34948] <= 16'b0000000000000010;
        weights1[34949] <= 16'b0000000000001011;
        weights1[34950] <= 16'b1111111111110011;
        weights1[34951] <= 16'b0000000000000011;
        weights1[34952] <= 16'b1111111111110001;
        weights1[34953] <= 16'b1111111111110010;
        weights1[34954] <= 16'b0000000000000011;
        weights1[34955] <= 16'b1111111111110011;
        weights1[34956] <= 16'b1111111111101110;
        weights1[34957] <= 16'b1111111111011010;
        weights1[34958] <= 16'b1111111111011111;
        weights1[34959] <= 16'b1111111111100101;
        weights1[34960] <= 16'b1111111111111011;
        weights1[34961] <= 16'b0000000000000110;
        weights1[34962] <= 16'b0000000000000000;
        weights1[34963] <= 16'b1111111111110110;
        weights1[34964] <= 16'b1111111111111100;
        weights1[34965] <= 16'b0000000000001100;
        weights1[34966] <= 16'b1111111111110110;
        weights1[34967] <= 16'b1111111111100010;
        weights1[34968] <= 16'b0000000000000000;
        weights1[34969] <= 16'b1111111111111110;
        weights1[34970] <= 16'b1111111111111111;
        weights1[34971] <= 16'b0000000000001010;
        weights1[34972] <= 16'b0000000000001111;
        weights1[34973] <= 16'b0000000000010100;
        weights1[34974] <= 16'b0000000000011100;
        weights1[34975] <= 16'b0000000000001111;
        weights1[34976] <= 16'b0000000000000110;
        weights1[34977] <= 16'b1111111111111110;
        weights1[34978] <= 16'b1111111111111110;
        weights1[34979] <= 16'b1111111111110100;
        weights1[34980] <= 16'b0000000000000001;
        weights1[34981] <= 16'b1111111111100001;
        weights1[34982] <= 16'b1111111111110111;
        weights1[34983] <= 16'b1111111111100010;
        weights1[34984] <= 16'b0000000000000010;
        weights1[34985] <= 16'b1111111111111100;
        weights1[34986] <= 16'b1111111111111100;
        weights1[34987] <= 16'b0000000000000100;
        weights1[34988] <= 16'b1111111111110111;
        weights1[34989] <= 16'b1111111111111110;
        weights1[34990] <= 16'b1111111111110011;
        weights1[34991] <= 16'b1111111111110010;
        weights1[34992] <= 16'b1111111111110111;
        weights1[34993] <= 16'b1111111111110100;
        weights1[34994] <= 16'b1111111111110001;
        weights1[34995] <= 16'b1111111111011100;
        weights1[34996] <= 16'b1111111111110101;
        weights1[34997] <= 16'b0000000000000000;
        weights1[34998] <= 16'b1111111111111101;
        weights1[34999] <= 16'b0000000000001100;
        weights1[35000] <= 16'b0000000000001110;
        weights1[35001] <= 16'b0000000000011010;
        weights1[35002] <= 16'b0000000000001001;
        weights1[35003] <= 16'b0000000000001000;
        weights1[35004] <= 16'b0000000000000100;
        weights1[35005] <= 16'b0000000000011100;
        weights1[35006] <= 16'b0000000000001011;
        weights1[35007] <= 16'b0000000000001100;
        weights1[35008] <= 16'b0000000000000000;
        weights1[35009] <= 16'b0000000000001110;
        weights1[35010] <= 16'b0000000000000101;
        weights1[35011] <= 16'b0000000000001011;
        weights1[35012] <= 16'b1111111111110100;
        weights1[35013] <= 16'b1111111111111000;
        weights1[35014] <= 16'b1111111111101000;
        weights1[35015] <= 16'b1111111111100000;
        weights1[35016] <= 16'b0000000000001001;
        weights1[35017] <= 16'b1111111111111111;
        weights1[35018] <= 16'b0000000000010010;
        weights1[35019] <= 16'b0000000000001011;
        weights1[35020] <= 16'b1111111111110111;
        weights1[35021] <= 16'b0000000000001001;
        weights1[35022] <= 16'b1111111111111000;
        weights1[35023] <= 16'b1111111111110110;
        weights1[35024] <= 16'b0000000000100010;
        weights1[35025] <= 16'b0000000000010100;
        weights1[35026] <= 16'b0000000000000110;
        weights1[35027] <= 16'b0000000000001001;
        weights1[35028] <= 16'b0000000000001100;
        weights1[35029] <= 16'b0000000000001110;
        weights1[35030] <= 16'b0000000000010000;
        weights1[35031] <= 16'b0000000000001110;
        weights1[35032] <= 16'b1111111111111010;
        weights1[35033] <= 16'b0000000000011001;
        weights1[35034] <= 16'b0000000000000011;
        weights1[35035] <= 16'b1111111111111111;
        weights1[35036] <= 16'b0000000000010000;
        weights1[35037] <= 16'b1111111111111000;
        weights1[35038] <= 16'b1111111111111001;
        weights1[35039] <= 16'b1111111111111000;
        weights1[35040] <= 16'b0000000000001110;
        weights1[35041] <= 16'b1111111111110100;
        weights1[35042] <= 16'b1111111111111100;
        weights1[35043] <= 16'b1111111111101011;
        weights1[35044] <= 16'b1111111111110101;
        weights1[35045] <= 16'b0000000000001111;
        weights1[35046] <= 16'b0000000000000010;
        weights1[35047] <= 16'b1111111111111010;
        weights1[35048] <= 16'b0000000000001101;
        weights1[35049] <= 16'b0000000000001010;
        weights1[35050] <= 16'b1111111111111011;
        weights1[35051] <= 16'b0000000000000110;
        weights1[35052] <= 16'b1111111111111100;
        weights1[35053] <= 16'b1111111111111110;
        weights1[35054] <= 16'b0000000000000110;
        weights1[35055] <= 16'b0000000000000100;
        weights1[35056] <= 16'b0000000000010010;
        weights1[35057] <= 16'b0000000000011011;
        weights1[35058] <= 16'b0000000000001001;
        weights1[35059] <= 16'b0000000000000001;
        weights1[35060] <= 16'b0000000000010111;
        weights1[35061] <= 16'b1111111111110011;
        weights1[35062] <= 16'b0000000000000000;
        weights1[35063] <= 16'b0000000000010111;
        weights1[35064] <= 16'b0000000000000000;
        weights1[35065] <= 16'b1111111111101100;
        weights1[35066] <= 16'b1111111111110111;
        weights1[35067] <= 16'b0000000000000001;
        weights1[35068] <= 16'b0000000000000000;
        weights1[35069] <= 16'b0000000000001000;
        weights1[35070] <= 16'b0000000000010000;
        weights1[35071] <= 16'b1111111111111001;
        weights1[35072] <= 16'b1111111111111000;
        weights1[35073] <= 16'b1111111111110110;
        weights1[35074] <= 16'b1111111111111110;
        weights1[35075] <= 16'b0000000000010011;
        weights1[35076] <= 16'b1111111111111011;
        weights1[35077] <= 16'b1111111111110101;
        weights1[35078] <= 16'b1111111111111100;
        weights1[35079] <= 16'b0000000000010011;
        weights1[35080] <= 16'b0000000000010111;
        weights1[35081] <= 16'b0000000000000001;
        weights1[35082] <= 16'b1111111111111000;
        weights1[35083] <= 16'b1111111111111110;
        weights1[35084] <= 16'b0000000000100000;
        weights1[35085] <= 16'b0000000000010011;
        weights1[35086] <= 16'b0000000000010100;
        weights1[35087] <= 16'b1111111111111110;
        weights1[35088] <= 16'b0000000000001100;
        weights1[35089] <= 16'b1111111111110111;
        weights1[35090] <= 16'b0000000000000111;
        weights1[35091] <= 16'b0000000000010001;
        weights1[35092] <= 16'b0000000000001100;
        weights1[35093] <= 16'b0000000000000000;
        weights1[35094] <= 16'b0000000000011001;
        weights1[35095] <= 16'b1111111111111101;
        weights1[35096] <= 16'b1111111111110000;
        weights1[35097] <= 16'b1111111111110101;
        weights1[35098] <= 16'b1111111111111010;
        weights1[35099] <= 16'b1111111111110000;
        weights1[35100] <= 16'b1111111111100101;
        weights1[35101] <= 16'b1111111111110010;
        weights1[35102] <= 16'b1111111111100110;
        weights1[35103] <= 16'b1111111111111111;
        weights1[35104] <= 16'b0000000000000010;
        weights1[35105] <= 16'b1111111111111001;
        weights1[35106] <= 16'b0000000000000011;
        weights1[35107] <= 16'b1111111111111000;
        weights1[35108] <= 16'b1111111111111110;
        weights1[35109] <= 16'b1111111111110011;
        weights1[35110] <= 16'b1111111111110110;
        weights1[35111] <= 16'b0000000000000101;
        weights1[35112] <= 16'b0000000000001110;
        weights1[35113] <= 16'b0000000000010000;
        weights1[35114] <= 16'b0000000000000010;
        weights1[35115] <= 16'b0000000000001000;
        weights1[35116] <= 16'b0000000000000001;
        weights1[35117] <= 16'b0000000000011110;
        weights1[35118] <= 16'b0000000000010100;
        weights1[35119] <= 16'b0000000000000010;
        weights1[35120] <= 16'b0000000000000001;
        weights1[35121] <= 16'b1111111111111010;
        weights1[35122] <= 16'b0000000000001111;
        weights1[35123] <= 16'b1111111111110101;
        weights1[35124] <= 16'b0000000000000110;
        weights1[35125] <= 16'b1111111111101101;
        weights1[35126] <= 16'b0000000000001110;
        weights1[35127] <= 16'b0000000000000111;
        weights1[35128] <= 16'b1111111111111000;
        weights1[35129] <= 16'b0000000000000111;
        weights1[35130] <= 16'b1111111111110111;
        weights1[35131] <= 16'b0000000000000000;
        weights1[35132] <= 16'b1111111111100011;
        weights1[35133] <= 16'b0000000000010010;
        weights1[35134] <= 16'b0000000000001111;
        weights1[35135] <= 16'b1111111111110110;
        weights1[35136] <= 16'b0000000000000000;
        weights1[35137] <= 16'b1111111111111111;
        weights1[35138] <= 16'b1111111111111101;
        weights1[35139] <= 16'b0000000000000011;
        weights1[35140] <= 16'b0000000000010011;
        weights1[35141] <= 16'b0000000000001100;
        weights1[35142] <= 16'b0000000000001100;
        weights1[35143] <= 16'b1111111111111011;
        weights1[35144] <= 16'b1111111111110101;
        weights1[35145] <= 16'b1111111111101010;
        weights1[35146] <= 16'b0000000000001101;
        weights1[35147] <= 16'b0000000000100101;
        weights1[35148] <= 16'b0000000000000111;
        weights1[35149] <= 16'b1111111111101100;
        weights1[35150] <= 16'b0000000000010100;
        weights1[35151] <= 16'b1111111111110101;
        weights1[35152] <= 16'b0000000000010000;
        weights1[35153] <= 16'b1111111111111110;
        weights1[35154] <= 16'b1111111111101000;
        weights1[35155] <= 16'b1111111111101011;
        weights1[35156] <= 16'b1111111111101101;
        weights1[35157] <= 16'b1111111111100100;
        weights1[35158] <= 16'b1111111111111000;
        weights1[35159] <= 16'b1111111111110010;
        weights1[35160] <= 16'b1111111111101100;
        weights1[35161] <= 16'b0000000000001010;
        weights1[35162] <= 16'b0000000000000110;
        weights1[35163] <= 16'b1111111111111101;
        weights1[35164] <= 16'b1111111111101011;
        weights1[35165] <= 16'b0000000000000011;
        weights1[35166] <= 16'b0000000000000100;
        weights1[35167] <= 16'b0000000000000110;
        weights1[35168] <= 16'b0000000000010010;
        weights1[35169] <= 16'b0000000000001110;
        weights1[35170] <= 16'b0000000000001011;
        weights1[35171] <= 16'b0000000000000001;
        weights1[35172] <= 16'b0000000000010011;
        weights1[35173] <= 16'b0000000000010110;
        weights1[35174] <= 16'b0000000000000011;
        weights1[35175] <= 16'b0000000000010001;
        weights1[35176] <= 16'b1111111111101001;
        weights1[35177] <= 16'b1111111111111011;
        weights1[35178] <= 16'b0000000000010010;
        weights1[35179] <= 16'b1111111111110110;
        weights1[35180] <= 16'b1111111111101110;
        weights1[35181] <= 16'b0000000000001101;
        weights1[35182] <= 16'b1111111111100111;
        weights1[35183] <= 16'b1111111111111100;
        weights1[35184] <= 16'b0000000000000111;
        weights1[35185] <= 16'b0000000000001111;
        weights1[35186] <= 16'b1111111111100110;
        weights1[35187] <= 16'b1111111111101110;
        weights1[35188] <= 16'b1111111111110111;
        weights1[35189] <= 16'b1111111111111111;
        weights1[35190] <= 16'b1111111111110001;
        weights1[35191] <= 16'b1111111111110111;
        weights1[35192] <= 16'b1111111111111001;
        weights1[35193] <= 16'b0000000000000111;
        weights1[35194] <= 16'b0000000000000011;
        weights1[35195] <= 16'b0000000000000011;
        weights1[35196] <= 16'b0000000000001010;
        weights1[35197] <= 16'b0000000000010101;
        weights1[35198] <= 16'b0000000000011001;
        weights1[35199] <= 16'b0000000000001000;
        weights1[35200] <= 16'b0000000000001010;
        weights1[35201] <= 16'b0000000000010001;
        weights1[35202] <= 16'b0000000000000100;
        weights1[35203] <= 16'b1111111111111101;
        weights1[35204] <= 16'b0000000000000010;
        weights1[35205] <= 16'b0000000000011001;
        weights1[35206] <= 16'b0000000000001110;
        weights1[35207] <= 16'b0000000000010111;
        weights1[35208] <= 16'b0000000000010101;
        weights1[35209] <= 16'b0000000000011010;
        weights1[35210] <= 16'b0000000000000011;
        weights1[35211] <= 16'b0000000000000000;
        weights1[35212] <= 16'b1111111111111110;
        weights1[35213] <= 16'b0000000000001110;
        weights1[35214] <= 16'b0000000000001010;
        weights1[35215] <= 16'b1111111111110100;
        weights1[35216] <= 16'b1111111111110010;
        weights1[35217] <= 16'b0000000000000111;
        weights1[35218] <= 16'b0000000000001010;
        weights1[35219] <= 16'b1111111111111000;
        weights1[35220] <= 16'b1111111111111101;
        weights1[35221] <= 16'b1111111111110111;
        weights1[35222] <= 16'b1111111111111111;
        weights1[35223] <= 16'b0000000000000001;
        weights1[35224] <= 16'b0000000000000101;
        weights1[35225] <= 16'b0000000000010010;
        weights1[35226] <= 16'b0000000000011000;
        weights1[35227] <= 16'b0000000000011001;
        weights1[35228] <= 16'b0000000000010101;
        weights1[35229] <= 16'b1111111111111000;
        weights1[35230] <= 16'b1111111111111100;
        weights1[35231] <= 16'b0000000000000110;
        weights1[35232] <= 16'b0000000000001010;
        weights1[35233] <= 16'b1111111111111001;
        weights1[35234] <= 16'b0000000000010110;
        weights1[35235] <= 16'b1111111111100111;
        weights1[35236] <= 16'b1111111111110011;
        weights1[35237] <= 16'b1111111111111101;
        weights1[35238] <= 16'b0000000000001111;
        weights1[35239] <= 16'b1111111111100010;
        weights1[35240] <= 16'b1111111111111101;
        weights1[35241] <= 16'b0000000000001001;
        weights1[35242] <= 16'b0000000000001001;
        weights1[35243] <= 16'b1111111111101111;
        weights1[35244] <= 16'b1111111111111001;
        weights1[35245] <= 16'b0000000000000101;
        weights1[35246] <= 16'b0000000000000110;
        weights1[35247] <= 16'b0000000000000010;
        weights1[35248] <= 16'b0000000000000000;
        weights1[35249] <= 16'b1111111111111011;
        weights1[35250] <= 16'b0000000000000000;
        weights1[35251] <= 16'b0000000000000010;
        weights1[35252] <= 16'b0000000000000001;
        weights1[35253] <= 16'b0000000000001011;
        weights1[35254] <= 16'b0000000000001010;
        weights1[35255] <= 16'b0000000000001111;
        weights1[35256] <= 16'b0000000000000011;
        weights1[35257] <= 16'b1111111111111001;
        weights1[35258] <= 16'b0000000000000101;
        weights1[35259] <= 16'b0000000000000111;
        weights1[35260] <= 16'b0000000000000110;
        weights1[35261] <= 16'b0000000000000100;
        weights1[35262] <= 16'b0000000000001111;
        weights1[35263] <= 16'b0000000000000010;
        weights1[35264] <= 16'b0000000000001111;
        weights1[35265] <= 16'b0000000000001000;
        weights1[35266] <= 16'b0000000000001001;
        weights1[35267] <= 16'b0000000000001111;
        weights1[35268] <= 16'b0000000000000011;
        weights1[35269] <= 16'b0000000000000000;
        weights1[35270] <= 16'b1111111111110101;
        weights1[35271] <= 16'b1111111111111101;
        weights1[35272] <= 16'b0000000000000000;
        weights1[35273] <= 16'b0000000000000000;
        weights1[35274] <= 16'b1111111111110100;
        weights1[35275] <= 16'b0000000000000000;
        weights1[35276] <= 16'b0000000000000001;
        weights1[35277] <= 16'b0000000000000000;
        weights1[35278] <= 16'b0000000000000011;
        weights1[35279] <= 16'b0000000000000010;
        weights1[35280] <= 16'b0000000000000000;
        weights1[35281] <= 16'b0000000000000000;
        weights1[35282] <= 16'b0000000000000000;
        weights1[35283] <= 16'b1111111111111111;
        weights1[35284] <= 16'b1111111111111111;
        weights1[35285] <= 16'b1111111111111001;
        weights1[35286] <= 16'b1111111111110101;
        weights1[35287] <= 16'b1111111111110100;
        weights1[35288] <= 16'b1111111111101110;
        weights1[35289] <= 16'b1111111111011101;
        weights1[35290] <= 16'b1111111111001011;
        weights1[35291] <= 16'b1111111111001010;
        weights1[35292] <= 16'b1111111111010000;
        weights1[35293] <= 16'b1111111111110010;
        weights1[35294] <= 16'b0000000000010001;
        weights1[35295] <= 16'b0000000000011001;
        weights1[35296] <= 16'b0000000000100111;
        weights1[35297] <= 16'b0000000000110000;
        weights1[35298] <= 16'b0000000000011110;
        weights1[35299] <= 16'b0000000000011110;
        weights1[35300] <= 16'b0000000000100001;
        weights1[35301] <= 16'b0000000000001001;
        weights1[35302] <= 16'b1111111111111111;
        weights1[35303] <= 16'b1111111111111101;
        weights1[35304] <= 16'b0000000000000001;
        weights1[35305] <= 16'b1111111111111110;
        weights1[35306] <= 16'b1111111111111101;
        weights1[35307] <= 16'b1111111111111100;
        weights1[35308] <= 16'b0000000000000000;
        weights1[35309] <= 16'b0000000000000000;
        weights1[35310] <= 16'b0000000000000000;
        weights1[35311] <= 16'b0000000000000001;
        weights1[35312] <= 16'b1111111111111011;
        weights1[35313] <= 16'b1111111111110101;
        weights1[35314] <= 16'b1111111111110100;
        weights1[35315] <= 16'b1111111111101000;
        weights1[35316] <= 16'b1111111111100000;
        weights1[35317] <= 16'b1111111111010101;
        weights1[35318] <= 16'b1111111111000111;
        weights1[35319] <= 16'b1111111110111111;
        weights1[35320] <= 16'b1111111111100101;
        weights1[35321] <= 16'b1111111111101100;
        weights1[35322] <= 16'b0000000000000110;
        weights1[35323] <= 16'b0000000000011010;
        weights1[35324] <= 16'b0000000000100101;
        weights1[35325] <= 16'b0000000000011011;
        weights1[35326] <= 16'b0000000000011101;
        weights1[35327] <= 16'b0000000000010010;
        weights1[35328] <= 16'b0000000000001110;
        weights1[35329] <= 16'b0000000000000111;
        weights1[35330] <= 16'b0000000000001001;
        weights1[35331] <= 16'b0000000000000100;
        weights1[35332] <= 16'b0000000000000000;
        weights1[35333] <= 16'b1111111111110110;
        weights1[35334] <= 16'b1111111111110110;
        weights1[35335] <= 16'b1111111111111100;
        weights1[35336] <= 16'b0000000000000000;
        weights1[35337] <= 16'b0000000000000000;
        weights1[35338] <= 16'b1111111111111110;
        weights1[35339] <= 16'b1111111111111111;
        weights1[35340] <= 16'b1111111111111011;
        weights1[35341] <= 16'b1111111111111000;
        weights1[35342] <= 16'b1111111111101010;
        weights1[35343] <= 16'b1111111111100001;
        weights1[35344] <= 16'b1111111111010001;
        weights1[35345] <= 16'b1111111111010011;
        weights1[35346] <= 16'b1111111111000000;
        weights1[35347] <= 16'b1111111111011101;
        weights1[35348] <= 16'b0000000000010001;
        weights1[35349] <= 16'b0000000000010110;
        weights1[35350] <= 16'b0000000000010110;
        weights1[35351] <= 16'b0000000000100000;
        weights1[35352] <= 16'b0000000000010111;
        weights1[35353] <= 16'b0000000000011010;
        weights1[35354] <= 16'b0000000000001011;
        weights1[35355] <= 16'b0000000000011100;
        weights1[35356] <= 16'b0000000000001111;
        weights1[35357] <= 16'b1111111111111101;
        weights1[35358] <= 16'b1111111111111000;
        weights1[35359] <= 16'b1111111111101111;
        weights1[35360] <= 16'b1111111111101011;
        weights1[35361] <= 16'b1111111111101111;
        weights1[35362] <= 16'b1111111111110010;
        weights1[35363] <= 16'b1111111111111000;
        weights1[35364] <= 16'b0000000000000000;
        weights1[35365] <= 16'b0000000000000000;
        weights1[35366] <= 16'b0000000000000000;
        weights1[35367] <= 16'b1111111111111011;
        weights1[35368] <= 16'b1111111111110101;
        weights1[35369] <= 16'b1111111111110000;
        weights1[35370] <= 16'b1111111111101011;
        weights1[35371] <= 16'b1111111111010111;
        weights1[35372] <= 16'b1111111111001100;
        weights1[35373] <= 16'b1111111111000011;
        weights1[35374] <= 16'b1111111110111010;
        weights1[35375] <= 16'b0000000000000010;
        weights1[35376] <= 16'b0000000000010001;
        weights1[35377] <= 16'b0000000000011010;
        weights1[35378] <= 16'b0000000000011000;
        weights1[35379] <= 16'b0000000000101011;
        weights1[35380] <= 16'b0000000000101011;
        weights1[35381] <= 16'b0000000000100111;
        weights1[35382] <= 16'b0000000000011000;
        weights1[35383] <= 16'b0000000000010011;
        weights1[35384] <= 16'b1111111111011100;
        weights1[35385] <= 16'b1111111111011000;
        weights1[35386] <= 16'b1111111111010101;
        weights1[35387] <= 16'b1111111111011000;
        weights1[35388] <= 16'b1111111111010001;
        weights1[35389] <= 16'b1111111111100011;
        weights1[35390] <= 16'b1111111111101000;
        weights1[35391] <= 16'b1111111111110101;
        weights1[35392] <= 16'b0000000000000000;
        weights1[35393] <= 16'b0000000000000000;
        weights1[35394] <= 16'b0000000000000000;
        weights1[35395] <= 16'b1111111111111010;
        weights1[35396] <= 16'b1111111111101111;
        weights1[35397] <= 16'b1111111111100100;
        weights1[35398] <= 16'b1111111111011010;
        weights1[35399] <= 16'b1111111111000111;
        weights1[35400] <= 16'b1111111110100110;
        weights1[35401] <= 16'b1111111110111110;
        weights1[35402] <= 16'b1111111111001010;
        weights1[35403] <= 16'b0000000000000101;
        weights1[35404] <= 16'b1111111111111010;
        weights1[35405] <= 16'b0000000000010100;
        weights1[35406] <= 16'b1111111111111101;
        weights1[35407] <= 16'b0000000000011001;
        weights1[35408] <= 16'b0000000000001110;
        weights1[35409] <= 16'b0000000000011111;
        weights1[35410] <= 16'b0000000000010000;
        weights1[35411] <= 16'b1111111111101101;
        weights1[35412] <= 16'b1111111111000100;
        weights1[35413] <= 16'b1111111111001110;
        weights1[35414] <= 16'b1111111110111000;
        weights1[35415] <= 16'b1111111110101001;
        weights1[35416] <= 16'b1111111111000001;
        weights1[35417] <= 16'b1111111111100000;
        weights1[35418] <= 16'b1111111111100110;
        weights1[35419] <= 16'b1111111111110101;
        weights1[35420] <= 16'b1111111111111111;
        weights1[35421] <= 16'b1111111111111011;
        weights1[35422] <= 16'b1111111111110110;
        weights1[35423] <= 16'b1111111111110100;
        weights1[35424] <= 16'b1111111111101011;
        weights1[35425] <= 16'b1111111111011011;
        weights1[35426] <= 16'b1111111111010100;
        weights1[35427] <= 16'b1111111110101001;
        weights1[35428] <= 16'b1111111110110100;
        weights1[35429] <= 16'b1111111111011010;
        weights1[35430] <= 16'b0000000000000100;
        weights1[35431] <= 16'b0000000001000010;
        weights1[35432] <= 16'b0000000000011010;
        weights1[35433] <= 16'b0000000000001000;
        weights1[35434] <= 16'b0000000000011001;
        weights1[35435] <= 16'b0000000000010110;
        weights1[35436] <= 16'b0000000000001010;
        weights1[35437] <= 16'b0000000000011101;
        weights1[35438] <= 16'b1111111111101101;
        weights1[35439] <= 16'b1111111111100011;
        weights1[35440] <= 16'b1111111111010100;
        weights1[35441] <= 16'b1111111111001000;
        weights1[35442] <= 16'b1111111110101010;
        weights1[35443] <= 16'b1111111111000011;
        weights1[35444] <= 16'b1111111111011010;
        weights1[35445] <= 16'b1111111111101010;
        weights1[35446] <= 16'b1111111111101111;
        weights1[35447] <= 16'b1111111111110100;
        weights1[35448] <= 16'b1111111111111110;
        weights1[35449] <= 16'b1111111111111001;
        weights1[35450] <= 16'b1111111111110010;
        weights1[35451] <= 16'b1111111111101011;
        weights1[35452] <= 16'b1111111111100011;
        weights1[35453] <= 16'b1111111111010100;
        weights1[35454] <= 16'b1111111110111110;
        weights1[35455] <= 16'b1111111110110000;
        weights1[35456] <= 16'b1111111110100000;
        weights1[35457] <= 16'b1111111111011010;
        weights1[35458] <= 16'b0000000000010100;
        weights1[35459] <= 16'b0000000000010100;
        weights1[35460] <= 16'b0000000000000001;
        weights1[35461] <= 16'b0000000000011101;
        weights1[35462] <= 16'b0000000000011101;
        weights1[35463] <= 16'b1111111111101111;
        weights1[35464] <= 16'b1111111111011101;
        weights1[35465] <= 16'b1111111111110100;
        weights1[35466] <= 16'b1111111110111101;
        weights1[35467] <= 16'b1111111111010110;
        weights1[35468] <= 16'b1111111111011010;
        weights1[35469] <= 16'b1111111111011101;
        weights1[35470] <= 16'b1111111111100110;
        weights1[35471] <= 16'b1111111111111001;
        weights1[35472] <= 16'b1111111111110110;
        weights1[35473] <= 16'b1111111111101000;
        weights1[35474] <= 16'b1111111111111101;
        weights1[35475] <= 16'b1111111111110000;
        weights1[35476] <= 16'b1111111111111110;
        weights1[35477] <= 16'b1111111111111010;
        weights1[35478] <= 16'b1111111111110110;
        weights1[35479] <= 16'b1111111111101101;
        weights1[35480] <= 16'b1111111111101110;
        weights1[35481] <= 16'b1111111111011010;
        weights1[35482] <= 16'b1111111110111111;
        weights1[35483] <= 16'b1111111110101011;
        weights1[35484] <= 16'b1111111110110001;
        weights1[35485] <= 16'b0000000000010110;
        weights1[35486] <= 16'b0000000000011101;
        weights1[35487] <= 16'b0000000000110010;
        weights1[35488] <= 16'b0000000000001101;
        weights1[35489] <= 16'b0000000000001111;
        weights1[35490] <= 16'b0000000000001110;
        weights1[35491] <= 16'b1111111111111101;
        weights1[35492] <= 16'b1111111111100111;
        weights1[35493] <= 16'b1111111111011010;
        weights1[35494] <= 16'b1111111111101000;
        weights1[35495] <= 16'b1111111111011110;
        weights1[35496] <= 16'b1111111111101101;
        weights1[35497] <= 16'b1111111111011110;
        weights1[35498] <= 16'b1111111111110011;
        weights1[35499] <= 16'b1111111111110001;
        weights1[35500] <= 16'b0000000000000110;
        weights1[35501] <= 16'b0000000000000100;
        weights1[35502] <= 16'b1111111111111101;
        weights1[35503] <= 16'b1111111111110111;
        weights1[35504] <= 16'b1111111111111101;
        weights1[35505] <= 16'b1111111111110110;
        weights1[35506] <= 16'b1111111111110001;
        weights1[35507] <= 16'b1111111111101001;
        weights1[35508] <= 16'b1111111111100111;
        weights1[35509] <= 16'b1111111111010011;
        weights1[35510] <= 16'b1111111111000001;
        weights1[35511] <= 16'b1111111110011001;
        weights1[35512] <= 16'b1111111111001100;
        weights1[35513] <= 16'b0000000000000111;
        weights1[35514] <= 16'b0000000000001010;
        weights1[35515] <= 16'b0000000000011101;
        weights1[35516] <= 16'b0000000000001111;
        weights1[35517] <= 16'b0000000000010101;
        weights1[35518] <= 16'b0000000000000111;
        weights1[35519] <= 16'b1111111111011010;
        weights1[35520] <= 16'b1111111111001111;
        weights1[35521] <= 16'b1111111111010010;
        weights1[35522] <= 16'b1111111111011001;
        weights1[35523] <= 16'b1111111111100001;
        weights1[35524] <= 16'b1111111111101111;
        weights1[35525] <= 16'b1111111111111011;
        weights1[35526] <= 16'b1111111111111101;
        weights1[35527] <= 16'b0000000000000101;
        weights1[35528] <= 16'b0000000000001110;
        weights1[35529] <= 16'b0000000000000000;
        weights1[35530] <= 16'b0000000000001000;
        weights1[35531] <= 16'b0000000000000000;
        weights1[35532] <= 16'b0000000000000000;
        weights1[35533] <= 16'b1111111111111100;
        weights1[35534] <= 16'b1111111111110011;
        weights1[35535] <= 16'b1111111111101010;
        weights1[35536] <= 16'b1111111111100101;
        weights1[35537] <= 16'b1111111111000110;
        weights1[35538] <= 16'b1111111110101001;
        weights1[35539] <= 16'b1111111110011100;
        weights1[35540] <= 16'b1111111111111001;
        weights1[35541] <= 16'b0000000000010001;
        weights1[35542] <= 16'b0000000000001110;
        weights1[35543] <= 16'b0000000000000100;
        weights1[35544] <= 16'b0000000000001111;
        weights1[35545] <= 16'b0000000000000111;
        weights1[35546] <= 16'b1111111111100100;
        weights1[35547] <= 16'b1111111111000100;
        weights1[35548] <= 16'b1111111111011101;
        weights1[35549] <= 16'b1111111111100101;
        weights1[35550] <= 16'b1111111111100001;
        weights1[35551] <= 16'b1111111111110010;
        weights1[35552] <= 16'b1111111111110010;
        weights1[35553] <= 16'b0000000000011101;
        weights1[35554] <= 16'b0000000000001011;
        weights1[35555] <= 16'b0000000000011001;
        weights1[35556] <= 16'b0000000000010001;
        weights1[35557] <= 16'b0000000000001010;
        weights1[35558] <= 16'b0000000000001011;
        weights1[35559] <= 16'b0000000000001000;
        weights1[35560] <= 16'b1111111111111110;
        weights1[35561] <= 16'b1111111111110110;
        weights1[35562] <= 16'b1111111111110010;
        weights1[35563] <= 16'b1111111111101100;
        weights1[35564] <= 16'b1111111111011010;
        weights1[35565] <= 16'b1111111111000101;
        weights1[35566] <= 16'b1111111110010111;
        weights1[35567] <= 16'b1111111111110010;
        weights1[35568] <= 16'b1111111111101001;
        weights1[35569] <= 16'b0000000000011001;
        weights1[35570] <= 16'b0000000000001011;
        weights1[35571] <= 16'b0000000000011110;
        weights1[35572] <= 16'b0000000000001001;
        weights1[35573] <= 16'b0000000000000111;
        weights1[35574] <= 16'b1111111111011010;
        weights1[35575] <= 16'b1111111111000101;
        weights1[35576] <= 16'b1111111111110101;
        weights1[35577] <= 16'b1111111111111111;
        weights1[35578] <= 16'b1111111111111111;
        weights1[35579] <= 16'b1111111111110100;
        weights1[35580] <= 16'b0000000000001100;
        weights1[35581] <= 16'b0000000000010100;
        weights1[35582] <= 16'b0000000000011001;
        weights1[35583] <= 16'b0000000000000100;
        weights1[35584] <= 16'b0000000000000011;
        weights1[35585] <= 16'b1111111111101011;
        weights1[35586] <= 16'b0000000000000111;
        weights1[35587] <= 16'b0000000000000100;
        weights1[35588] <= 16'b1111111111111111;
        weights1[35589] <= 16'b1111111111111010;
        weights1[35590] <= 16'b1111111111110011;
        weights1[35591] <= 16'b1111111111110010;
        weights1[35592] <= 16'b1111111111010110;
        weights1[35593] <= 16'b1111111110111101;
        weights1[35594] <= 16'b1111111111001100;
        weights1[35595] <= 16'b1111111111101100;
        weights1[35596] <= 16'b1111111111110110;
        weights1[35597] <= 16'b0000000000001010;
        weights1[35598] <= 16'b0000000000000010;
        weights1[35599] <= 16'b0000000000011110;
        weights1[35600] <= 16'b0000000000100100;
        weights1[35601] <= 16'b1111111111101100;
        weights1[35602] <= 16'b1111111111000001;
        weights1[35603] <= 16'b1111111111001011;
        weights1[35604] <= 16'b0000000000001000;
        weights1[35605] <= 16'b1111111111101000;
        weights1[35606] <= 16'b1111111111111100;
        weights1[35607] <= 16'b0000000000010011;
        weights1[35608] <= 16'b0000000000001100;
        weights1[35609] <= 16'b1111111111111100;
        weights1[35610] <= 16'b0000000000001111;
        weights1[35611] <= 16'b0000000000001011;
        weights1[35612] <= 16'b1111111111110001;
        weights1[35613] <= 16'b0000000000001010;
        weights1[35614] <= 16'b0000000000010011;
        weights1[35615] <= 16'b0000000000001001;
        weights1[35616] <= 16'b1111111111111111;
        weights1[35617] <= 16'b1111111111111011;
        weights1[35618] <= 16'b1111111111110100;
        weights1[35619] <= 16'b1111111111100111;
        weights1[35620] <= 16'b1111111111010010;
        weights1[35621] <= 16'b1111111111000111;
        weights1[35622] <= 16'b1111111111100101;
        weights1[35623] <= 16'b1111111111101110;
        weights1[35624] <= 16'b0000000000001011;
        weights1[35625] <= 16'b0000000000001110;
        weights1[35626] <= 16'b1111111111111110;
        weights1[35627] <= 16'b0000000000101110;
        weights1[35628] <= 16'b0000000000010010;
        weights1[35629] <= 16'b1111111111101111;
        weights1[35630] <= 16'b1111111111000010;
        weights1[35631] <= 16'b1111111111110001;
        weights1[35632] <= 16'b1111111111111101;
        weights1[35633] <= 16'b0000000000000000;
        weights1[35634] <= 16'b1111111111111110;
        weights1[35635] <= 16'b1111111111110101;
        weights1[35636] <= 16'b1111111111111001;
        weights1[35637] <= 16'b0000000000000010;
        weights1[35638] <= 16'b0000000000000001;
        weights1[35639] <= 16'b1111111111111111;
        weights1[35640] <= 16'b0000000000010001;
        weights1[35641] <= 16'b1111111111101100;
        weights1[35642] <= 16'b0000000000000000;
        weights1[35643] <= 16'b0000000000001100;
        weights1[35644] <= 16'b1111111111111110;
        weights1[35645] <= 16'b1111111111110101;
        weights1[35646] <= 16'b1111111111101111;
        weights1[35647] <= 16'b1111111111100001;
        weights1[35648] <= 16'b1111111111100100;
        weights1[35649] <= 16'b1111111111010100;
        weights1[35650] <= 16'b1111111111110100;
        weights1[35651] <= 16'b0000000000011001;
        weights1[35652] <= 16'b1111111111111011;
        weights1[35653] <= 16'b0000000000000001;
        weights1[35654] <= 16'b0000000000011000;
        weights1[35655] <= 16'b0000000000101000;
        weights1[35656] <= 16'b0000000000000110;
        weights1[35657] <= 16'b1111111111100100;
        weights1[35658] <= 16'b1111111111001101;
        weights1[35659] <= 16'b1111111111110111;
        weights1[35660] <= 16'b1111111111110111;
        weights1[35661] <= 16'b0000000000000010;
        weights1[35662] <= 16'b1111111111110101;
        weights1[35663] <= 16'b0000000000011011;
        weights1[35664] <= 16'b1111111111111101;
        weights1[35665] <= 16'b0000000000011111;
        weights1[35666] <= 16'b0000000000001101;
        weights1[35667] <= 16'b1111111111110000;
        weights1[35668] <= 16'b0000000000001111;
        weights1[35669] <= 16'b0000000000001011;
        weights1[35670] <= 16'b0000000000000110;
        weights1[35671] <= 16'b1111111111111111;
        weights1[35672] <= 16'b1111111111111000;
        weights1[35673] <= 16'b1111111111110100;
        weights1[35674] <= 16'b1111111111110000;
        weights1[35675] <= 16'b1111111111100000;
        weights1[35676] <= 16'b1111111111001011;
        weights1[35677] <= 16'b1111111111100111;
        weights1[35678] <= 16'b0000000000000110;
        weights1[35679] <= 16'b0000000000001100;
        weights1[35680] <= 16'b0000000000001011;
        weights1[35681] <= 16'b0000000000010000;
        weights1[35682] <= 16'b0000000000010110;
        weights1[35683] <= 16'b0000000000100110;
        weights1[35684] <= 16'b0000000000000011;
        weights1[35685] <= 16'b1111111111101010;
        weights1[35686] <= 16'b1111111111100101;
        weights1[35687] <= 16'b1111111111111010;
        weights1[35688] <= 16'b0000000000011010;
        weights1[35689] <= 16'b0000000000001000;
        weights1[35690] <= 16'b1111111111111001;
        weights1[35691] <= 16'b1111111111110000;
        weights1[35692] <= 16'b0000000000100001;
        weights1[35693] <= 16'b0000000000001011;
        weights1[35694] <= 16'b0000000000011001;
        weights1[35695] <= 16'b1111111111111100;
        weights1[35696] <= 16'b0000000000011001;
        weights1[35697] <= 16'b1111111111101011;
        weights1[35698] <= 16'b0000000000010100;
        weights1[35699] <= 16'b0000000000001000;
        weights1[35700] <= 16'b1111111111110100;
        weights1[35701] <= 16'b1111111111101111;
        weights1[35702] <= 16'b1111111111101010;
        weights1[35703] <= 16'b1111111111100000;
        weights1[35704] <= 16'b1111111111100101;
        weights1[35705] <= 16'b1111111111101101;
        weights1[35706] <= 16'b1111111111111100;
        weights1[35707] <= 16'b0000000000001001;
        weights1[35708] <= 16'b0000000000100110;
        weights1[35709] <= 16'b0000000000100001;
        weights1[35710] <= 16'b0000000000010111;
        weights1[35711] <= 16'b0000000000101110;
        weights1[35712] <= 16'b1111111111111101;
        weights1[35713] <= 16'b1111111111101010;
        weights1[35714] <= 16'b1111111111110110;
        weights1[35715] <= 16'b1111111111101000;
        weights1[35716] <= 16'b1111111111111100;
        weights1[35717] <= 16'b1111111111111011;
        weights1[35718] <= 16'b1111111111111110;
        weights1[35719] <= 16'b0000000000001101;
        weights1[35720] <= 16'b1111111111111111;
        weights1[35721] <= 16'b0000000000100100;
        weights1[35722] <= 16'b0000000000001111;
        weights1[35723] <= 16'b0000000000100011;
        weights1[35724] <= 16'b0000000000000111;
        weights1[35725] <= 16'b0000000000001110;
        weights1[35726] <= 16'b1111111111111101;
        weights1[35727] <= 16'b0000000000010011;
        weights1[35728] <= 16'b1111111111110101;
        weights1[35729] <= 16'b1111111111110000;
        weights1[35730] <= 16'b1111111111110001;
        weights1[35731] <= 16'b1111111111011110;
        weights1[35732] <= 16'b1111111111110010;
        weights1[35733] <= 16'b0000000000010101;
        weights1[35734] <= 16'b0000000000001111;
        weights1[35735] <= 16'b0000000000001110;
        weights1[35736] <= 16'b0000000000001110;
        weights1[35737] <= 16'b1111111111111100;
        weights1[35738] <= 16'b1111111111111010;
        weights1[35739] <= 16'b0000000000100010;
        weights1[35740] <= 16'b1111111111111000;
        weights1[35741] <= 16'b1111111111111000;
        weights1[35742] <= 16'b0000000000001001;
        weights1[35743] <= 16'b0000000000000100;
        weights1[35744] <= 16'b1111111111100010;
        weights1[35745] <= 16'b1111111111111000;
        weights1[35746] <= 16'b0000000000000010;
        weights1[35747] <= 16'b0000000000000101;
        weights1[35748] <= 16'b0000000000001101;
        weights1[35749] <= 16'b0000000000001010;
        weights1[35750] <= 16'b0000000000000100;
        weights1[35751] <= 16'b1111111111111010;
        weights1[35752] <= 16'b1111111111110000;
        weights1[35753] <= 16'b0000000000000100;
        weights1[35754] <= 16'b0000000000001011;
        weights1[35755] <= 16'b0000000000010000;
        weights1[35756] <= 16'b1111111111110111;
        weights1[35757] <= 16'b1111111111110001;
        weights1[35758] <= 16'b1111111111101110;
        weights1[35759] <= 16'b1111111111100011;
        weights1[35760] <= 16'b1111111111110111;
        weights1[35761] <= 16'b0000000000010001;
        weights1[35762] <= 16'b0000000000000101;
        weights1[35763] <= 16'b0000000000001001;
        weights1[35764] <= 16'b0000000000001100;
        weights1[35765] <= 16'b0000000000000110;
        weights1[35766] <= 16'b1111111111111100;
        weights1[35767] <= 16'b0000000000011011;
        weights1[35768] <= 16'b0000000000001010;
        weights1[35769] <= 16'b0000000000000101;
        weights1[35770] <= 16'b0000000000000000;
        weights1[35771] <= 16'b1111111111100111;
        weights1[35772] <= 16'b1111111111111010;
        weights1[35773] <= 16'b0000000000001111;
        weights1[35774] <= 16'b1111111111111110;
        weights1[35775] <= 16'b0000000000001010;
        weights1[35776] <= 16'b0000000000000100;
        weights1[35777] <= 16'b1111111111111111;
        weights1[35778] <= 16'b0000000000010001;
        weights1[35779] <= 16'b0000000000000010;
        weights1[35780] <= 16'b0000000000000010;
        weights1[35781] <= 16'b0000000000000111;
        weights1[35782] <= 16'b0000000000000111;
        weights1[35783] <= 16'b0000000000001100;
        weights1[35784] <= 16'b1111111111111101;
        weights1[35785] <= 16'b1111111111110001;
        weights1[35786] <= 16'b1111111111101110;
        weights1[35787] <= 16'b1111111111101010;
        weights1[35788] <= 16'b1111111111111101;
        weights1[35789] <= 16'b1111111111111001;
        weights1[35790] <= 16'b1111111111110100;
        weights1[35791] <= 16'b1111111111111110;
        weights1[35792] <= 16'b0000000000011001;
        weights1[35793] <= 16'b0000000000001011;
        weights1[35794] <= 16'b1111111111111111;
        weights1[35795] <= 16'b0000000000000010;
        weights1[35796] <= 16'b1111111111111100;
        weights1[35797] <= 16'b1111111111111010;
        weights1[35798] <= 16'b0000000000000100;
        weights1[35799] <= 16'b0000000000001010;
        weights1[35800] <= 16'b1111111111101111;
        weights1[35801] <= 16'b1111111111111000;
        weights1[35802] <= 16'b1111111111110100;
        weights1[35803] <= 16'b1111111111011100;
        weights1[35804] <= 16'b1111111111100111;
        weights1[35805] <= 16'b1111111111001101;
        weights1[35806] <= 16'b0000000000000100;
        weights1[35807] <= 16'b1111111111101010;
        weights1[35808] <= 16'b0000000000000010;
        weights1[35809] <= 16'b0000000000000001;
        weights1[35810] <= 16'b0000000000000110;
        weights1[35811] <= 16'b1111111111110101;
        weights1[35812] <= 16'b1111111111111111;
        weights1[35813] <= 16'b1111111111110100;
        weights1[35814] <= 16'b1111111111100111;
        weights1[35815] <= 16'b1111111111101000;
        weights1[35816] <= 16'b1111111111110001;
        weights1[35817] <= 16'b0000000000000011;
        weights1[35818] <= 16'b1111111111101011;
        weights1[35819] <= 16'b1111111111111011;
        weights1[35820] <= 16'b1111111111111110;
        weights1[35821] <= 16'b0000000000001000;
        weights1[35822] <= 16'b0000000000010001;
        weights1[35823] <= 16'b0000000000100000;
        weights1[35824] <= 16'b0000000000011000;
        weights1[35825] <= 16'b0000000000001110;
        weights1[35826] <= 16'b1111111111111100;
        weights1[35827] <= 16'b0000000000000001;
        weights1[35828] <= 16'b1111111111110001;
        weights1[35829] <= 16'b1111111111101000;
        weights1[35830] <= 16'b0000000000010101;
        weights1[35831] <= 16'b0000000000000110;
        weights1[35832] <= 16'b1111111111111101;
        weights1[35833] <= 16'b0000000000000101;
        weights1[35834] <= 16'b1111111111011100;
        weights1[35835] <= 16'b1111111111110110;
        weights1[35836] <= 16'b1111111111111100;
        weights1[35837] <= 16'b1111111111110010;
        weights1[35838] <= 16'b1111111111111001;
        weights1[35839] <= 16'b1111111111110111;
        weights1[35840] <= 16'b1111111111111010;
        weights1[35841] <= 16'b1111111111111001;
        weights1[35842] <= 16'b1111111111101000;
        weights1[35843] <= 16'b1111111111101010;
        weights1[35844] <= 16'b1111111111111110;
        weights1[35845] <= 16'b0000000000001001;
        weights1[35846] <= 16'b0000000000000111;
        weights1[35847] <= 16'b1111111111110001;
        weights1[35848] <= 16'b0000000000000101;
        weights1[35849] <= 16'b0000000000001001;
        weights1[35850] <= 16'b0000000000010111;
        weights1[35851] <= 16'b0000000000010001;
        weights1[35852] <= 16'b0000000000011111;
        weights1[35853] <= 16'b0000000000010100;
        weights1[35854] <= 16'b1111111111111101;
        weights1[35855] <= 16'b0000000000001010;
        weights1[35856] <= 16'b1111111111110011;
        weights1[35857] <= 16'b1111111111110111;
        weights1[35858] <= 16'b1111111111110010;
        weights1[35859] <= 16'b1111111111110111;
        weights1[35860] <= 16'b0000000000000001;
        weights1[35861] <= 16'b0000000000000100;
        weights1[35862] <= 16'b1111111111101101;
        weights1[35863] <= 16'b1111111111101011;
        weights1[35864] <= 16'b1111111111101111;
        weights1[35865] <= 16'b1111111111101100;
        weights1[35866] <= 16'b1111111111110011;
        weights1[35867] <= 16'b1111111111110001;
        weights1[35868] <= 16'b1111111111111011;
        weights1[35869] <= 16'b1111111111111000;
        weights1[35870] <= 16'b1111111111101101;
        weights1[35871] <= 16'b1111111111011111;
        weights1[35872] <= 16'b1111111111101001;
        weights1[35873] <= 16'b0000000000000010;
        weights1[35874] <= 16'b1111111111110111;
        weights1[35875] <= 16'b0000000000001001;
        weights1[35876] <= 16'b0000000000000001;
        weights1[35877] <= 16'b0000000000000110;
        weights1[35878] <= 16'b0000000000001110;
        weights1[35879] <= 16'b0000000000011001;
        weights1[35880] <= 16'b0000000000011011;
        weights1[35881] <= 16'b0000000000010011;
        weights1[35882] <= 16'b0000000000000111;
        weights1[35883] <= 16'b0000000000010110;
        weights1[35884] <= 16'b1111111111110011;
        weights1[35885] <= 16'b1111111111110110;
        weights1[35886] <= 16'b1111111111111111;
        weights1[35887] <= 16'b1111111111100100;
        weights1[35888] <= 16'b0000000000001100;
        weights1[35889] <= 16'b1111111111101010;
        weights1[35890] <= 16'b1111111111100111;
        weights1[35891] <= 16'b0000000000000100;
        weights1[35892] <= 16'b1111111111110100;
        weights1[35893] <= 16'b1111111111110110;
        weights1[35894] <= 16'b1111111111111000;
        weights1[35895] <= 16'b1111111111101110;
        weights1[35896] <= 16'b1111111111111000;
        weights1[35897] <= 16'b1111111111110110;
        weights1[35898] <= 16'b1111111111110010;
        weights1[35899] <= 16'b1111111111100101;
        weights1[35900] <= 16'b1111111111011111;
        weights1[35901] <= 16'b1111111111110011;
        weights1[35902] <= 16'b1111111111110011;
        weights1[35903] <= 16'b0000000000001100;
        weights1[35904] <= 16'b1111111111110001;
        weights1[35905] <= 16'b0000000000010011;
        weights1[35906] <= 16'b0000000000000100;
        weights1[35907] <= 16'b0000000000010000;
        weights1[35908] <= 16'b0000000000010100;
        weights1[35909] <= 16'b0000000000001010;
        weights1[35910] <= 16'b0000000000001000;
        weights1[35911] <= 16'b0000000000001010;
        weights1[35912] <= 16'b0000000000000001;
        weights1[35913] <= 16'b1111111111110000;
        weights1[35914] <= 16'b0000000000001100;
        weights1[35915] <= 16'b0000000000000111;
        weights1[35916] <= 16'b1111111111111010;
        weights1[35917] <= 16'b1111111111101101;
        weights1[35918] <= 16'b1111111111110110;
        weights1[35919] <= 16'b1111111111110000;
        weights1[35920] <= 16'b1111111111101111;
        weights1[35921] <= 16'b1111111111101111;
        weights1[35922] <= 16'b1111111111111000;
        weights1[35923] <= 16'b1111111111110101;
        weights1[35924] <= 16'b1111111111111101;
        weights1[35925] <= 16'b1111111111110111;
        weights1[35926] <= 16'b1111111111110000;
        weights1[35927] <= 16'b1111111111110111;
        weights1[35928] <= 16'b1111111111101101;
        weights1[35929] <= 16'b1111111111110001;
        weights1[35930] <= 16'b1111111111110010;
        weights1[35931] <= 16'b1111111111110010;
        weights1[35932] <= 16'b0000000000011111;
        weights1[35933] <= 16'b0000000000000100;
        weights1[35934] <= 16'b0000000000000111;
        weights1[35935] <= 16'b0000000000101000;
        weights1[35936] <= 16'b0000000000010110;
        weights1[35937] <= 16'b0000000000011011;
        weights1[35938] <= 16'b0000000000000100;
        weights1[35939] <= 16'b0000000000101011;
        weights1[35940] <= 16'b0000000000010000;
        weights1[35941] <= 16'b0000000000000000;
        weights1[35942] <= 16'b0000000000001010;
        weights1[35943] <= 16'b0000000000100000;
        weights1[35944] <= 16'b0000000000000001;
        weights1[35945] <= 16'b1111111111111010;
        weights1[35946] <= 16'b1111111111101111;
        weights1[35947] <= 16'b1111111111110110;
        weights1[35948] <= 16'b1111111111101001;
        weights1[35949] <= 16'b1111111111111001;
        weights1[35950] <= 16'b1111111111111001;
        weights1[35951] <= 16'b1111111111110101;
        weights1[35952] <= 16'b0000000000000000;
        weights1[35953] <= 16'b0000000000000001;
        weights1[35954] <= 16'b1111111111111001;
        weights1[35955] <= 16'b1111111111110010;
        weights1[35956] <= 16'b1111111111110101;
        weights1[35957] <= 16'b1111111111100110;
        weights1[35958] <= 16'b1111111111101000;
        weights1[35959] <= 16'b1111111111110110;
        weights1[35960] <= 16'b1111111111110001;
        weights1[35961] <= 16'b0000000000010100;
        weights1[35962] <= 16'b0000000000010101;
        weights1[35963] <= 16'b0000000000010011;
        weights1[35964] <= 16'b0000000000011010;
        weights1[35965] <= 16'b0000000000011010;
        weights1[35966] <= 16'b0000000000010000;
        weights1[35967] <= 16'b0000000000100011;
        weights1[35968] <= 16'b0000000000011100;
        weights1[35969] <= 16'b1111111111110001;
        weights1[35970] <= 16'b1111111111101010;
        weights1[35971] <= 16'b1111111111110010;
        weights1[35972] <= 16'b1111111111101001;
        weights1[35973] <= 16'b1111111111110111;
        weights1[35974] <= 16'b0000000000000110;
        weights1[35975] <= 16'b1111111111110111;
        weights1[35976] <= 16'b1111111111110101;
        weights1[35977] <= 16'b1111111111110101;
        weights1[35978] <= 16'b1111111111110111;
        weights1[35979] <= 16'b1111111111110100;
        weights1[35980] <= 16'b0000000000000000;
        weights1[35981] <= 16'b1111111111111111;
        weights1[35982] <= 16'b1111111111111100;
        weights1[35983] <= 16'b1111111111110101;
        weights1[35984] <= 16'b1111111111110001;
        weights1[35985] <= 16'b1111111111010111;
        weights1[35986] <= 16'b1111111111010111;
        weights1[35987] <= 16'b1111111111001110;
        weights1[35988] <= 16'b1111111111101110;
        weights1[35989] <= 16'b1111111111100010;
        weights1[35990] <= 16'b1111111111110001;
        weights1[35991] <= 16'b1111111111110010;
        weights1[35992] <= 16'b1111111111111010;
        weights1[35993] <= 16'b1111111111101101;
        weights1[35994] <= 16'b0000000000000000;
        weights1[35995] <= 16'b1111111111111101;
        weights1[35996] <= 16'b1111111111111001;
        weights1[35997] <= 16'b0000000000010010;
        weights1[35998] <= 16'b1111111111111101;
        weights1[35999] <= 16'b1111111111110101;
        weights1[36000] <= 16'b1111111111110101;
        weights1[36001] <= 16'b1111111111110011;
        weights1[36002] <= 16'b1111111111111010;
        weights1[36003] <= 16'b1111111111111101;
        weights1[36004] <= 16'b1111111111110001;
        weights1[36005] <= 16'b1111111111110110;
        weights1[36006] <= 16'b1111111111110100;
        weights1[36007] <= 16'b1111111111110110;
        weights1[36008] <= 16'b0000000000000000;
        weights1[36009] <= 16'b0000000000000001;
        weights1[36010] <= 16'b1111111111111100;
        weights1[36011] <= 16'b1111111111110101;
        weights1[36012] <= 16'b1111111111110001;
        weights1[36013] <= 16'b1111111111101110;
        weights1[36014] <= 16'b1111111111010011;
        weights1[36015] <= 16'b1111111111001111;
        weights1[36016] <= 16'b1111111111010001;
        weights1[36017] <= 16'b1111111111010111;
        weights1[36018] <= 16'b1111111111011011;
        weights1[36019] <= 16'b1111111111101011;
        weights1[36020] <= 16'b1111111111110001;
        weights1[36021] <= 16'b1111111111101011;
        weights1[36022] <= 16'b1111111111101011;
        weights1[36023] <= 16'b1111111111101001;
        weights1[36024] <= 16'b1111111111100110;
        weights1[36025] <= 16'b1111111111100100;
        weights1[36026] <= 16'b1111111111111110;
        weights1[36027] <= 16'b1111111111110000;
        weights1[36028] <= 16'b1111111111110000;
        weights1[36029] <= 16'b1111111111101010;
        weights1[36030] <= 16'b1111111111110001;
        weights1[36031] <= 16'b1111111111110011;
        weights1[36032] <= 16'b1111111111110011;
        weights1[36033] <= 16'b1111111111111001;
        weights1[36034] <= 16'b1111111111110111;
        weights1[36035] <= 16'b1111111111111010;
        weights1[36036] <= 16'b1111111111111111;
        weights1[36037] <= 16'b1111111111111110;
        weights1[36038] <= 16'b1111111111111000;
        weights1[36039] <= 16'b1111111111111001;
        weights1[36040] <= 16'b1111111111101101;
        weights1[36041] <= 16'b1111111111100101;
        weights1[36042] <= 16'b1111111111100111;
        weights1[36043] <= 16'b1111111111011100;
        weights1[36044] <= 16'b1111111111001111;
        weights1[36045] <= 16'b1111111111001011;
        weights1[36046] <= 16'b1111111111011011;
        weights1[36047] <= 16'b1111111111000101;
        weights1[36048] <= 16'b1111111111001000;
        weights1[36049] <= 16'b1111111111000011;
        weights1[36050] <= 16'b1111111110111100;
        weights1[36051] <= 16'b1111111111001101;
        weights1[36052] <= 16'b1111111111001011;
        weights1[36053] <= 16'b1111111111100000;
        weights1[36054] <= 16'b1111111111100000;
        weights1[36055] <= 16'b1111111111011110;
        weights1[36056] <= 16'b1111111111101011;
        weights1[36057] <= 16'b1111111111100110;
        weights1[36058] <= 16'b1111111111110001;
        weights1[36059] <= 16'b1111111111110011;
        weights1[36060] <= 16'b1111111111110110;
        weights1[36061] <= 16'b1111111111111101;
        weights1[36062] <= 16'b1111111111111100;
        weights1[36063] <= 16'b1111111111111101;
        weights1[36064] <= 16'b0000000000000000;
        weights1[36065] <= 16'b0000000000000000;
        weights1[36066] <= 16'b0000000000000000;
        weights1[36067] <= 16'b0000000000000000;
        weights1[36068] <= 16'b0000000000000000;
        weights1[36069] <= 16'b0000000000000001;
        weights1[36070] <= 16'b1111111111111111;
        weights1[36071] <= 16'b1111111111111000;
        weights1[36072] <= 16'b1111111111110100;
        weights1[36073] <= 16'b1111111111101101;
        weights1[36074] <= 16'b1111111111101101;
        weights1[36075] <= 16'b1111111111100111;
        weights1[36076] <= 16'b1111111111101000;
        weights1[36077] <= 16'b1111111111100110;
        weights1[36078] <= 16'b1111111111100011;
        weights1[36079] <= 16'b1111111111100000;
        weights1[36080] <= 16'b1111111111010110;
        weights1[36081] <= 16'b1111111111011101;
        weights1[36082] <= 16'b1111111111010101;
        weights1[36083] <= 16'b1111111111101000;
        weights1[36084] <= 16'b1111111111110011;
        weights1[36085] <= 16'b1111111111111110;
        weights1[36086] <= 16'b0000000000001010;
        weights1[36087] <= 16'b0000000000001000;
        weights1[36088] <= 16'b0000000000000001;
        weights1[36089] <= 16'b0000000000000110;
        weights1[36090] <= 16'b0000000000000111;
        weights1[36091] <= 16'b0000000000000000;
        weights1[36092] <= 16'b0000000000000000;
        weights1[36093] <= 16'b0000000000000000;
        weights1[36094] <= 16'b1111111111111110;
        weights1[36095] <= 16'b1111111111111110;
        weights1[36096] <= 16'b1111111111111100;
        weights1[36097] <= 16'b1111111111111110;
        weights1[36098] <= 16'b1111111111111011;
        weights1[36099] <= 16'b1111111111111010;
        weights1[36100] <= 16'b1111111111110100;
        weights1[36101] <= 16'b1111111111111110;
        weights1[36102] <= 16'b1111111111110101;
        weights1[36103] <= 16'b1111111111011101;
        weights1[36104] <= 16'b1111111111011110;
        weights1[36105] <= 16'b1111111111100100;
        weights1[36106] <= 16'b1111111111100010;
        weights1[36107] <= 16'b1111111111010001;
        weights1[36108] <= 16'b1111111111100011;
        weights1[36109] <= 16'b1111111111011000;
        weights1[36110] <= 16'b1111111111011110;
        weights1[36111] <= 16'b1111111111110011;
        weights1[36112] <= 16'b1111111111111001;
        weights1[36113] <= 16'b1111111111101111;
        weights1[36114] <= 16'b0000000000000011;
        weights1[36115] <= 16'b0000000000001000;
        weights1[36116] <= 16'b0000000000000010;
        weights1[36117] <= 16'b0000000000000101;
        weights1[36118] <= 16'b0000000000000101;
        weights1[36119] <= 16'b1111111111111110;
        weights1[36120] <= 16'b0000000000000000;
        weights1[36121] <= 16'b0000000000000000;
        weights1[36122] <= 16'b1111111111111111;
        weights1[36123] <= 16'b1111111111111110;
        weights1[36124] <= 16'b1111111111111011;
        weights1[36125] <= 16'b1111111111111001;
        weights1[36126] <= 16'b1111111111111001;
        weights1[36127] <= 16'b1111111111111110;
        weights1[36128] <= 16'b0000000000000010;
        weights1[36129] <= 16'b1111111111110101;
        weights1[36130] <= 16'b1111111111110100;
        weights1[36131] <= 16'b1111111111110111;
        weights1[36132] <= 16'b1111111111100110;
        weights1[36133] <= 16'b1111111111101100;
        weights1[36134] <= 16'b1111111111100011;
        weights1[36135] <= 16'b1111111111111001;
        weights1[36136] <= 16'b1111111111111000;
        weights1[36137] <= 16'b1111111111100010;
        weights1[36138] <= 16'b0000000000000101;
        weights1[36139] <= 16'b1111111111101110;
        weights1[36140] <= 16'b1111111111110100;
        weights1[36141] <= 16'b1111111111111101;
        weights1[36142] <= 16'b0000000000010000;
        weights1[36143] <= 16'b0000000000000100;
        weights1[36144] <= 16'b0000000000000000;
        weights1[36145] <= 16'b0000000000011011;
        weights1[36146] <= 16'b0000000000010110;
        weights1[36147] <= 16'b0000000000001110;
        weights1[36148] <= 16'b1111111111111110;
        weights1[36149] <= 16'b1111111111111110;
        weights1[36150] <= 16'b1111111111111101;
        weights1[36151] <= 16'b1111111111111010;
        weights1[36152] <= 16'b1111111111111001;
        weights1[36153] <= 16'b1111111111111111;
        weights1[36154] <= 16'b1111111111110010;
        weights1[36155] <= 16'b0000000000000001;
        weights1[36156] <= 16'b1111111111111010;
        weights1[36157] <= 16'b0000000000000100;
        weights1[36158] <= 16'b1111111111101001;
        weights1[36159] <= 16'b0000000000000100;
        weights1[36160] <= 16'b1111111111101100;
        weights1[36161] <= 16'b1111111111111001;
        weights1[36162] <= 16'b1111111111111101;
        weights1[36163] <= 16'b0000000000000100;
        weights1[36164] <= 16'b0000000000000100;
        weights1[36165] <= 16'b1111111111111001;
        weights1[36166] <= 16'b0000000000011000;
        weights1[36167] <= 16'b0000000000101001;
        weights1[36168] <= 16'b0000000000011101;
        weights1[36169] <= 16'b0000000000011100;
        weights1[36170] <= 16'b0000000000010100;
        weights1[36171] <= 16'b0000000000010100;
        weights1[36172] <= 16'b1111111111111101;
        weights1[36173] <= 16'b0000000000010110;
        weights1[36174] <= 16'b0000000000101000;
        weights1[36175] <= 16'b0000000000011011;
        weights1[36176] <= 16'b1111111111111110;
        weights1[36177] <= 16'b1111111111111110;
        weights1[36178] <= 16'b0000000000000001;
        weights1[36179] <= 16'b1111111111111111;
        weights1[36180] <= 16'b1111111111101111;
        weights1[36181] <= 16'b1111111111110011;
        weights1[36182] <= 16'b1111111111110111;
        weights1[36183] <= 16'b1111111111111011;
        weights1[36184] <= 16'b1111111111111000;
        weights1[36185] <= 16'b1111111111110101;
        weights1[36186] <= 16'b1111111111101110;
        weights1[36187] <= 16'b1111111111111110;
        weights1[36188] <= 16'b1111111111110010;
        weights1[36189] <= 16'b1111111111110001;
        weights1[36190] <= 16'b1111111111111101;
        weights1[36191] <= 16'b0000000000000111;
        weights1[36192] <= 16'b1111111111111100;
        weights1[36193] <= 16'b0000000000010001;
        weights1[36194] <= 16'b0000000000011100;
        weights1[36195] <= 16'b0000000000011111;
        weights1[36196] <= 16'b1111111111110110;
        weights1[36197] <= 16'b0000000000010100;
        weights1[36198] <= 16'b0000000000010011;
        weights1[36199] <= 16'b0000000000011111;
        weights1[36200] <= 16'b0000000000100110;
        weights1[36201] <= 16'b0000000000010010;
        weights1[36202] <= 16'b0000000000011011;
        weights1[36203] <= 16'b0000000000100100;
        weights1[36204] <= 16'b1111111111111001;
        weights1[36205] <= 16'b1111111111111011;
        weights1[36206] <= 16'b1111111111111000;
        weights1[36207] <= 16'b1111111111110110;
        weights1[36208] <= 16'b1111111111101111;
        weights1[36209] <= 16'b1111111111011110;
        weights1[36210] <= 16'b1111111111111101;
        weights1[36211] <= 16'b1111111111100000;
        weights1[36212] <= 16'b0000000000001000;
        weights1[36213] <= 16'b1111111111111010;
        weights1[36214] <= 16'b0000000000010010;
        weights1[36215] <= 16'b0000000000000001;
        weights1[36216] <= 16'b1111111111111100;
        weights1[36217] <= 16'b0000000000001001;
        weights1[36218] <= 16'b0000000000001000;
        weights1[36219] <= 16'b0000000000000100;
        weights1[36220] <= 16'b0000000000100011;
        weights1[36221] <= 16'b0000000000001000;
        weights1[36222] <= 16'b0000000000011011;
        weights1[36223] <= 16'b0000000000001000;
        weights1[36224] <= 16'b0000000000011010;
        weights1[36225] <= 16'b0000000000100001;
        weights1[36226] <= 16'b0000000000101001;
        weights1[36227] <= 16'b0000000000110110;
        weights1[36228] <= 16'b0000000000101001;
        weights1[36229] <= 16'b0000000000100010;
        weights1[36230] <= 16'b0000000000010111;
        weights1[36231] <= 16'b0000000000101110;
        weights1[36232] <= 16'b1111111111111010;
        weights1[36233] <= 16'b1111111111110101;
        weights1[36234] <= 16'b1111111111111000;
        weights1[36235] <= 16'b1111111111111010;
        weights1[36236] <= 16'b1111111111100010;
        weights1[36237] <= 16'b1111111111101010;
        weights1[36238] <= 16'b1111111111101111;
        weights1[36239] <= 16'b0000000000010110;
        weights1[36240] <= 16'b1111111111110111;
        weights1[36241] <= 16'b0000000000000011;
        weights1[36242] <= 16'b1111111111110101;
        weights1[36243] <= 16'b0000000000000100;
        weights1[36244] <= 16'b0000000000001011;
        weights1[36245] <= 16'b1111111111111111;
        weights1[36246] <= 16'b0000000000010000;
        weights1[36247] <= 16'b0000000000000100;
        weights1[36248] <= 16'b1111111111110111;
        weights1[36249] <= 16'b0000000000000101;
        weights1[36250] <= 16'b0000000000000110;
        weights1[36251] <= 16'b0000000000100110;
        weights1[36252] <= 16'b0000000000100111;
        weights1[36253] <= 16'b0000000000011100;
        weights1[36254] <= 16'b0000000000011000;
        weights1[36255] <= 16'b0000000000101100;
        weights1[36256] <= 16'b0000000001011110;
        weights1[36257] <= 16'b0000000000101110;
        weights1[36258] <= 16'b0000000000101110;
        weights1[36259] <= 16'b0000000000100100;
        weights1[36260] <= 16'b1111111111111100;
        weights1[36261] <= 16'b1111111111110111;
        weights1[36262] <= 16'b1111111111101000;
        weights1[36263] <= 16'b0000000000000010;
        weights1[36264] <= 16'b1111111111110011;
        weights1[36265] <= 16'b1111111111111110;
        weights1[36266] <= 16'b0000000000000100;
        weights1[36267] <= 16'b0000000000001101;
        weights1[36268] <= 16'b1111111111110011;
        weights1[36269] <= 16'b1111111111110101;
        weights1[36270] <= 16'b0000000000001100;
        weights1[36271] <= 16'b1111111111111110;
        weights1[36272] <= 16'b0000000000001100;
        weights1[36273] <= 16'b0000000000000100;
        weights1[36274] <= 16'b0000000000011101;
        weights1[36275] <= 16'b0000000000010011;
        weights1[36276] <= 16'b0000000000101000;
        weights1[36277] <= 16'b0000000000110010;
        weights1[36278] <= 16'b0000000000110111;
        weights1[36279] <= 16'b0000000000111111;
        weights1[36280] <= 16'b0000000001010101;
        weights1[36281] <= 16'b0000000001001000;
        weights1[36282] <= 16'b0000000001000011;
        weights1[36283] <= 16'b0000000001101010;
        weights1[36284] <= 16'b0000000001010011;
        weights1[36285] <= 16'b0000000000100101;
        weights1[36286] <= 16'b0000000000011000;
        weights1[36287] <= 16'b1111111111111011;
        weights1[36288] <= 16'b1111111111111101;
        weights1[36289] <= 16'b1111111111110000;
        weights1[36290] <= 16'b1111111111110011;
        weights1[36291] <= 16'b0000000000000101;
        weights1[36292] <= 16'b1111111111100010;
        weights1[36293] <= 16'b1111111111111010;
        weights1[36294] <= 16'b1111111111110111;
        weights1[36295] <= 16'b1111111111111100;
        weights1[36296] <= 16'b1111111111110111;
        weights1[36297] <= 16'b0000000000000001;
        weights1[36298] <= 16'b1111111111111110;
        weights1[36299] <= 16'b0000000000010000;
        weights1[36300] <= 16'b0000000000001111;
        weights1[36301] <= 16'b0000000000010100;
        weights1[36302] <= 16'b0000000000011000;
        weights1[36303] <= 16'b0000000000001111;
        weights1[36304] <= 16'b0000000000101010;
        weights1[36305] <= 16'b0000000000101000;
        weights1[36306] <= 16'b0000000000100110;
        weights1[36307] <= 16'b0000000000110000;
        weights1[36308] <= 16'b0000000001000100;
        weights1[36309] <= 16'b0000000000110000;
        weights1[36310] <= 16'b0000000000010111;
        weights1[36311] <= 16'b0000000001000010;
        weights1[36312] <= 16'b0000000000010101;
        weights1[36313] <= 16'b1111111111001011;
        weights1[36314] <= 16'b1111111111001000;
        weights1[36315] <= 16'b1111111111000101;
        weights1[36316] <= 16'b1111111111110100;
        weights1[36317] <= 16'b1111111111111001;
        weights1[36318] <= 16'b0000000000001100;
        weights1[36319] <= 16'b1111111111111100;
        weights1[36320] <= 16'b1111111111111011;
        weights1[36321] <= 16'b1111111111101000;
        weights1[36322] <= 16'b1111111111111100;
        weights1[36323] <= 16'b1111111111110100;
        weights1[36324] <= 16'b0000000000000001;
        weights1[36325] <= 16'b1111111111111101;
        weights1[36326] <= 16'b0000000000000011;
        weights1[36327] <= 16'b1111111111110100;
        weights1[36328] <= 16'b1111111111110110;
        weights1[36329] <= 16'b1111111111101111;
        weights1[36330] <= 16'b1111111111011111;
        weights1[36331] <= 16'b1111111111010011;
        weights1[36332] <= 16'b1111111110111010;
        weights1[36333] <= 16'b1111111111000001;
        weights1[36334] <= 16'b1111111110101000;
        weights1[36335] <= 16'b1111111110100000;
        weights1[36336] <= 16'b1111111110000010;
        weights1[36337] <= 16'b1111111110000111;
        weights1[36338] <= 16'b1111111110010000;
        weights1[36339] <= 16'b1111111101101010;
        weights1[36340] <= 16'b1111111101110010;
        weights1[36341] <= 16'b1111111110101000;
        weights1[36342] <= 16'b1111111110100010;
        weights1[36343] <= 16'b1111111110100000;
        weights1[36344] <= 16'b1111111111110110;
        weights1[36345] <= 16'b1111111111110101;
        weights1[36346] <= 16'b0000000000000010;
        weights1[36347] <= 16'b1111111111111011;
        weights1[36348] <= 16'b1111111111111001;
        weights1[36349] <= 16'b1111111111101111;
        weights1[36350] <= 16'b1111111111111000;
        weights1[36351] <= 16'b0000000000000101;
        weights1[36352] <= 16'b1111111111101110;
        weights1[36353] <= 16'b1111111111111111;
        weights1[36354] <= 16'b1111111111110011;
        weights1[36355] <= 16'b1111111111110101;
        weights1[36356] <= 16'b1111111111001011;
        weights1[36357] <= 16'b1111111111001110;
        weights1[36358] <= 16'b1111111110110101;
        weights1[36359] <= 16'b1111111110100010;
        weights1[36360] <= 16'b1111111101110110;
        weights1[36361] <= 16'b1111111100011100;
        weights1[36362] <= 16'b1111111011101101;
        weights1[36363] <= 16'b1111111011001111;
        weights1[36364] <= 16'b1111111100000011;
        weights1[36365] <= 16'b1111111100100001;
        weights1[36366] <= 16'b1111111100110011;
        weights1[36367] <= 16'b1111111101010100;
        weights1[36368] <= 16'b1111111101001000;
        weights1[36369] <= 16'b1111111110000001;
        weights1[36370] <= 16'b1111111110011001;
        weights1[36371] <= 16'b1111111110010100;
        weights1[36372] <= 16'b1111111111111010;
        weights1[36373] <= 16'b0000000000000001;
        weights1[36374] <= 16'b1111111111111000;
        weights1[36375] <= 16'b1111111111110110;
        weights1[36376] <= 16'b0000000000001110;
        weights1[36377] <= 16'b0000000000000001;
        weights1[36378] <= 16'b0000000000001000;
        weights1[36379] <= 16'b0000000000001100;
        weights1[36380] <= 16'b1111111111101111;
        weights1[36381] <= 16'b1111111111101001;
        weights1[36382] <= 16'b1111111111110000;
        weights1[36383] <= 16'b1111111111101011;
        weights1[36384] <= 16'b1111111111110101;
        weights1[36385] <= 16'b1111111111011011;
        weights1[36386] <= 16'b1111111111110000;
        weights1[36387] <= 16'b1111111111110101;
        weights1[36388] <= 16'b1111111111101110;
        weights1[36389] <= 16'b1111111111101001;
        weights1[36390] <= 16'b1111111111000110;
        weights1[36391] <= 16'b1111111110000101;
        weights1[36392] <= 16'b1111111100110110;
        weights1[36393] <= 16'b1111111100100000;
        weights1[36394] <= 16'b1111111100110011;
        weights1[36395] <= 16'b1111111101000010;
        weights1[36396] <= 16'b1111111101010100;
        weights1[36397] <= 16'b1111111101111100;
        weights1[36398] <= 16'b1111111110101000;
        weights1[36399] <= 16'b1111111110011011;
        weights1[36400] <= 16'b0000000000000010;
        weights1[36401] <= 16'b1111111111111001;
        weights1[36402] <= 16'b1111111111111110;
        weights1[36403] <= 16'b0000000000000101;
        weights1[36404] <= 16'b1111111111110000;
        weights1[36405] <= 16'b0000000000000001;
        weights1[36406] <= 16'b1111111111101110;
        weights1[36407] <= 16'b1111111111110011;
        weights1[36408] <= 16'b0000000000010000;
        weights1[36409] <= 16'b1111111111110101;
        weights1[36410] <= 16'b1111111111110110;
        weights1[36411] <= 16'b1111111111111101;
        weights1[36412] <= 16'b0000000000000100;
        weights1[36413] <= 16'b0000000000000011;
        weights1[36414] <= 16'b0000000000000010;
        weights1[36415] <= 16'b1111111111111101;
        weights1[36416] <= 16'b0000000000010011;
        weights1[36417] <= 16'b0000000000010110;
        weights1[36418] <= 16'b0000000000010000;
        weights1[36419] <= 16'b1111111111111111;
        weights1[36420] <= 16'b1111111111100001;
        weights1[36421] <= 16'b1111111110110000;
        weights1[36422] <= 16'b1111111101111110;
        weights1[36423] <= 16'b1111111101111011;
        weights1[36424] <= 16'b1111111101101100;
        weights1[36425] <= 16'b1111111101111011;
        weights1[36426] <= 16'b1111111110011111;
        weights1[36427] <= 16'b1111111110010110;
        weights1[36428] <= 16'b1111111111111111;
        weights1[36429] <= 16'b0000000000000000;
        weights1[36430] <= 16'b0000000000001010;
        weights1[36431] <= 16'b1111111111111000;
        weights1[36432] <= 16'b0000000000000110;
        weights1[36433] <= 16'b1111111111110101;
        weights1[36434] <= 16'b0000000000010010;
        weights1[36435] <= 16'b1111111111111010;
        weights1[36436] <= 16'b1111111111101101;
        weights1[36437] <= 16'b1111111111110111;
        weights1[36438] <= 16'b0000000000000010;
        weights1[36439] <= 16'b0000000000000000;
        weights1[36440] <= 16'b0000000000001100;
        weights1[36441] <= 16'b0000000000000010;
        weights1[36442] <= 16'b1111111111111100;
        weights1[36443] <= 16'b0000000000000110;
        weights1[36444] <= 16'b1111111111110001;
        weights1[36445] <= 16'b0000000000010100;
        weights1[36446] <= 16'b1111111111111100;
        weights1[36447] <= 16'b0000000000001111;
        weights1[36448] <= 16'b0000000000010100;
        weights1[36449] <= 16'b0000000000000101;
        weights1[36450] <= 16'b0000000000010101;
        weights1[36451] <= 16'b1111111111010001;
        weights1[36452] <= 16'b1111111111011000;
        weights1[36453] <= 16'b1111111110111001;
        weights1[36454] <= 16'b1111111110100111;
        weights1[36455] <= 16'b1111111110100101;
        weights1[36456] <= 16'b1111111111110111;
        weights1[36457] <= 16'b0000000000000111;
        weights1[36458] <= 16'b0000000000010000;
        weights1[36459] <= 16'b0000000000000010;
        weights1[36460] <= 16'b0000000000010001;
        weights1[36461] <= 16'b1111111111101001;
        weights1[36462] <= 16'b0000000000011001;
        weights1[36463] <= 16'b0000000000010000;
        weights1[36464] <= 16'b0000000000010011;
        weights1[36465] <= 16'b1111111111111111;
        weights1[36466] <= 16'b0000000000000001;
        weights1[36467] <= 16'b0000000000001110;
        weights1[36468] <= 16'b1111111111111101;
        weights1[36469] <= 16'b0000000000001010;
        weights1[36470] <= 16'b1111111111111111;
        weights1[36471] <= 16'b0000000000001010;
        weights1[36472] <= 16'b0000000000001001;
        weights1[36473] <= 16'b1111111111111010;
        weights1[36474] <= 16'b0000000000010000;
        weights1[36475] <= 16'b0000000000010001;
        weights1[36476] <= 16'b0000000000100000;
        weights1[36477] <= 16'b0000000000010001;
        weights1[36478] <= 16'b0000000000011101;
        weights1[36479] <= 16'b0000000000100100;
        weights1[36480] <= 16'b0000000000100010;
        weights1[36481] <= 16'b1111111111110110;
        weights1[36482] <= 16'b1111111111100000;
        weights1[36483] <= 16'b1111111111010011;
        weights1[36484] <= 16'b1111111111111101;
        weights1[36485] <= 16'b0000000000001011;
        weights1[36486] <= 16'b0000000000000010;
        weights1[36487] <= 16'b0000000000000010;
        weights1[36488] <= 16'b0000000000010110;
        weights1[36489] <= 16'b0000000000001101;
        weights1[36490] <= 16'b0000000000000101;
        weights1[36491] <= 16'b1111111111110100;
        weights1[36492] <= 16'b0000000000010100;
        weights1[36493] <= 16'b1111111111111011;
        weights1[36494] <= 16'b0000000000001111;
        weights1[36495] <= 16'b0000000000000001;
        weights1[36496] <= 16'b1111111111110100;
        weights1[36497] <= 16'b1111111111111111;
        weights1[36498] <= 16'b1111111111101011;
        weights1[36499] <= 16'b0000000000001001;
        weights1[36500] <= 16'b0000000000000111;
        weights1[36501] <= 16'b0000000000000111;
        weights1[36502] <= 16'b0000000000001001;
        weights1[36503] <= 16'b0000000000000000;
        weights1[36504] <= 16'b0000000000011010;
        weights1[36505] <= 16'b0000000000010101;
        weights1[36506] <= 16'b0000000000000001;
        weights1[36507] <= 16'b0000000000101001;
        weights1[36508] <= 16'b0000000000011011;
        weights1[36509] <= 16'b0000000000000110;
        weights1[36510] <= 16'b0000000000000001;
        weights1[36511] <= 16'b1111111111110110;
        weights1[36512] <= 16'b1111111111111110;
        weights1[36513] <= 16'b0000000000010000;
        weights1[36514] <= 16'b0000000000001111;
        weights1[36515] <= 16'b1111111111111010;
        weights1[36516] <= 16'b0000000000000001;
        weights1[36517] <= 16'b1111111111111100;
        weights1[36518] <= 16'b1111111111111101;
        weights1[36519] <= 16'b0000000000001010;
        weights1[36520] <= 16'b1111111111111010;
        weights1[36521] <= 16'b0000000000001001;
        weights1[36522] <= 16'b0000000000000011;
        weights1[36523] <= 16'b0000000000000100;
        weights1[36524] <= 16'b1111111111111100;
        weights1[36525] <= 16'b0000000000000110;
        weights1[36526] <= 16'b0000000000001100;
        weights1[36527] <= 16'b0000000000000101;
        weights1[36528] <= 16'b1111111111111110;
        weights1[36529] <= 16'b0000000000010110;
        weights1[36530] <= 16'b0000000000000001;
        weights1[36531] <= 16'b0000000000000101;
        weights1[36532] <= 16'b1111111111111110;
        weights1[36533] <= 16'b0000000000001011;
        weights1[36534] <= 16'b0000000000100000;
        weights1[36535] <= 16'b0000000000001010;
        weights1[36536] <= 16'b0000000000010001;
        weights1[36537] <= 16'b1111111111111011;
        weights1[36538] <= 16'b0000000000000110;
        weights1[36539] <= 16'b0000000000000100;
        weights1[36540] <= 16'b0000000000000100;
        weights1[36541] <= 16'b1111111111111100;
        weights1[36542] <= 16'b1111111111111010;
        weights1[36543] <= 16'b1111111111111110;
        weights1[36544] <= 16'b1111111111110011;
        weights1[36545] <= 16'b0000000000001101;
        weights1[36546] <= 16'b1111111111111010;
        weights1[36547] <= 16'b0000000000000011;
        weights1[36548] <= 16'b0000000000010100;
        weights1[36549] <= 16'b1111111111110011;
        weights1[36550] <= 16'b0000000000000100;
        weights1[36551] <= 16'b0000000000000111;
        weights1[36552] <= 16'b1111111111111010;
        weights1[36553] <= 16'b0000000000000000;
        weights1[36554] <= 16'b1111111111110010;
        weights1[36555] <= 16'b1111111111111000;
        weights1[36556] <= 16'b1111111111111011;
        weights1[36557] <= 16'b1111111111111010;
        weights1[36558] <= 16'b0000000000010100;
        weights1[36559] <= 16'b0000000000000011;
        weights1[36560] <= 16'b0000000000001110;
        weights1[36561] <= 16'b1111111111101110;
        weights1[36562] <= 16'b1111111111111111;
        weights1[36563] <= 16'b0000000000000101;
        weights1[36564] <= 16'b0000000000010010;
        weights1[36565] <= 16'b1111111111111101;
        weights1[36566] <= 16'b0000000000010000;
        weights1[36567] <= 16'b1111111111110101;
        weights1[36568] <= 16'b1111111111111111;
        weights1[36569] <= 16'b1111111111110101;
        weights1[36570] <= 16'b1111111111111101;
        weights1[36571] <= 16'b0000000000010010;
        weights1[36572] <= 16'b0000000000000100;
        weights1[36573] <= 16'b1111111111111111;
        weights1[36574] <= 16'b0000000000000001;
        weights1[36575] <= 16'b0000000000000011;
        weights1[36576] <= 16'b1111111111110111;
        weights1[36577] <= 16'b0000000000000110;
        weights1[36578] <= 16'b0000000000000000;
        weights1[36579] <= 16'b1111111111111000;
        weights1[36580] <= 16'b0000000000001001;
        weights1[36581] <= 16'b0000000000001110;
        weights1[36582] <= 16'b1111111111110100;
        weights1[36583] <= 16'b0000000000000111;
        weights1[36584] <= 16'b0000000000001010;
        weights1[36585] <= 16'b1111111111111111;
        weights1[36586] <= 16'b1111111111111100;
        weights1[36587] <= 16'b0000000000011001;
        weights1[36588] <= 16'b0000000000000101;
        weights1[36589] <= 16'b1111111111111101;
        weights1[36590] <= 16'b0000000000000110;
        weights1[36591] <= 16'b0000000000001010;
        weights1[36592] <= 16'b1111111111111000;
        weights1[36593] <= 16'b0000000000000110;
        weights1[36594] <= 16'b0000000000000011;
        weights1[36595] <= 16'b1111111111111000;
        weights1[36596] <= 16'b1111111111111000;
        weights1[36597] <= 16'b0000000000000011;
        weights1[36598] <= 16'b0000000000000100;
        weights1[36599] <= 16'b1111111111110000;
        weights1[36600] <= 16'b0000000000000110;
        weights1[36601] <= 16'b0000000000001100;
        weights1[36602] <= 16'b1111111111111001;
        weights1[36603] <= 16'b1111111111101100;
        weights1[36604] <= 16'b0000000000010001;
        weights1[36605] <= 16'b0000000000000001;
        weights1[36606] <= 16'b0000000000000000;
        weights1[36607] <= 16'b1111111111110101;
        weights1[36608] <= 16'b0000000000011100;
        weights1[36609] <= 16'b1111111111110110;
        weights1[36610] <= 16'b0000000000010010;
        weights1[36611] <= 16'b0000000000000100;
        weights1[36612] <= 16'b0000000000000011;
        weights1[36613] <= 16'b0000000000001000;
        weights1[36614] <= 16'b0000000000000110;
        weights1[36615] <= 16'b0000000000000000;
        weights1[36616] <= 16'b1111111111111110;
        weights1[36617] <= 16'b0000000000000110;
        weights1[36618] <= 16'b0000000000010011;
        weights1[36619] <= 16'b1111111111101111;
        weights1[36620] <= 16'b0000000000011010;
        weights1[36621] <= 16'b0000000000000110;
        weights1[36622] <= 16'b0000000000001011;
        weights1[36623] <= 16'b0000000000010000;
        weights1[36624] <= 16'b1111111111111111;
        weights1[36625] <= 16'b1111111111111011;
        weights1[36626] <= 16'b1111111111111110;
        weights1[36627] <= 16'b1111111111111101;
        weights1[36628] <= 16'b1111111111110001;
        weights1[36629] <= 16'b0000000000000101;
        weights1[36630] <= 16'b0000000000000001;
        weights1[36631] <= 16'b1111111111101011;
        weights1[36632] <= 16'b1111111111111010;
        weights1[36633] <= 16'b0000000000000010;
        weights1[36634] <= 16'b1111111111111001;
        weights1[36635] <= 16'b0000000000010100;
        weights1[36636] <= 16'b1111111111111111;
        weights1[36637] <= 16'b1111111111110011;
        weights1[36638] <= 16'b1111111111111111;
        weights1[36639] <= 16'b0000000000001000;
        weights1[36640] <= 16'b1111111111111111;
        weights1[36641] <= 16'b0000000000001010;
        weights1[36642] <= 16'b1111111111111100;
        weights1[36643] <= 16'b1111111111101011;
        weights1[36644] <= 16'b0000000000001000;
        weights1[36645] <= 16'b0000000000001110;
        weights1[36646] <= 16'b0000000000000011;
        weights1[36647] <= 16'b0000000000010001;
        weights1[36648] <= 16'b1111111111110111;
        weights1[36649] <= 16'b0000000000010000;
        weights1[36650] <= 16'b0000000000001011;
        weights1[36651] <= 16'b0000000000001110;
        weights1[36652] <= 16'b1111111111111111;
        weights1[36653] <= 16'b0000000000001001;
        weights1[36654] <= 16'b0000000000001111;
        weights1[36655] <= 16'b0000000000010011;
        weights1[36656] <= 16'b0000000000010001;
        weights1[36657] <= 16'b0000000000010001;
        weights1[36658] <= 16'b1111111111111100;
        weights1[36659] <= 16'b0000000000010111;
        weights1[36660] <= 16'b1111111111110010;
        weights1[36661] <= 16'b0000000000001010;
        weights1[36662] <= 16'b0000000000001101;
        weights1[36663] <= 16'b0000000000000000;
        weights1[36664] <= 16'b0000000000000110;
        weights1[36665] <= 16'b0000000000010111;
        weights1[36666] <= 16'b1111111111111010;
        weights1[36667] <= 16'b0000000000001110;
        weights1[36668] <= 16'b0000000000001101;
        weights1[36669] <= 16'b0000000000010000;
        weights1[36670] <= 16'b0000000000000110;
        weights1[36671] <= 16'b0000000000001111;
        weights1[36672] <= 16'b1111111111111100;
        weights1[36673] <= 16'b1111111111110100;
        weights1[36674] <= 16'b0000000000011010;
        weights1[36675] <= 16'b0000000000011101;
        weights1[36676] <= 16'b0000000000000001;
        weights1[36677] <= 16'b0000000000011110;
        weights1[36678] <= 16'b0000000000000000;
        weights1[36679] <= 16'b0000000000000010;
        weights1[36680] <= 16'b1111111111110100;
        weights1[36681] <= 16'b1111111111111111;
        weights1[36682] <= 16'b0000000000001011;
        weights1[36683] <= 16'b1111111111111111;
        weights1[36684] <= 16'b1111111111111001;
        weights1[36685] <= 16'b1111111111111001;
        weights1[36686] <= 16'b1111111111111110;
        weights1[36687] <= 16'b1111111111111110;
        weights1[36688] <= 16'b0000000000001001;
        weights1[36689] <= 16'b1111111111101101;
        weights1[36690] <= 16'b0000000000010000;
        weights1[36691] <= 16'b1111111111110000;
        weights1[36692] <= 16'b0000000000001100;
        weights1[36693] <= 16'b1111111111111100;
        weights1[36694] <= 16'b0000000000000110;
        weights1[36695] <= 16'b0000000000000100;
        weights1[36696] <= 16'b1111111111111010;
        weights1[36697] <= 16'b1111111111111110;
        weights1[36698] <= 16'b0000000000011000;
        weights1[36699] <= 16'b1111111111110110;
        weights1[36700] <= 16'b0000000000010010;
        weights1[36701] <= 16'b1111111111110010;
        weights1[36702] <= 16'b0000000000010001;
        weights1[36703] <= 16'b0000000000001101;
        weights1[36704] <= 16'b1111111111111101;
        weights1[36705] <= 16'b0000000000001011;
        weights1[36706] <= 16'b1111111111111101;
        weights1[36707] <= 16'b0000000000000111;
        weights1[36708] <= 16'b1111111111111100;
        weights1[36709] <= 16'b1111111111111010;
        weights1[36710] <= 16'b1111111111110001;
        weights1[36711] <= 16'b1111111111101111;
        weights1[36712] <= 16'b1111111111111010;
        weights1[36713] <= 16'b0000000000000011;
        weights1[36714] <= 16'b1111111111101011;
        weights1[36715] <= 16'b1111111111111100;
        weights1[36716] <= 16'b1111111111111110;
        weights1[36717] <= 16'b0000000000001111;
        weights1[36718] <= 16'b1111111111110001;
        weights1[36719] <= 16'b1111111111101101;
        weights1[36720] <= 16'b1111111111111100;
        weights1[36721] <= 16'b1111111111110101;
        weights1[36722] <= 16'b0000000000001000;
        weights1[36723] <= 16'b0000000000000110;
        weights1[36724] <= 16'b0000000000001010;
        weights1[36725] <= 16'b1111111111111010;
        weights1[36726] <= 16'b1111111111111110;
        weights1[36727] <= 16'b0000000000001101;
        weights1[36728] <= 16'b0000000000001010;
        weights1[36729] <= 16'b0000000000000011;
        weights1[36730] <= 16'b1111111111111111;
        weights1[36731] <= 16'b0000000000001101;
        weights1[36732] <= 16'b0000000000001101;
        weights1[36733] <= 16'b0000000000000010;
        weights1[36734] <= 16'b0000000000000110;
        weights1[36735] <= 16'b1111111111111100;
        weights1[36736] <= 16'b1111111111111010;
        weights1[36737] <= 16'b0000000000000001;
        weights1[36738] <= 16'b1111111111111010;
        weights1[36739] <= 16'b0000000000000010;
        weights1[36740] <= 16'b1111111111111010;
        weights1[36741] <= 16'b0000000000010100;
        weights1[36742] <= 16'b0000000000000000;
        weights1[36743] <= 16'b0000000000001010;
        weights1[36744] <= 16'b1111111111101011;
        weights1[36745] <= 16'b0000000000001110;
        weights1[36746] <= 16'b1111111111111000;
        weights1[36747] <= 16'b0000000000000111;
        weights1[36748] <= 16'b0000000000000100;
        weights1[36749] <= 16'b1111111111110000;
        weights1[36750] <= 16'b1111111111111010;
        weights1[36751] <= 16'b0000000000000101;
        weights1[36752] <= 16'b1111111111110001;
        weights1[36753] <= 16'b0000000000000101;
        weights1[36754] <= 16'b1111111111111100;
        weights1[36755] <= 16'b1111111111110000;
        weights1[36756] <= 16'b0000000000001010;
        weights1[36757] <= 16'b0000000000000000;
        weights1[36758] <= 16'b1111111111111111;
        weights1[36759] <= 16'b0000000000000110;
        weights1[36760] <= 16'b0000000000000111;
        weights1[36761] <= 16'b1111111111111000;
        weights1[36762] <= 16'b1111111111111101;
        weights1[36763] <= 16'b1111111111111100;
        weights1[36764] <= 16'b1111111111111011;
        weights1[36765] <= 16'b0000000000000000;
        weights1[36766] <= 16'b1111111111111111;
        weights1[36767] <= 16'b0000000000000101;
        weights1[36768] <= 16'b1111111111111111;
        weights1[36769] <= 16'b0000000000000100;
        weights1[36770] <= 16'b0000000000000010;
        weights1[36771] <= 16'b0000000000000011;
        weights1[36772] <= 16'b1111111111111001;
        weights1[36773] <= 16'b0000000000010100;
        weights1[36774] <= 16'b1111111111110111;
        weights1[36775] <= 16'b1111111111110000;
        weights1[36776] <= 16'b0000000000010100;
        weights1[36777] <= 16'b0000000000000000;
        weights1[36778] <= 16'b0000000000001011;
        weights1[36779] <= 16'b0000000000001110;
        weights1[36780] <= 16'b0000000000000101;
        weights1[36781] <= 16'b0000000000010001;
        weights1[36782] <= 16'b0000000000001100;
        weights1[36783] <= 16'b1111111111111000;
        weights1[36784] <= 16'b0000000000011001;
        weights1[36785] <= 16'b0000000000000111;
        weights1[36786] <= 16'b0000000000001111;
        weights1[36787] <= 16'b0000000000001011;
        weights1[36788] <= 16'b0000000000000000;
        weights1[36789] <= 16'b1111111111111100;
        weights1[36790] <= 16'b1111111111110111;
        weights1[36791] <= 16'b1111111111111011;
        weights1[36792] <= 16'b1111111111111111;
        weights1[36793] <= 16'b1111111111111110;
        weights1[36794] <= 16'b1111111111111101;
        weights1[36795] <= 16'b1111111111111000;
        weights1[36796] <= 16'b1111111111110111;
        weights1[36797] <= 16'b1111111111100111;
        weights1[36798] <= 16'b1111111111101010;
        weights1[36799] <= 16'b1111111111111001;
        weights1[36800] <= 16'b0000000000000011;
        weights1[36801] <= 16'b0000000000000001;
        weights1[36802] <= 16'b1111111111111111;
        weights1[36803] <= 16'b0000000000000111;
        weights1[36804] <= 16'b1111111111110111;
        weights1[36805] <= 16'b0000000000000011;
        weights1[36806] <= 16'b1111111111110010;
        weights1[36807] <= 16'b1111111111110000;
        weights1[36808] <= 16'b1111111111111010;
        weights1[36809] <= 16'b1111111111111010;
        weights1[36810] <= 16'b0000000000001010;
        weights1[36811] <= 16'b0000000000001000;
        weights1[36812] <= 16'b1111111111111010;
        weights1[36813] <= 16'b1111111111110010;
        weights1[36814] <= 16'b1111111111111010;
        weights1[36815] <= 16'b1111111111111010;
        weights1[36816] <= 16'b0000000000001000;
        weights1[36817] <= 16'b0000000000000001;
        weights1[36818] <= 16'b0000000000000001;
        weights1[36819] <= 16'b0000000000000000;
        weights1[36820] <= 16'b1111111111111111;
        weights1[36821] <= 16'b1111111111111101;
        weights1[36822] <= 16'b1111111111111101;
        weights1[36823] <= 16'b1111111111111010;
        weights1[36824] <= 16'b1111111111111110;
        weights1[36825] <= 16'b0000000000000001;
        weights1[36826] <= 16'b1111111111111100;
        weights1[36827] <= 16'b1111111111110010;
        weights1[36828] <= 16'b1111111111101100;
        weights1[36829] <= 16'b0000000000000000;
        weights1[36830] <= 16'b1111111111101001;
        weights1[36831] <= 16'b1111111111111011;
        weights1[36832] <= 16'b1111111111110100;
        weights1[36833] <= 16'b1111111111101110;
        weights1[36834] <= 16'b1111111111110100;
        weights1[36835] <= 16'b0000000000000101;
        weights1[36836] <= 16'b1111111111111011;
        weights1[36837] <= 16'b1111111111111001;
        weights1[36838] <= 16'b1111111111101001;
        weights1[36839] <= 16'b1111111111101100;
        weights1[36840] <= 16'b1111111111111010;
        weights1[36841] <= 16'b1111111111100010;
        weights1[36842] <= 16'b1111111111111000;
        weights1[36843] <= 16'b0000000000000110;
        weights1[36844] <= 16'b0000000000000110;
        weights1[36845] <= 16'b0000000000000000;
        weights1[36846] <= 16'b0000000000000010;
        weights1[36847] <= 16'b0000000000000000;
        weights1[36848] <= 16'b0000000000000000;
        weights1[36849] <= 16'b0000000000000000;
        weights1[36850] <= 16'b0000000000000011;
        weights1[36851] <= 16'b0000000000000100;
        weights1[36852] <= 16'b0000000000001001;
        weights1[36853] <= 16'b0000000000001110;
        weights1[36854] <= 16'b0000000000001101;
        weights1[36855] <= 16'b0000000000001111;
        weights1[36856] <= 16'b0000000000011000;
        weights1[36857] <= 16'b0000000000100000;
        weights1[36858] <= 16'b0000000000100001;
        weights1[36859] <= 16'b0000000000010111;
        weights1[36860] <= 16'b0000000000000001;
        weights1[36861] <= 16'b0000000000001110;
        weights1[36862] <= 16'b0000000000010011;
        weights1[36863] <= 16'b0000000000010000;
        weights1[36864] <= 16'b0000000000010110;
        weights1[36865] <= 16'b0000000000000100;
        weights1[36866] <= 16'b0000000000000100;
        weights1[36867] <= 16'b1111111111111100;
        weights1[36868] <= 16'b0000000000000000;
        weights1[36869] <= 16'b0000000000001001;
        weights1[36870] <= 16'b0000000000000001;
        weights1[36871] <= 16'b1111111111111010;
        weights1[36872] <= 16'b0000000000000001;
        weights1[36873] <= 16'b0000000000001111;
        weights1[36874] <= 16'b0000000000000111;
        weights1[36875] <= 16'b1111111111111100;
        weights1[36876] <= 16'b0000000000000000;
        weights1[36877] <= 16'b0000000000000011;
        weights1[36878] <= 16'b0000000000001000;
        weights1[36879] <= 16'b0000000000001010;
        weights1[36880] <= 16'b0000000000011011;
        weights1[36881] <= 16'b0000000000011101;
        weights1[36882] <= 16'b0000000000100000;
        weights1[36883] <= 16'b0000000000100010;
        weights1[36884] <= 16'b0000000000011011;
        weights1[36885] <= 16'b0000000000001101;
        weights1[36886] <= 16'b0000000000011100;
        weights1[36887] <= 16'b0000000000000010;
        weights1[36888] <= 16'b0000000000000101;
        weights1[36889] <= 16'b0000000000001000;
        weights1[36890] <= 16'b1111111111111001;
        weights1[36891] <= 16'b1111111111111100;
        weights1[36892] <= 16'b0000000000001001;
        weights1[36893] <= 16'b0000000000000100;
        weights1[36894] <= 16'b0000000000000101;
        weights1[36895] <= 16'b1111111111110011;
        weights1[36896] <= 16'b1111111111111111;
        weights1[36897] <= 16'b1111111111110010;
        weights1[36898] <= 16'b1111111111111010;
        weights1[36899] <= 16'b1111111111110100;
        weights1[36900] <= 16'b0000000000000110;
        weights1[36901] <= 16'b0000000000001010;
        weights1[36902] <= 16'b0000000000010010;
        weights1[36903] <= 16'b0000000000000011;
        weights1[36904] <= 16'b0000000000000010;
        weights1[36905] <= 16'b0000000000001000;
        weights1[36906] <= 16'b0000000000000001;
        weights1[36907] <= 16'b0000000000010000;
        weights1[36908] <= 16'b0000000000011010;
        weights1[36909] <= 16'b0000000000010100;
        weights1[36910] <= 16'b0000000000010101;
        weights1[36911] <= 16'b0000000000100011;
        weights1[36912] <= 16'b0000000000010000;
        weights1[36913] <= 16'b0000000000011110;
        weights1[36914] <= 16'b0000000000001011;
        weights1[36915] <= 16'b0000000000001111;
        weights1[36916] <= 16'b0000000000010000;
        weights1[36917] <= 16'b0000000000011010;
        weights1[36918] <= 16'b0000000000000011;
        weights1[36919] <= 16'b0000000000000101;
        weights1[36920] <= 16'b1111111111111111;
        weights1[36921] <= 16'b0000000000000101;
        weights1[36922] <= 16'b0000000000000010;
        weights1[36923] <= 16'b1111111111111010;
        weights1[36924] <= 16'b1111111111111101;
        weights1[36925] <= 16'b0000000000000101;
        weights1[36926] <= 16'b0000000000000010;
        weights1[36927] <= 16'b1111111111111111;
        weights1[36928] <= 16'b0000000000000010;
        weights1[36929] <= 16'b1111111111111100;
        weights1[36930] <= 16'b0000000000000000;
        weights1[36931] <= 16'b1111111111111101;
        weights1[36932] <= 16'b0000000000000011;
        weights1[36933] <= 16'b0000000000001010;
        weights1[36934] <= 16'b0000000000000001;
        weights1[36935] <= 16'b0000000000010000;
        weights1[36936] <= 16'b0000000000001111;
        weights1[36937] <= 16'b0000000000010011;
        weights1[36938] <= 16'b0000000000010001;
        weights1[36939] <= 16'b0000000000011100;
        weights1[36940] <= 16'b0000000000001111;
        weights1[36941] <= 16'b0000000000000111;
        weights1[36942] <= 16'b0000000000001100;
        weights1[36943] <= 16'b0000000000000111;
        weights1[36944] <= 16'b0000000000001110;
        weights1[36945] <= 16'b0000000000000111;
        weights1[36946] <= 16'b1111111111111011;
        weights1[36947] <= 16'b0000000000011000;
        weights1[36948] <= 16'b0000000000001100;
        weights1[36949] <= 16'b1111111111110110;
        weights1[36950] <= 16'b0000000000000110;
        weights1[36951] <= 16'b0000000000001100;
        weights1[36952] <= 16'b0000000000001010;
        weights1[36953] <= 16'b0000000000000001;
        weights1[36954] <= 16'b0000000000000001;
        weights1[36955] <= 16'b1111111111110100;
        weights1[36956] <= 16'b0000000000000000;
        weights1[36957] <= 16'b1111111111111001;
        weights1[36958] <= 16'b0000000000001011;
        weights1[36959] <= 16'b0000000000001100;
        weights1[36960] <= 16'b0000000000000110;
        weights1[36961] <= 16'b0000000000000111;
        weights1[36962] <= 16'b0000000000000111;
        weights1[36963] <= 16'b1111111111111001;
        weights1[36964] <= 16'b1111111111110010;
        weights1[36965] <= 16'b0000000000000010;
        weights1[36966] <= 16'b0000000000001000;
        weights1[36967] <= 16'b0000000000010011;
        weights1[36968] <= 16'b0000000000001010;
        weights1[36969] <= 16'b0000000000010101;
        weights1[36970] <= 16'b0000000000011000;
        weights1[36971] <= 16'b0000000000110000;
        weights1[36972] <= 16'b0000000000001100;
        weights1[36973] <= 16'b0000000000010011;
        weights1[36974] <= 16'b0000000000010100;
        weights1[36975] <= 16'b1111111111110100;
        weights1[36976] <= 16'b0000000000011010;
        weights1[36977] <= 16'b1111111111111110;
        weights1[36978] <= 16'b0000000000000101;
        weights1[36979] <= 16'b1111111111110111;
        weights1[36980] <= 16'b0000000000000011;
        weights1[36981] <= 16'b1111111111111010;
        weights1[36982] <= 16'b1111111111111101;
        weights1[36983] <= 16'b0000000000001001;
        weights1[36984] <= 16'b0000000000001001;
        weights1[36985] <= 16'b0000000000001011;
        weights1[36986] <= 16'b0000000000000011;
        weights1[36987] <= 16'b0000000000000101;
        weights1[36988] <= 16'b0000000000000101;
        weights1[36989] <= 16'b0000000000001001;
        weights1[36990] <= 16'b0000000000000001;
        weights1[36991] <= 16'b1111111111101110;
        weights1[36992] <= 16'b1111111111111011;
        weights1[36993] <= 16'b0000000000001010;
        weights1[36994] <= 16'b0000000000001010;
        weights1[36995] <= 16'b1111111111110100;
        weights1[36996] <= 16'b0000000000011011;
        weights1[36997] <= 16'b0000000000010001;
        weights1[36998] <= 16'b0000000000000110;
        weights1[36999] <= 16'b0000000000000110;
        weights1[37000] <= 16'b0000000000011000;
        weights1[37001] <= 16'b0000000000011101;
        weights1[37002] <= 16'b0000000000010010;
        weights1[37003] <= 16'b0000000000001101;
        weights1[37004] <= 16'b0000000000010011;
        weights1[37005] <= 16'b0000000000011001;
        weights1[37006] <= 16'b0000000000001100;
        weights1[37007] <= 16'b0000000000000010;
        weights1[37008] <= 16'b0000000000000110;
        weights1[37009] <= 16'b0000000000001111;
        weights1[37010] <= 16'b0000000000001101;
        weights1[37011] <= 16'b0000000000000010;
        weights1[37012] <= 16'b1111111111111000;
        weights1[37013] <= 16'b0000000000000001;
        weights1[37014] <= 16'b0000000000001001;
        weights1[37015] <= 16'b0000000000000010;
        weights1[37016] <= 16'b0000000000000101;
        weights1[37017] <= 16'b1111111111111010;
        weights1[37018] <= 16'b1111111111110010;
        weights1[37019] <= 16'b1111111111101100;
        weights1[37020] <= 16'b1111111111101000;
        weights1[37021] <= 16'b1111111111101000;
        weights1[37022] <= 16'b0000000000000000;
        weights1[37023] <= 16'b1111111111101111;
        weights1[37024] <= 16'b1111111111101100;
        weights1[37025] <= 16'b1111111111110000;
        weights1[37026] <= 16'b1111111111101100;
        weights1[37027] <= 16'b1111111111111001;
        weights1[37028] <= 16'b1111111111111011;
        weights1[37029] <= 16'b0000000000001001;
        weights1[37030] <= 16'b0000000000000011;
        weights1[37031] <= 16'b0000000000001010;
        weights1[37032] <= 16'b0000000000000011;
        weights1[37033] <= 16'b1111111111110111;
        weights1[37034] <= 16'b0000000000010001;
        weights1[37035] <= 16'b0000000000000110;
        weights1[37036] <= 16'b0000000000001010;
        weights1[37037] <= 16'b0000000000000100;
        weights1[37038] <= 16'b0000000000001010;
        weights1[37039] <= 16'b0000000000001100;
        weights1[37040] <= 16'b0000000000010001;
        weights1[37041] <= 16'b0000000000000100;
        weights1[37042] <= 16'b0000000000000001;
        weights1[37043] <= 16'b0000000000001001;
        weights1[37044] <= 16'b1111111111110101;
        weights1[37045] <= 16'b1111111111100101;
        weights1[37046] <= 16'b1111111111100100;
        weights1[37047] <= 16'b1111111111011011;
        weights1[37048] <= 16'b1111111111011101;
        weights1[37049] <= 16'b1111111111001010;
        weights1[37050] <= 16'b1111111111100000;
        weights1[37051] <= 16'b1111111111011000;
        weights1[37052] <= 16'b1111111111100011;
        weights1[37053] <= 16'b1111111111101100;
        weights1[37054] <= 16'b1111111111101011;
        weights1[37055] <= 16'b1111111111101000;
        weights1[37056] <= 16'b1111111111100111;
        weights1[37057] <= 16'b1111111111101011;
        weights1[37058] <= 16'b1111111111110101;
        weights1[37059] <= 16'b1111111111101001;
        weights1[37060] <= 16'b0000000000000010;
        weights1[37061] <= 16'b1111111111110100;
        weights1[37062] <= 16'b1111111111111100;
        weights1[37063] <= 16'b1111111111111010;
        weights1[37064] <= 16'b1111111111111110;
        weights1[37065] <= 16'b1111111111111001;
        weights1[37066] <= 16'b1111111111111011;
        weights1[37067] <= 16'b1111111111111011;
        weights1[37068] <= 16'b1111111111110111;
        weights1[37069] <= 16'b0000000000000000;
        weights1[37070] <= 16'b0000000000001110;
        weights1[37071] <= 16'b0000000000001110;
        weights1[37072] <= 16'b1111111111110001;
        weights1[37073] <= 16'b1111111111011000;
        weights1[37074] <= 16'b1111111111011011;
        weights1[37075] <= 16'b1111111111010011;
        weights1[37076] <= 16'b1111111111001111;
        weights1[37077] <= 16'b1111111111010011;
        weights1[37078] <= 16'b1111111111011001;
        weights1[37079] <= 16'b1111111111101011;
        weights1[37080] <= 16'b1111111111010101;
        weights1[37081] <= 16'b1111111111101111;
        weights1[37082] <= 16'b1111111111111110;
        weights1[37083] <= 16'b1111111111110100;
        weights1[37084] <= 16'b1111111111100001;
        weights1[37085] <= 16'b0000000000001110;
        weights1[37086] <= 16'b1111111111110001;
        weights1[37087] <= 16'b0000000000001100;
        weights1[37088] <= 16'b1111111111101011;
        weights1[37089] <= 16'b0000000000000001;
        weights1[37090] <= 16'b0000000000000010;
        weights1[37091] <= 16'b1111111111101000;
        weights1[37092] <= 16'b0000000000000100;
        weights1[37093] <= 16'b1111111111111001;
        weights1[37094] <= 16'b0000000000010010;
        weights1[37095] <= 16'b0000000000000110;
        weights1[37096] <= 16'b1111111111101110;
        weights1[37097] <= 16'b0000000000000010;
        weights1[37098] <= 16'b1111111111111001;
        weights1[37099] <= 16'b0000000000000111;
        weights1[37100] <= 16'b1111111111100110;
        weights1[37101] <= 16'b1111111111010011;
        weights1[37102] <= 16'b1111111111010110;
        weights1[37103] <= 16'b1111111111010111;
        weights1[37104] <= 16'b1111111111101100;
        weights1[37105] <= 16'b1111111111110010;
        weights1[37106] <= 16'b0000000000000010;
        weights1[37107] <= 16'b0000000000000110;
        weights1[37108] <= 16'b1111111111101110;
        weights1[37109] <= 16'b1111111111110000;
        weights1[37110] <= 16'b1111111111111110;
        weights1[37111] <= 16'b0000000000001111;
        weights1[37112] <= 16'b0000000000000101;
        weights1[37113] <= 16'b0000000000001110;
        weights1[37114] <= 16'b0000000000001010;
        weights1[37115] <= 16'b0000000000000100;
        weights1[37116] <= 16'b0000000000010001;
        weights1[37117] <= 16'b0000000000000101;
        weights1[37118] <= 16'b0000000000000110;
        weights1[37119] <= 16'b1111111111111000;
        weights1[37120] <= 16'b1111111111110100;
        weights1[37121] <= 16'b1111111111111010;
        weights1[37122] <= 16'b1111111111101101;
        weights1[37123] <= 16'b1111111111111101;
        weights1[37124] <= 16'b1111111111111010;
        weights1[37125] <= 16'b0000000000000001;
        weights1[37126] <= 16'b0000000000000011;
        weights1[37127] <= 16'b0000000000000101;
        weights1[37128] <= 16'b1111111111011110;
        weights1[37129] <= 16'b1111111111000101;
        weights1[37130] <= 16'b1111111111000101;
        weights1[37131] <= 16'b1111111111001100;
        weights1[37132] <= 16'b1111111111011111;
        weights1[37133] <= 16'b1111111111111101;
        weights1[37134] <= 16'b0000000000000000;
        weights1[37135] <= 16'b0000000000010011;
        weights1[37136] <= 16'b0000000000000110;
        weights1[37137] <= 16'b0000000000100101;
        weights1[37138] <= 16'b0000000000001111;
        weights1[37139] <= 16'b0000000000010101;
        weights1[37140] <= 16'b0000000000100101;
        weights1[37141] <= 16'b0000000000011100;
        weights1[37142] <= 16'b0000000000001101;
        weights1[37143] <= 16'b0000000000010010;
        weights1[37144] <= 16'b1111111111111100;
        weights1[37145] <= 16'b0000000000001011;
        weights1[37146] <= 16'b0000000000001000;
        weights1[37147] <= 16'b0000000000000101;
        weights1[37148] <= 16'b0000000000001001;
        weights1[37149] <= 16'b0000000000010000;
        weights1[37150] <= 16'b1111111111111110;
        weights1[37151] <= 16'b0000000000000100;
        weights1[37152] <= 16'b1111111111111110;
        weights1[37153] <= 16'b1111111111110111;
        weights1[37154] <= 16'b1111111111110011;
        weights1[37155] <= 16'b0000000000000000;
        weights1[37156] <= 16'b1111111111100000;
        weights1[37157] <= 16'b1111111111000101;
        weights1[37158] <= 16'b1111111110110100;
        weights1[37159] <= 16'b1111111110101001;
        weights1[37160] <= 16'b1111111110111010;
        weights1[37161] <= 16'b1111111111000111;
        weights1[37162] <= 16'b1111111111101001;
        weights1[37163] <= 16'b0000000000000100;
        weights1[37164] <= 16'b0000000000111010;
        weights1[37165] <= 16'b0000000000100010;
        weights1[37166] <= 16'b0000000000110110;
        weights1[37167] <= 16'b0000000000100011;
        weights1[37168] <= 16'b0000000000100111;
        weights1[37169] <= 16'b0000000000011011;
        weights1[37170] <= 16'b0000000000011110;
        weights1[37171] <= 16'b0000000000010111;
        weights1[37172] <= 16'b0000000000010111;
        weights1[37173] <= 16'b0000000000011010;
        weights1[37174] <= 16'b0000000000000011;
        weights1[37175] <= 16'b0000000000001001;
        weights1[37176] <= 16'b0000000000001000;
        weights1[37177] <= 16'b0000000000001010;
        weights1[37178] <= 16'b1111111111111101;
        weights1[37179] <= 16'b0000000000010001;
        weights1[37180] <= 16'b1111111111111100;
        weights1[37181] <= 16'b1111111111101011;
        weights1[37182] <= 16'b0000000000000101;
        weights1[37183] <= 16'b1111111111111100;
        weights1[37184] <= 16'b1111111111011010;
        weights1[37185] <= 16'b1111111111000000;
        weights1[37186] <= 16'b1111111110011101;
        weights1[37187] <= 16'b1111111110101000;
        weights1[37188] <= 16'b1111111110001001;
        weights1[37189] <= 16'b1111111110000010;
        weights1[37190] <= 16'b1111111101111110;
        weights1[37191] <= 16'b1111111110110100;
        weights1[37192] <= 16'b1111111111011100;
        weights1[37193] <= 16'b1111111111111110;
        weights1[37194] <= 16'b0000000000100000;
        weights1[37195] <= 16'b0000000000100101;
        weights1[37196] <= 16'b0000000000101010;
        weights1[37197] <= 16'b0000000000101111;
        weights1[37198] <= 16'b0000000000010011;
        weights1[37199] <= 16'b0000000000010010;
        weights1[37200] <= 16'b0000000000000111;
        weights1[37201] <= 16'b0000000000000000;
        weights1[37202] <= 16'b0000000000000010;
        weights1[37203] <= 16'b1111111111101111;
        weights1[37204] <= 16'b1111111111110111;
        weights1[37205] <= 16'b1111111111110110;
        weights1[37206] <= 16'b1111111111101101;
        weights1[37207] <= 16'b1111111111110110;
        weights1[37208] <= 16'b1111111111110110;
        weights1[37209] <= 16'b1111111111101110;
        weights1[37210] <= 16'b1111111111111010;
        weights1[37211] <= 16'b1111111111111100;
        weights1[37212] <= 16'b1111111111011111;
        weights1[37213] <= 16'b1111111111000010;
        weights1[37214] <= 16'b1111111110101111;
        weights1[37215] <= 16'b1111111110001111;
        weights1[37216] <= 16'b1111111110000010;
        weights1[37217] <= 16'b1111111101010111;
        weights1[37218] <= 16'b1111111100110110;
        weights1[37219] <= 16'b1111111100101101;
        weights1[37220] <= 16'b1111111100100000;
        weights1[37221] <= 16'b1111111101110101;
        weights1[37222] <= 16'b1111111110110100;
        weights1[37223] <= 16'b1111111111010100;
        weights1[37224] <= 16'b1111111111110111;
        weights1[37225] <= 16'b0000000000010000;
        weights1[37226] <= 16'b1111111111111011;
        weights1[37227] <= 16'b0000000000001001;
        weights1[37228] <= 16'b1111111111110000;
        weights1[37229] <= 16'b1111111111111110;
        weights1[37230] <= 16'b1111111111110100;
        weights1[37231] <= 16'b0000000000001011;
        weights1[37232] <= 16'b1111111111110101;
        weights1[37233] <= 16'b1111111111111001;
        weights1[37234] <= 16'b0000000000000101;
        weights1[37235] <= 16'b1111111111110000;
        weights1[37236] <= 16'b1111111111111011;
        weights1[37237] <= 16'b1111111111111111;
        weights1[37238] <= 16'b1111111111111101;
        weights1[37239] <= 16'b1111111111100111;
        weights1[37240] <= 16'b1111111111110111;
        weights1[37241] <= 16'b1111111111100100;
        weights1[37242] <= 16'b1111111111010110;
        weights1[37243] <= 16'b1111111111000110;
        weights1[37244] <= 16'b1111111110111110;
        weights1[37245] <= 16'b1111111110011111;
        weights1[37246] <= 16'b1111111101110011;
        weights1[37247] <= 16'b1111111101001010;
        weights1[37248] <= 16'b1111111100001001;
        weights1[37249] <= 16'b1111111011101110;
        weights1[37250] <= 16'b1111111011110100;
        weights1[37251] <= 16'b1111111100010000;
        weights1[37252] <= 16'b1111111101011000;
        weights1[37253] <= 16'b1111111110011000;
        weights1[37254] <= 16'b1111111110110001;
        weights1[37255] <= 16'b1111111111001110;
        weights1[37256] <= 16'b1111111111011111;
        weights1[37257] <= 16'b1111111111100111;
        weights1[37258] <= 16'b1111111111010101;
        weights1[37259] <= 16'b1111111111101000;
        weights1[37260] <= 16'b1111111111111111;
        weights1[37261] <= 16'b0000000000000011;
        weights1[37262] <= 16'b1111111111111111;
        weights1[37263] <= 16'b1111111111111011;
        weights1[37264] <= 16'b0000000000010000;
        weights1[37265] <= 16'b0000000000001100;
        weights1[37266] <= 16'b1111111111110010;
        weights1[37267] <= 16'b1111111111101100;
        weights1[37268] <= 16'b0000000000010000;
        weights1[37269] <= 16'b1111111111110100;
        weights1[37270] <= 16'b0000000000010001;
        weights1[37271] <= 16'b0000000000000010;
        weights1[37272] <= 16'b0000000000000010;
        weights1[37273] <= 16'b1111111111111010;
        weights1[37274] <= 16'b0000000000001010;
        weights1[37275] <= 16'b1111111111010001;
        weights1[37276] <= 16'b1111111111000100;
        weights1[37277] <= 16'b1111111110010101;
        weights1[37278] <= 16'b1111111101011111;
        weights1[37279] <= 16'b1111111101001001;
        weights1[37280] <= 16'b1111111101011011;
        weights1[37281] <= 16'b1111111101100011;
        weights1[37282] <= 16'b1111111110010000;
        weights1[37283] <= 16'b1111111110010101;
        weights1[37284] <= 16'b1111111111000000;
        weights1[37285] <= 16'b1111111110111000;
        weights1[37286] <= 16'b1111111111110100;
        weights1[37287] <= 16'b1111111111110111;
        weights1[37288] <= 16'b1111111111101111;
        weights1[37289] <= 16'b1111111111111101;
        weights1[37290] <= 16'b0000000000000100;
        weights1[37291] <= 16'b1111111111111001;
        weights1[37292] <= 16'b0000000000000111;
        weights1[37293] <= 16'b0000000000010101;
        weights1[37294] <= 16'b0000000000010001;
        weights1[37295] <= 16'b1111111111101111;
        weights1[37296] <= 16'b0000000000011101;
        weights1[37297] <= 16'b0000000000010011;
        weights1[37298] <= 16'b0000000000100101;
        weights1[37299] <= 16'b0000000000010111;
        weights1[37300] <= 16'b0000000000111011;
        weights1[37301] <= 16'b0000000000100100;
        weights1[37302] <= 16'b0000000000101010;
        weights1[37303] <= 16'b0000000001000011;
        weights1[37304] <= 16'b0000000000101001;
        weights1[37305] <= 16'b0000000000101001;
        weights1[37306] <= 16'b0000000000001101;
        weights1[37307] <= 16'b0000000000001110;
        weights1[37308] <= 16'b1111111111110100;
        weights1[37309] <= 16'b1111111111110101;
        weights1[37310] <= 16'b1111111111011110;
        weights1[37311] <= 16'b1111111111100000;
        weights1[37312] <= 16'b1111111111010100;
        weights1[37313] <= 16'b1111111111011011;
        weights1[37314] <= 16'b1111111111101001;
        weights1[37315] <= 16'b1111111111110000;
        weights1[37316] <= 16'b1111111111111011;
        weights1[37317] <= 16'b1111111111110010;
        weights1[37318] <= 16'b0000000000000010;
        weights1[37319] <= 16'b0000000000000000;
        weights1[37320] <= 16'b0000000000001000;
        weights1[37321] <= 16'b0000000000000000;
        weights1[37322] <= 16'b1111111111111100;
        weights1[37323] <= 16'b1111111111110011;
        weights1[37324] <= 16'b0000000000100010;
        weights1[37325] <= 16'b0000000000100110;
        weights1[37326] <= 16'b0000000000100111;
        weights1[37327] <= 16'b0000000000101000;
        weights1[37328] <= 16'b0000000000101110;
        weights1[37329] <= 16'b0000000000111000;
        weights1[37330] <= 16'b0000000000110110;
        weights1[37331] <= 16'b0000000001000001;
        weights1[37332] <= 16'b0000000001011110;
        weights1[37333] <= 16'b0000000001000001;
        weights1[37334] <= 16'b0000000001001110;
        weights1[37335] <= 16'b0000000001010001;
        weights1[37336] <= 16'b0000000000101010;
        weights1[37337] <= 16'b0000000000100100;
        weights1[37338] <= 16'b1111111111111110;
        weights1[37339] <= 16'b0000000000001011;
        weights1[37340] <= 16'b0000000000000100;
        weights1[37341] <= 16'b0000000000001100;
        weights1[37342] <= 16'b1111111111101111;
        weights1[37343] <= 16'b0000000000001001;
        weights1[37344] <= 16'b1111111111101000;
        weights1[37345] <= 16'b1111111111110001;
        weights1[37346] <= 16'b1111111111110110;
        weights1[37347] <= 16'b1111111111111010;
        weights1[37348] <= 16'b1111111111110000;
        weights1[37349] <= 16'b1111111111110101;
        weights1[37350] <= 16'b1111111111101110;
        weights1[37351] <= 16'b1111111111111011;
        weights1[37352] <= 16'b0000000000101000;
        weights1[37353] <= 16'b0000000000011100;
        weights1[37354] <= 16'b0000000000101110;
        weights1[37355] <= 16'b0000000000111110;
        weights1[37356] <= 16'b0000000000100000;
        weights1[37357] <= 16'b1111111111111111;
        weights1[37358] <= 16'b0000000000110011;
        weights1[37359] <= 16'b0000000000101100;
        weights1[37360] <= 16'b0000000000100011;
        weights1[37361] <= 16'b0000000000101100;
        weights1[37362] <= 16'b0000000000101101;
        weights1[37363] <= 16'b0000000000110011;
        weights1[37364] <= 16'b0000000000101010;
        weights1[37365] <= 16'b0000000000001111;
        weights1[37366] <= 16'b0000000000010011;
        weights1[37367] <= 16'b0000000000011100;
        weights1[37368] <= 16'b1111111111111000;
        weights1[37369] <= 16'b0000000000000010;
        weights1[37370] <= 16'b1111111111110101;
        weights1[37371] <= 16'b1111111111110000;
        weights1[37372] <= 16'b1111111111110110;
        weights1[37373] <= 16'b1111111111111110;
        weights1[37374] <= 16'b1111111111111100;
        weights1[37375] <= 16'b1111111111111001;
        weights1[37376] <= 16'b0000000000001110;
        weights1[37377] <= 16'b0000000000000010;
        weights1[37378] <= 16'b1111111111110000;
        weights1[37379] <= 16'b0000000000001010;
        weights1[37380] <= 16'b0000000000001011;
        weights1[37381] <= 16'b0000000000000101;
        weights1[37382] <= 16'b0000000000011000;
        weights1[37383] <= 16'b0000000000101110;
        weights1[37384] <= 16'b0000000000011000;
        weights1[37385] <= 16'b0000000000001101;
        weights1[37386] <= 16'b0000000000100110;
        weights1[37387] <= 16'b0000000000011000;
        weights1[37388] <= 16'b0000000000001010;
        weights1[37389] <= 16'b0000000000011010;
        weights1[37390] <= 16'b0000000000100001;
        weights1[37391] <= 16'b0000000000011001;
        weights1[37392] <= 16'b0000000000100010;
        weights1[37393] <= 16'b0000000000011111;
        weights1[37394] <= 16'b0000000000010011;
        weights1[37395] <= 16'b0000000000001011;
        weights1[37396] <= 16'b0000000000010100;
        weights1[37397] <= 16'b0000000000010011;
        weights1[37398] <= 16'b0000000000000111;
        weights1[37399] <= 16'b0000000000001001;
        weights1[37400] <= 16'b1111111111110111;
        weights1[37401] <= 16'b1111111111111100;
        weights1[37402] <= 16'b1111111111011111;
        weights1[37403] <= 16'b1111111111110101;
        weights1[37404] <= 16'b1111111111100111;
        weights1[37405] <= 16'b1111111111101000;
        weights1[37406] <= 16'b1111111111110001;
        weights1[37407] <= 16'b1111111111111111;
        weights1[37408] <= 16'b0000000000000010;
        weights1[37409] <= 16'b0000000000001000;
        weights1[37410] <= 16'b0000000000000111;
        weights1[37411] <= 16'b1111111111111000;
        weights1[37412] <= 16'b1111111111001101;
        weights1[37413] <= 16'b0000000000000100;
        weights1[37414] <= 16'b1111111111111000;
        weights1[37415] <= 16'b0000000000011101;
        weights1[37416] <= 16'b0000000000101111;
        weights1[37417] <= 16'b0000000000000100;
        weights1[37418] <= 16'b0000000000000111;
        weights1[37419] <= 16'b0000000000000110;
        weights1[37420] <= 16'b0000000000001110;
        weights1[37421] <= 16'b0000000000010101;
        weights1[37422] <= 16'b0000000000000110;
        weights1[37423] <= 16'b0000000000010010;
        weights1[37424] <= 16'b0000000000010000;
        weights1[37425] <= 16'b1111111111111001;
        weights1[37426] <= 16'b0000000000000101;
        weights1[37427] <= 16'b0000000000001101;
        weights1[37428] <= 16'b0000000000001000;
        weights1[37429] <= 16'b0000000000001001;
        weights1[37430] <= 16'b0000000000001001;
        weights1[37431] <= 16'b1111111111110010;
        weights1[37432] <= 16'b1111111111110001;
        weights1[37433] <= 16'b1111111111110011;
        weights1[37434] <= 16'b1111111111111100;
        weights1[37435] <= 16'b1111111111111010;
        weights1[37436] <= 16'b0000000000000100;
        weights1[37437] <= 16'b0000000000000101;
        weights1[37438] <= 16'b0000000000001101;
        weights1[37439] <= 16'b1111111111101101;
        weights1[37440] <= 16'b1111111111100011;
        weights1[37441] <= 16'b1111111111100101;
        weights1[37442] <= 16'b1111111111100001;
        weights1[37443] <= 16'b1111111111111000;
        weights1[37444] <= 16'b0000000000000001;
        weights1[37445] <= 16'b1111111111111101;
        weights1[37446] <= 16'b1111111111101111;
        weights1[37447] <= 16'b0000000000000000;
        weights1[37448] <= 16'b0000000000000100;
        weights1[37449] <= 16'b1111111111110110;
        weights1[37450] <= 16'b1111111111110101;
        weights1[37451] <= 16'b1111111111111110;
        weights1[37452] <= 16'b1111111111110010;
        weights1[37453] <= 16'b0000000000011010;
        weights1[37454] <= 16'b1111111111111110;
        weights1[37455] <= 16'b0000000000001000;
        weights1[37456] <= 16'b1111111111110101;
        weights1[37457] <= 16'b1111111111111111;
        weights1[37458] <= 16'b1111111111110110;
        weights1[37459] <= 16'b0000000000000010;
        weights1[37460] <= 16'b0000000000000110;
        weights1[37461] <= 16'b0000000000000000;
        weights1[37462] <= 16'b0000000000000001;
        weights1[37463] <= 16'b1111111111111011;
        weights1[37464] <= 16'b1111111111111000;
        weights1[37465] <= 16'b0000000000000011;
        weights1[37466] <= 16'b0000000000001100;
        weights1[37467] <= 16'b0000000000001110;
        weights1[37468] <= 16'b1111111111101101;
        weights1[37469] <= 16'b1111111111100011;
        weights1[37470] <= 16'b1111111111101110;
        weights1[37471] <= 16'b1111111111101111;
        weights1[37472] <= 16'b1111111111110001;
        weights1[37473] <= 16'b0000000000000000;
        weights1[37474] <= 16'b1111111111111110;
        weights1[37475] <= 16'b1111111111110100;
        weights1[37476] <= 16'b1111111111110111;
        weights1[37477] <= 16'b0000000000001001;
        weights1[37478] <= 16'b0000000000000000;
        weights1[37479] <= 16'b0000000000011000;
        weights1[37480] <= 16'b0000000000001000;
        weights1[37481] <= 16'b1111111111111011;
        weights1[37482] <= 16'b1111111111110110;
        weights1[37483] <= 16'b1111111111110101;
        weights1[37484] <= 16'b1111111111111010;
        weights1[37485] <= 16'b0000000000001001;
        weights1[37486] <= 16'b0000000000001001;
        weights1[37487] <= 16'b0000000000001011;
        weights1[37488] <= 16'b0000000000000100;
        weights1[37489] <= 16'b0000000000001101;
        weights1[37490] <= 16'b0000000000000011;
        weights1[37491] <= 16'b0000000000000110;
        weights1[37492] <= 16'b1111111111111101;
        weights1[37493] <= 16'b0000000000000011;
        weights1[37494] <= 16'b0000000000000101;
        weights1[37495] <= 16'b0000000000000100;
        weights1[37496] <= 16'b1111111111110010;
        weights1[37497] <= 16'b1111111111101001;
        weights1[37498] <= 16'b1111111111011111;
        weights1[37499] <= 16'b1111111111000011;
        weights1[37500] <= 16'b1111111111100011;
        weights1[37501] <= 16'b1111111111101001;
        weights1[37502] <= 16'b1111111111110100;
        weights1[37503] <= 16'b0000000000000100;
        weights1[37504] <= 16'b0000000000000100;
        weights1[37505] <= 16'b1111111111111101;
        weights1[37506] <= 16'b1111111111100101;
        weights1[37507] <= 16'b1111111111101101;
        weights1[37508] <= 16'b0000000000000000;
        weights1[37509] <= 16'b1111111111110011;
        weights1[37510] <= 16'b1111111111111011;
        weights1[37511] <= 16'b0000000000100010;
        weights1[37512] <= 16'b0000000000001101;
        weights1[37513] <= 16'b0000000000010001;
        weights1[37514] <= 16'b0000000000011010;
        weights1[37515] <= 16'b0000000000010010;
        weights1[37516] <= 16'b0000000000011011;
        weights1[37517] <= 16'b0000000000011101;
        weights1[37518] <= 16'b0000000000000101;
        weights1[37519] <= 16'b0000000000000100;
        weights1[37520] <= 16'b0000000000000000;
        weights1[37521] <= 16'b1111111111111101;
        weights1[37522] <= 16'b0000000000000111;
        weights1[37523] <= 16'b1111111111111101;
        weights1[37524] <= 16'b1111111111111110;
        weights1[37525] <= 16'b0000000000000100;
        weights1[37526] <= 16'b1111111111101011;
        weights1[37527] <= 16'b1111111111011010;
        weights1[37528] <= 16'b1111111111001101;
        weights1[37529] <= 16'b1111111111001111;
        weights1[37530] <= 16'b1111111111001101;
        weights1[37531] <= 16'b1111111111011100;
        weights1[37532] <= 16'b1111111111011010;
        weights1[37533] <= 16'b1111111111100100;
        weights1[37534] <= 16'b1111111111111010;
        weights1[37535] <= 16'b1111111111101100;
        weights1[37536] <= 16'b1111111111110010;
        weights1[37537] <= 16'b1111111111111001;
        weights1[37538] <= 16'b0000000000011000;
        weights1[37539] <= 16'b0000000000010001;
        weights1[37540] <= 16'b1111111111111101;
        weights1[37541] <= 16'b0000000000001101;
        weights1[37542] <= 16'b0000000000001100;
        weights1[37543] <= 16'b0000000000001000;
        weights1[37544] <= 16'b0000000000100011;
        weights1[37545] <= 16'b0000000000010110;
        weights1[37546] <= 16'b0000000000001110;
        weights1[37547] <= 16'b0000000000000010;
        weights1[37548] <= 16'b1111111111111111;
        weights1[37549] <= 16'b1111111111111100;
        weights1[37550] <= 16'b0000000000000110;
        weights1[37551] <= 16'b1111111111111100;
        weights1[37552] <= 16'b0000000000001110;
        weights1[37553] <= 16'b1111111111110101;
        weights1[37554] <= 16'b1111111111111000;
        weights1[37555] <= 16'b1111111111111110;
        weights1[37556] <= 16'b1111111111110100;
        weights1[37557] <= 16'b0000000000000110;
        weights1[37558] <= 16'b1111111111101011;
        weights1[37559] <= 16'b1111111111101111;
        weights1[37560] <= 16'b1111111111111010;
        weights1[37561] <= 16'b1111111111101110;
        weights1[37562] <= 16'b1111111111110110;
        weights1[37563] <= 16'b0000000000001110;
        weights1[37564] <= 16'b1111111111111100;
        weights1[37565] <= 16'b0000000000001101;
        weights1[37566] <= 16'b1111111111111101;
        weights1[37567] <= 16'b0000000000000111;
        weights1[37568] <= 16'b0000000000001000;
        weights1[37569] <= 16'b0000000000000000;
        weights1[37570] <= 16'b0000000000001010;
        weights1[37571] <= 16'b0000000000001110;
        weights1[37572] <= 16'b0000000000010001;
        weights1[37573] <= 16'b0000000000001100;
        weights1[37574] <= 16'b1111111111111111;
        weights1[37575] <= 16'b0000000000000001;
        weights1[37576] <= 16'b0000000000000110;
        weights1[37577] <= 16'b0000000000000100;
        weights1[37578] <= 16'b0000000000000100;
        weights1[37579] <= 16'b0000000000000011;
        weights1[37580] <= 16'b0000000000001111;
        weights1[37581] <= 16'b1111111111110111;
        weights1[37582] <= 16'b0000000000011110;
        weights1[37583] <= 16'b0000000000000111;
        weights1[37584] <= 16'b0000000000011000;
        weights1[37585] <= 16'b0000000000100010;
        weights1[37586] <= 16'b0000000000101100;
        weights1[37587] <= 16'b0000000000110010;
        weights1[37588] <= 16'b0000000000010100;
        weights1[37589] <= 16'b0000000000010110;
        weights1[37590] <= 16'b0000000000010001;
        weights1[37591] <= 16'b0000000000010101;
        weights1[37592] <= 16'b0000000000001000;
        weights1[37593] <= 16'b0000000000001011;
        weights1[37594] <= 16'b0000000000010101;
        weights1[37595] <= 16'b1111111111110100;
        weights1[37596] <= 16'b1111111111110111;
        weights1[37597] <= 16'b0000000000001110;
        weights1[37598] <= 16'b0000000000011000;
        weights1[37599] <= 16'b0000000000000110;
        weights1[37600] <= 16'b0000000000000010;
        weights1[37601] <= 16'b0000000000000011;
        weights1[37602] <= 16'b0000000000000000;
        weights1[37603] <= 16'b1111111111111111;
        weights1[37604] <= 16'b0000000000000100;
        weights1[37605] <= 16'b0000000000000010;
        weights1[37606] <= 16'b0000000000000100;
        weights1[37607] <= 16'b0000000000010011;
        weights1[37608] <= 16'b0000000000011000;
        weights1[37609] <= 16'b0000000000010111;
        weights1[37610] <= 16'b0000000000101101;
        weights1[37611] <= 16'b0000000000101011;
        weights1[37612] <= 16'b0000000000100100;
        weights1[37613] <= 16'b0000000000101011;
        weights1[37614] <= 16'b0000000000100110;
        weights1[37615] <= 16'b0000000000010110;
        weights1[37616] <= 16'b0000000000011111;
        weights1[37617] <= 16'b0000000000011101;
        weights1[37618] <= 16'b0000000000011111;
        weights1[37619] <= 16'b0000000000011000;
        weights1[37620] <= 16'b0000000000001101;
        weights1[37621] <= 16'b0000000000011001;
        weights1[37622] <= 16'b0000000000001101;
        weights1[37623] <= 16'b0000000000000111;
        weights1[37624] <= 16'b0000000000001010;
        weights1[37625] <= 16'b0000000000011010;
        weights1[37626] <= 16'b0000000000010001;
        weights1[37627] <= 16'b0000000000001000;
        weights1[37628] <= 16'b0000000000000001;
        weights1[37629] <= 16'b0000000000000001;
        weights1[37630] <= 16'b1111111111111111;
        weights1[37631] <= 16'b0000000000000000;
        weights1[37632] <= 16'b1111111111111111;
        weights1[37633] <= 16'b1111111111111110;
        weights1[37634] <= 16'b1111111111111110;
        weights1[37635] <= 16'b1111111111111100;
        weights1[37636] <= 16'b1111111111111110;
        weights1[37637] <= 16'b1111111111111101;
        weights1[37638] <= 16'b0000000000000101;
        weights1[37639] <= 16'b0000000000010011;
        weights1[37640] <= 16'b0000000000000110;
        weights1[37641] <= 16'b0000000000000111;
        weights1[37642] <= 16'b1111111111111010;
        weights1[37643] <= 16'b0000000000000010;
        weights1[37644] <= 16'b1111111111111100;
        weights1[37645] <= 16'b1111111111111110;
        weights1[37646] <= 16'b1111111111111001;
        weights1[37647] <= 16'b1111111111111000;
        weights1[37648] <= 16'b1111111111101111;
        weights1[37649] <= 16'b1111111111110111;
        weights1[37650] <= 16'b1111111111111011;
        weights1[37651] <= 16'b1111111111111011;
        weights1[37652] <= 16'b0000000000000000;
        weights1[37653] <= 16'b0000000000000101;
        weights1[37654] <= 16'b0000000000000010;
        weights1[37655] <= 16'b0000000000000001;
        weights1[37656] <= 16'b0000000000000000;
        weights1[37657] <= 16'b1111111111111000;
        weights1[37658] <= 16'b1111111111111101;
        weights1[37659] <= 16'b0000000000000000;
        weights1[37660] <= 16'b0000000000000001;
        weights1[37661] <= 16'b1111111111111111;
        weights1[37662] <= 16'b1111111111111100;
        weights1[37663] <= 16'b1111111111111011;
        weights1[37664] <= 16'b0000000000000011;
        weights1[37665] <= 16'b0000000000000010;
        weights1[37666] <= 16'b0000000000000100;
        weights1[37667] <= 16'b0000000000001100;
        weights1[37668] <= 16'b0000000000010000;
        weights1[37669] <= 16'b0000000000001011;
        weights1[37670] <= 16'b1111111111110100;
        weights1[37671] <= 16'b0000000000000000;
        weights1[37672] <= 16'b1111111111111100;
        weights1[37673] <= 16'b1111111111100110;
        weights1[37674] <= 16'b0000000000000110;
        weights1[37675] <= 16'b1111111111111001;
        weights1[37676] <= 16'b1111111111101011;
        weights1[37677] <= 16'b1111111111110000;
        weights1[37678] <= 16'b0000000000000111;
        weights1[37679] <= 16'b0000000000000100;
        weights1[37680] <= 16'b1111111111111101;
        weights1[37681] <= 16'b1111111111111111;
        weights1[37682] <= 16'b0000000000001100;
        weights1[37683] <= 16'b0000000000001000;
        weights1[37684] <= 16'b1111111111110100;
        weights1[37685] <= 16'b1111111111110100;
        weights1[37686] <= 16'b1111111111111100;
        weights1[37687] <= 16'b0000000000000000;
        weights1[37688] <= 16'b1111111111111111;
        weights1[37689] <= 16'b1111111111111110;
        weights1[37690] <= 16'b1111111111111010;
        weights1[37691] <= 16'b0000000000001000;
        weights1[37692] <= 16'b0000000000000001;
        weights1[37693] <= 16'b0000000000000000;
        weights1[37694] <= 16'b1111111111111011;
        weights1[37695] <= 16'b0000000000001100;
        weights1[37696] <= 16'b0000000000000101;
        weights1[37697] <= 16'b1111111111111101;
        weights1[37698] <= 16'b0000000000000111;
        weights1[37699] <= 16'b1111111111111010;
        weights1[37700] <= 16'b1111111111111011;
        weights1[37701] <= 16'b1111111111100111;
        weights1[37702] <= 16'b1111111111101001;
        weights1[37703] <= 16'b1111111111110001;
        weights1[37704] <= 16'b0000000000000100;
        weights1[37705] <= 16'b0000000000000010;
        weights1[37706] <= 16'b0000000000001100;
        weights1[37707] <= 16'b1111111111101000;
        weights1[37708] <= 16'b0000000000001000;
        weights1[37709] <= 16'b1111111111111101;
        weights1[37710] <= 16'b0000000000000001;
        weights1[37711] <= 16'b1111111111111101;
        weights1[37712] <= 16'b1111111111110101;
        weights1[37713] <= 16'b1111111111110101;
        weights1[37714] <= 16'b1111111111111111;
        weights1[37715] <= 16'b1111111111111111;
        weights1[37716] <= 16'b1111111111111101;
        weights1[37717] <= 16'b1111111111111100;
        weights1[37718] <= 16'b0000000000000001;
        weights1[37719] <= 16'b0000000000000000;
        weights1[37720] <= 16'b1111111111111101;
        weights1[37721] <= 16'b0000000000001010;
        weights1[37722] <= 16'b0000000000000001;
        weights1[37723] <= 16'b1111111111110110;
        weights1[37724] <= 16'b1111111111110100;
        weights1[37725] <= 16'b1111111111111101;
        weights1[37726] <= 16'b1111111111011111;
        weights1[37727] <= 16'b0000000000000100;
        weights1[37728] <= 16'b1111111111110111;
        weights1[37729] <= 16'b0000000000000010;
        weights1[37730] <= 16'b0000000000010000;
        weights1[37731] <= 16'b0000000000000010;
        weights1[37732] <= 16'b0000000000001001;
        weights1[37733] <= 16'b1111111111111010;
        weights1[37734] <= 16'b0000000000010001;
        weights1[37735] <= 16'b0000000000001000;
        weights1[37736] <= 16'b0000000000010011;
        weights1[37737] <= 16'b0000000000001100;
        weights1[37738] <= 16'b0000000000000001;
        weights1[37739] <= 16'b1111111111111101;
        weights1[37740] <= 16'b0000000000000101;
        weights1[37741] <= 16'b0000000000001101;
        weights1[37742] <= 16'b0000000000001010;
        weights1[37743] <= 16'b0000000000000101;
        weights1[37744] <= 16'b1111111111111011;
        weights1[37745] <= 16'b1111111111111011;
        weights1[37746] <= 16'b1111111111111101;
        weights1[37747] <= 16'b0000000000000101;
        weights1[37748] <= 16'b1111111111111010;
        weights1[37749] <= 16'b0000000000001010;
        weights1[37750] <= 16'b0000000000001000;
        weights1[37751] <= 16'b0000000000000100;
        weights1[37752] <= 16'b1111111111111110;
        weights1[37753] <= 16'b0000000000000110;
        weights1[37754] <= 16'b1111111111111101;
        weights1[37755] <= 16'b1111111111111001;
        weights1[37756] <= 16'b1111111111111110;
        weights1[37757] <= 16'b1111111111111100;
        weights1[37758] <= 16'b1111111111101010;
        weights1[37759] <= 16'b0000000000000001;
        weights1[37760] <= 16'b1111111111111000;
        weights1[37761] <= 16'b0000000000000001;
        weights1[37762] <= 16'b0000000000001100;
        weights1[37763] <= 16'b0000000000001000;
        weights1[37764] <= 16'b1111111111101111;
        weights1[37765] <= 16'b1111111111111101;
        weights1[37766] <= 16'b1111111111110111;
        weights1[37767] <= 16'b0000000000001010;
        weights1[37768] <= 16'b1111111111110101;
        weights1[37769] <= 16'b1111111111111110;
        weights1[37770] <= 16'b0000000000000100;
        weights1[37771] <= 16'b1111111111111101;
        weights1[37772] <= 16'b1111111111111010;
        weights1[37773] <= 16'b1111111111110110;
        weights1[37774] <= 16'b0000000000001010;
        weights1[37775] <= 16'b1111111111110111;
        weights1[37776] <= 16'b0000000000000011;
        weights1[37777] <= 16'b1111111111110111;
        weights1[37778] <= 16'b1111111111100101;
        weights1[37779] <= 16'b1111111111111100;
        weights1[37780] <= 16'b1111111111101111;
        weights1[37781] <= 16'b0000000000010010;
        weights1[37782] <= 16'b0000000000100001;
        weights1[37783] <= 16'b1111111111111100;
        weights1[37784] <= 16'b1111111111101111;
        weights1[37785] <= 16'b1111111111110100;
        weights1[37786] <= 16'b0000000000000001;
        weights1[37787] <= 16'b1111111111100001;
        weights1[37788] <= 16'b0000000000000001;
        weights1[37789] <= 16'b1111111111110100;
        weights1[37790] <= 16'b1111111111111111;
        weights1[37791] <= 16'b1111111111111001;
        weights1[37792] <= 16'b0000000000001010;
        weights1[37793] <= 16'b1111111111111000;
        weights1[37794] <= 16'b1111111111111110;
        weights1[37795] <= 16'b1111111111110100;
        weights1[37796] <= 16'b1111111111100101;
        weights1[37797] <= 16'b0000000000010010;
        weights1[37798] <= 16'b0000000000000001;
        weights1[37799] <= 16'b1111111111111110;
        weights1[37800] <= 16'b0000000000000000;
        weights1[37801] <= 16'b1111111111111100;
        weights1[37802] <= 16'b0000000000001010;
        weights1[37803] <= 16'b0000000000000000;
        weights1[37804] <= 16'b1111111111111101;
        weights1[37805] <= 16'b0000000000000011;
        weights1[37806] <= 16'b1111111111111000;
        weights1[37807] <= 16'b0000000000001010;
        weights1[37808] <= 16'b1111111111110111;
        weights1[37809] <= 16'b1111111111100011;
        weights1[37810] <= 16'b1111111111111001;
        weights1[37811] <= 16'b1111111111011101;
        weights1[37812] <= 16'b1111111111111010;
        weights1[37813] <= 16'b1111111111110111;
        weights1[37814] <= 16'b1111111111111110;
        weights1[37815] <= 16'b0000000000001001;
        weights1[37816] <= 16'b1111111111110100;
        weights1[37817] <= 16'b1111111111111001;
        weights1[37818] <= 16'b0000000000000010;
        weights1[37819] <= 16'b1111111111111001;
        weights1[37820] <= 16'b1111111111111111;
        weights1[37821] <= 16'b1111111111111010;
        weights1[37822] <= 16'b1111111111111100;
        weights1[37823] <= 16'b0000000000001100;
        weights1[37824] <= 16'b0000000000000101;
        weights1[37825] <= 16'b1111111111111100;
        weights1[37826] <= 16'b1111111111111111;
        weights1[37827] <= 16'b0000000000000011;
        weights1[37828] <= 16'b1111111111110110;
        weights1[37829] <= 16'b1111111111110110;
        weights1[37830] <= 16'b0000000000001000;
        weights1[37831] <= 16'b1111111111110001;
        weights1[37832] <= 16'b0000000000010001;
        weights1[37833] <= 16'b0000000000001000;
        weights1[37834] <= 16'b0000000000000111;
        weights1[37835] <= 16'b1111111111101010;
        weights1[37836] <= 16'b0000000000000100;
        weights1[37837] <= 16'b1111111111110111;
        weights1[37838] <= 16'b1111111111111010;
        weights1[37839] <= 16'b0000000000001010;
        weights1[37840] <= 16'b1111111111110100;
        weights1[37841] <= 16'b1111111111111111;
        weights1[37842] <= 16'b1111111111111010;
        weights1[37843] <= 16'b1111111111110100;
        weights1[37844] <= 16'b0000000000000010;
        weights1[37845] <= 16'b0000000000000100;
        weights1[37846] <= 16'b1111111111110101;
        weights1[37847] <= 16'b0000000000000110;
        weights1[37848] <= 16'b1111111111110101;
        weights1[37849] <= 16'b1111111111110101;
        weights1[37850] <= 16'b0000000000001110;
        weights1[37851] <= 16'b1111111111111100;
        weights1[37852] <= 16'b1111111111110101;
        weights1[37853] <= 16'b1111111111101111;
        weights1[37854] <= 16'b0000000000000001;
        weights1[37855] <= 16'b0000000000000010;
        weights1[37856] <= 16'b1111111111111001;
        weights1[37857] <= 16'b1111111111110100;
        weights1[37858] <= 16'b1111111111110101;
        weights1[37859] <= 16'b0000000000000010;
        weights1[37860] <= 16'b0000000000001101;
        weights1[37861] <= 16'b1111111111111010;
        weights1[37862] <= 16'b0000000000000010;
        weights1[37863] <= 16'b1111111111111111;
        weights1[37864] <= 16'b1111111111110111;
        weights1[37865] <= 16'b0000000000010000;
        weights1[37866] <= 16'b1111111111110111;
        weights1[37867] <= 16'b1111111111101111;
        weights1[37868] <= 16'b0000000000001000;
        weights1[37869] <= 16'b1111111111110111;
        weights1[37870] <= 16'b0000000000010101;
        weights1[37871] <= 16'b0000000000001111;
        weights1[37872] <= 16'b1111111111111101;
        weights1[37873] <= 16'b0000000000000011;
        weights1[37874] <= 16'b1111111111110111;
        weights1[37875] <= 16'b1111111111111101;
        weights1[37876] <= 16'b0000000000001111;
        weights1[37877] <= 16'b1111111111010100;
        weights1[37878] <= 16'b0000000000000110;
        weights1[37879] <= 16'b1111111111111011;
        weights1[37880] <= 16'b1111111111101110;
        weights1[37881] <= 16'b1111111111110001;
        weights1[37882] <= 16'b1111111111111010;
        weights1[37883] <= 16'b1111111111111101;
        weights1[37884] <= 16'b1111111111111100;
        weights1[37885] <= 16'b0000000000000001;
        weights1[37886] <= 16'b1111111111111111;
        weights1[37887] <= 16'b1111111111111011;
        weights1[37888] <= 16'b1111111111110100;
        weights1[37889] <= 16'b1111111111111100;
        weights1[37890] <= 16'b1111111111111110;
        weights1[37891] <= 16'b0000000000000100;
        weights1[37892] <= 16'b0000000000000001;
        weights1[37893] <= 16'b1111111111111110;
        weights1[37894] <= 16'b1111111111111100;
        weights1[37895] <= 16'b1111111111111011;
        weights1[37896] <= 16'b1111111111110101;
        weights1[37897] <= 16'b1111111111111101;
        weights1[37898] <= 16'b1111111111100010;
        weights1[37899] <= 16'b1111111111111101;
        weights1[37900] <= 16'b1111111111111111;
        weights1[37901] <= 16'b1111111111101100;
        weights1[37902] <= 16'b1111111111111100;
        weights1[37903] <= 16'b1111111111110111;
        weights1[37904] <= 16'b0000000000000010;
        weights1[37905] <= 16'b1111111111101101;
        weights1[37906] <= 16'b0000000000010101;
        weights1[37907] <= 16'b1111111111110011;
        weights1[37908] <= 16'b1111111111111010;
        weights1[37909] <= 16'b0000000000000001;
        weights1[37910] <= 16'b1111111111101111;
        weights1[37911] <= 16'b0000000000000000;
        weights1[37912] <= 16'b1111111111111010;
        weights1[37913] <= 16'b0000000000011000;
        weights1[37914] <= 16'b0000000000000001;
        weights1[37915] <= 16'b0000000000000001;
        weights1[37916] <= 16'b1111111111110110;
        weights1[37917] <= 16'b1111111111110010;
        weights1[37918] <= 16'b0000000000000101;
        weights1[37919] <= 16'b1111111111110000;
        weights1[37920] <= 16'b1111111111111010;
        weights1[37921] <= 16'b1111111111110000;
        weights1[37922] <= 16'b1111111111111000;
        weights1[37923] <= 16'b1111111111110111;
        weights1[37924] <= 16'b0000000000001000;
        weights1[37925] <= 16'b1111111111111101;
        weights1[37926] <= 16'b1111111111111011;
        weights1[37927] <= 16'b1111111111101110;
        weights1[37928] <= 16'b1111111111111110;
        weights1[37929] <= 16'b1111111111111110;
        weights1[37930] <= 16'b0000000000000001;
        weights1[37931] <= 16'b1111111111101111;
        weights1[37932] <= 16'b0000000000000101;
        weights1[37933] <= 16'b1111111111111100;
        weights1[37934] <= 16'b1111111111101111;
        weights1[37935] <= 16'b1111111111101011;
        weights1[37936] <= 16'b1111111111101110;
        weights1[37937] <= 16'b1111111111010100;
        weights1[37938] <= 16'b1111111111110111;
        weights1[37939] <= 16'b1111111111101011;
        weights1[37940] <= 16'b1111111111110111;
        weights1[37941] <= 16'b1111111111111110;
        weights1[37942] <= 16'b1111111111110101;
        weights1[37943] <= 16'b1111111111111110;
        weights1[37944] <= 16'b1111111111111111;
        weights1[37945] <= 16'b1111111111101010;
        weights1[37946] <= 16'b0000000000000110;
        weights1[37947] <= 16'b1111111111111010;
        weights1[37948] <= 16'b1111111111111100;
        weights1[37949] <= 16'b1111111111101000;
        weights1[37950] <= 16'b0000000000000110;
        weights1[37951] <= 16'b1111111111110111;
        weights1[37952] <= 16'b1111111111111010;
        weights1[37953] <= 16'b0000000000000000;
        weights1[37954] <= 16'b0000000000000010;
        weights1[37955] <= 16'b0000000000000001;
        weights1[37956] <= 16'b1111111111101011;
        weights1[37957] <= 16'b1111111111111111;
        weights1[37958] <= 16'b1111111111101111;
        weights1[37959] <= 16'b1111111111111110;
        weights1[37960] <= 16'b1111111111011011;
        weights1[37961] <= 16'b1111111111100110;
        weights1[37962] <= 16'b1111111111100000;
        weights1[37963] <= 16'b1111111111011001;
        weights1[37964] <= 16'b1111111111001111;
        weights1[37965] <= 16'b1111111111101011;
        weights1[37966] <= 16'b1111111111110101;
        weights1[37967] <= 16'b1111111111100001;
        weights1[37968] <= 16'b1111111111110100;
        weights1[37969] <= 16'b1111111111111011;
        weights1[37970] <= 16'b1111111111101011;
        weights1[37971] <= 16'b0000000000000110;
        weights1[37972] <= 16'b1111111111101111;
        weights1[37973] <= 16'b1111111111111001;
        weights1[37974] <= 16'b1111111111111011;
        weights1[37975] <= 16'b0000000000000011;
        weights1[37976] <= 16'b1111111111111101;
        weights1[37977] <= 16'b0000000000001000;
        weights1[37978] <= 16'b0000000000000110;
        weights1[37979] <= 16'b0000000000001011;
        weights1[37980] <= 16'b0000000000010010;
        weights1[37981] <= 16'b1111111111111010;
        weights1[37982] <= 16'b1111111111111101;
        weights1[37983] <= 16'b0000000000000000;
        weights1[37984] <= 16'b0000000000000000;
        weights1[37985] <= 16'b1111111111101110;
        weights1[37986] <= 16'b1111111111101101;
        weights1[37987] <= 16'b1111111111110011;
        weights1[37988] <= 16'b1111111111110010;
        weights1[37989] <= 16'b0000000000000101;
        weights1[37990] <= 16'b0000000000000100;
        weights1[37991] <= 16'b1111111111110000;
        weights1[37992] <= 16'b1111111111101101;
        weights1[37993] <= 16'b1111111111100100;
        weights1[37994] <= 16'b1111111111101010;
        weights1[37995] <= 16'b1111111111101001;
        weights1[37996] <= 16'b1111111111110111;
        weights1[37997] <= 16'b0000000000001011;
        weights1[37998] <= 16'b1111111111101101;
        weights1[37999] <= 16'b0000000000000011;
        weights1[38000] <= 16'b1111111111110001;
        weights1[38001] <= 16'b0000000000000101;
        weights1[38002] <= 16'b1111111111111000;
        weights1[38003] <= 16'b1111111111111000;
        weights1[38004] <= 16'b1111111111110110;
        weights1[38005] <= 16'b0000000000000000;
        weights1[38006] <= 16'b1111111111111011;
        weights1[38007] <= 16'b1111111111110010;
        weights1[38008] <= 16'b1111111111111110;
        weights1[38009] <= 16'b1111111111111111;
        weights1[38010] <= 16'b0000000000000101;
        weights1[38011] <= 16'b1111111111111101;
        weights1[38012] <= 16'b1111111111101011;
        weights1[38013] <= 16'b0000000000001001;
        weights1[38014] <= 16'b1111111111110100;
        weights1[38015] <= 16'b1111111111100110;
        weights1[38016] <= 16'b1111111111110111;
        weights1[38017] <= 16'b1111111111101100;
        weights1[38018] <= 16'b1111111111011100;
        weights1[38019] <= 16'b1111111111110100;
        weights1[38020] <= 16'b1111111111110011;
        weights1[38021] <= 16'b1111111111101111;
        weights1[38022] <= 16'b1111111111101110;
        weights1[38023] <= 16'b1111111111101000;
        weights1[38024] <= 16'b0000000000000001;
        weights1[38025] <= 16'b0000000000000101;
        weights1[38026] <= 16'b1111111111110110;
        weights1[38027] <= 16'b0000000000000100;
        weights1[38028] <= 16'b1111111111101110;
        weights1[38029] <= 16'b1111111111110011;
        weights1[38030] <= 16'b0000000000000011;
        weights1[38031] <= 16'b0000000000000010;
        weights1[38032] <= 16'b0000000000000010;
        weights1[38033] <= 16'b0000000000000100;
        weights1[38034] <= 16'b0000000000000010;
        weights1[38035] <= 16'b1111111111110100;
        weights1[38036] <= 16'b0000000000000001;
        weights1[38037] <= 16'b1111111111110110;
        weights1[38038] <= 16'b1111111111110010;
        weights1[38039] <= 16'b1111111111111011;
        weights1[38040] <= 16'b1111111111110100;
        weights1[38041] <= 16'b1111111111110111;
        weights1[38042] <= 16'b0000000000010110;
        weights1[38043] <= 16'b1111111111110100;
        weights1[38044] <= 16'b1111111111101001;
        weights1[38045] <= 16'b0000000000001010;
        weights1[38046] <= 16'b0000000000000011;
        weights1[38047] <= 16'b0000000000000011;
        weights1[38048] <= 16'b0000000000001101;
        weights1[38049] <= 16'b0000000000000000;
        weights1[38050] <= 16'b0000000000000010;
        weights1[38051] <= 16'b1111111111111010;
        weights1[38052] <= 16'b0000000000000000;
        weights1[38053] <= 16'b0000000000001001;
        weights1[38054] <= 16'b0000000000000111;
        weights1[38055] <= 16'b0000000000000011;
        weights1[38056] <= 16'b0000000000000100;
        weights1[38057] <= 16'b0000000000001111;
        weights1[38058] <= 16'b0000000000000100;
        weights1[38059] <= 16'b0000000000000000;
        weights1[38060] <= 16'b1111111111111100;
        weights1[38061] <= 16'b1111111111101111;
        weights1[38062] <= 16'b0000000000000111;
        weights1[38063] <= 16'b1111111111101011;
        weights1[38064] <= 16'b1111111111110000;
        weights1[38065] <= 16'b1111111111100100;
        weights1[38066] <= 16'b0000000000000000;
        weights1[38067] <= 16'b1111111111110110;
        weights1[38068] <= 16'b1111111111110011;
        weights1[38069] <= 16'b0000000000001100;
        weights1[38070] <= 16'b1111111111101010;
        weights1[38071] <= 16'b0000000000001010;
        weights1[38072] <= 16'b1111111111111101;
        weights1[38073] <= 16'b1111111111111000;
        weights1[38074] <= 16'b1111111111101011;
        weights1[38075] <= 16'b0000000000010000;
        weights1[38076] <= 16'b0000000000001100;
        weights1[38077] <= 16'b0000000000011000;
        weights1[38078] <= 16'b0000000000001011;
        weights1[38079] <= 16'b0000000000001000;
        weights1[38080] <= 16'b0000000000000100;
        weights1[38081] <= 16'b0000000000000001;
        weights1[38082] <= 16'b0000000000000111;
        weights1[38083] <= 16'b1111111111101110;
        weights1[38084] <= 16'b1111111111111100;
        weights1[38085] <= 16'b0000000000010111;
        weights1[38086] <= 16'b0000000000000100;
        weights1[38087] <= 16'b1111111111110111;
        weights1[38088] <= 16'b0000000000000101;
        weights1[38089] <= 16'b0000000000001010;
        weights1[38090] <= 16'b1111111111111111;
        weights1[38091] <= 16'b0000000000000101;
        weights1[38092] <= 16'b1111111111110011;
        weights1[38093] <= 16'b1111111111111010;
        weights1[38094] <= 16'b1111111111111101;
        weights1[38095] <= 16'b1111111111111010;
        weights1[38096] <= 16'b1111111111110100;
        weights1[38097] <= 16'b0000000000000010;
        weights1[38098] <= 16'b1111111111110000;
        weights1[38099] <= 16'b0000000000001100;
        weights1[38100] <= 16'b1111111111111010;
        weights1[38101] <= 16'b0000000000000101;
        weights1[38102] <= 16'b0000000000010010;
        weights1[38103] <= 16'b0000000000010101;
        weights1[38104] <= 16'b0000000000111100;
        weights1[38105] <= 16'b0000000000100000;
        weights1[38106] <= 16'b0000000000001100;
        weights1[38107] <= 16'b0000000000000100;
        weights1[38108] <= 16'b0000000000000100;
        weights1[38109] <= 16'b1111111111111000;
        weights1[38110] <= 16'b0000000000000101;
        weights1[38111] <= 16'b1111111111111000;
        weights1[38112] <= 16'b0000000000000101;
        weights1[38113] <= 16'b0000000000010000;
        weights1[38114] <= 16'b0000000000000010;
        weights1[38115] <= 16'b1111111111100100;
        weights1[38116] <= 16'b1111111111111010;
        weights1[38117] <= 16'b1111111111100111;
        weights1[38118] <= 16'b0000000000000001;
        weights1[38119] <= 16'b1111111111111000;
        weights1[38120] <= 16'b1111111111110111;
        weights1[38121] <= 16'b1111111111111011;
        weights1[38122] <= 16'b1111111111011101;
        weights1[38123] <= 16'b1111111111110011;
        weights1[38124] <= 16'b1111111111010100;
        weights1[38125] <= 16'b1111111111100111;
        weights1[38126] <= 16'b1111111111111011;
        weights1[38127] <= 16'b0000000000000110;
        weights1[38128] <= 16'b1111111111111111;
        weights1[38129] <= 16'b0000000000011110;
        weights1[38130] <= 16'b0000000000101100;
        weights1[38131] <= 16'b0000000000001100;
        weights1[38132] <= 16'b0000000000011100;
        weights1[38133] <= 16'b0000000000110101;
        weights1[38134] <= 16'b0000000000100001;
        weights1[38135] <= 16'b0000000000001000;
        weights1[38136] <= 16'b0000000000001011;
        weights1[38137] <= 16'b1111111111111010;
        weights1[38138] <= 16'b0000000000000010;
        weights1[38139] <= 16'b1111111111111101;
        weights1[38140] <= 16'b1111111111111111;
        weights1[38141] <= 16'b1111111111110001;
        weights1[38142] <= 16'b1111111111011010;
        weights1[38143] <= 16'b0000000000000010;
        weights1[38144] <= 16'b0000000000001001;
        weights1[38145] <= 16'b1111111111101001;
        weights1[38146] <= 16'b1111111111110100;
        weights1[38147] <= 16'b1111111111101110;
        weights1[38148] <= 16'b1111111111110010;
        weights1[38149] <= 16'b1111111111101011;
        weights1[38150] <= 16'b1111111111100011;
        weights1[38151] <= 16'b1111111111101110;
        weights1[38152] <= 16'b0000000000000000;
        weights1[38153] <= 16'b0000000000000001;
        weights1[38154] <= 16'b0000000000000011;
        weights1[38155] <= 16'b0000000000101000;
        weights1[38156] <= 16'b0000000000010011;
        weights1[38157] <= 16'b0000000000100001;
        weights1[38158] <= 16'b0000000000011000;
        weights1[38159] <= 16'b0000000000100100;
        weights1[38160] <= 16'b0000000000100001;
        weights1[38161] <= 16'b0000000000110001;
        weights1[38162] <= 16'b0000000000010101;
        weights1[38163] <= 16'b0000000000000000;
        weights1[38164] <= 16'b0000000000011100;
        weights1[38165] <= 16'b0000000000010011;
        weights1[38166] <= 16'b0000000000000000;
        weights1[38167] <= 16'b0000000000001011;
        weights1[38168] <= 16'b0000000000000010;
        weights1[38169] <= 16'b0000000000000101;
        weights1[38170] <= 16'b1111111111101101;
        weights1[38171] <= 16'b1111111111100100;
        weights1[38172] <= 16'b1111111111110101;
        weights1[38173] <= 16'b1111111111100110;
        weights1[38174] <= 16'b1111111111111110;
        weights1[38175] <= 16'b1111111111111110;
        weights1[38176] <= 16'b1111111111111111;
        weights1[38177] <= 16'b0000000000001101;
        weights1[38178] <= 16'b0000000000010010;
        weights1[38179] <= 16'b0000000000010111;
        weights1[38180] <= 16'b0000000000011011;
        weights1[38181] <= 16'b0000000000100001;
        weights1[38182] <= 16'b0000000000011100;
        weights1[38183] <= 16'b1111111111110111;
        weights1[38184] <= 16'b0000000000110110;
        weights1[38185] <= 16'b0000000000100001;
        weights1[38186] <= 16'b0000000000011100;
        weights1[38187] <= 16'b0000000000100101;
        weights1[38188] <= 16'b0000000000100000;
        weights1[38189] <= 16'b0000000000001010;
        weights1[38190] <= 16'b0000000000000110;
        weights1[38191] <= 16'b1111111111111011;
        weights1[38192] <= 16'b0000000000101100;
        weights1[38193] <= 16'b0000000000011010;
        weights1[38194] <= 16'b0000000000011110;
        weights1[38195] <= 16'b0000000000101110;
        weights1[38196] <= 16'b0000000000011111;
        weights1[38197] <= 16'b0000000000011101;
        weights1[38198] <= 16'b0000000000001101;
        weights1[38199] <= 16'b0000000000001110;
        weights1[38200] <= 16'b0000000000011000;
        weights1[38201] <= 16'b0000000000011100;
        weights1[38202] <= 16'b0000000000010000;
        weights1[38203] <= 16'b0000000000010011;
        weights1[38204] <= 16'b0000000000101010;
        weights1[38205] <= 16'b0000000000100001;
        weights1[38206] <= 16'b0000000000111001;
        weights1[38207] <= 16'b0000000000110111;
        weights1[38208] <= 16'b0000000000101101;
        weights1[38209] <= 16'b0000000000101001;
        weights1[38210] <= 16'b0000000000100100;
        weights1[38211] <= 16'b0000000000110011;
        weights1[38212] <= 16'b0000000000011010;
        weights1[38213] <= 16'b0000000000011001;
        weights1[38214] <= 16'b0000000000010011;
        weights1[38215] <= 16'b0000000000010111;
        weights1[38216] <= 16'b0000000000010000;
        weights1[38217] <= 16'b1111111111110101;
        weights1[38218] <= 16'b1111111111101011;
        weights1[38219] <= 16'b1111111111011111;
        weights1[38220] <= 16'b0000000000101001;
        weights1[38221] <= 16'b0000000000101011;
        weights1[38222] <= 16'b0000000000011111;
        weights1[38223] <= 16'b0000000000110110;
        weights1[38224] <= 16'b0000000000100100;
        weights1[38225] <= 16'b0000000000011011;
        weights1[38226] <= 16'b0000000000011000;
        weights1[38227] <= 16'b0000000000110011;
        weights1[38228] <= 16'b0000000000011101;
        weights1[38229] <= 16'b0000000000110010;
        weights1[38230] <= 16'b0000000000110000;
        weights1[38231] <= 16'b0000000000100111;
        weights1[38232] <= 16'b0000000000110000;
        weights1[38233] <= 16'b0000000000111101;
        weights1[38234] <= 16'b0000000000010100;
        weights1[38235] <= 16'b0000000000100010;
        weights1[38236] <= 16'b0000000000100110;
        weights1[38237] <= 16'b0000000000001011;
        weights1[38238] <= 16'b0000000000100011;
        weights1[38239] <= 16'b0000000000100001;
        weights1[38240] <= 16'b0000000000011000;
        weights1[38241] <= 16'b0000000000100000;
        weights1[38242] <= 16'b0000000000010100;
        weights1[38243] <= 16'b1111111111111000;
        weights1[38244] <= 16'b1111111111110000;
        weights1[38245] <= 16'b1111111111001000;
        weights1[38246] <= 16'b1111111111001010;
        weights1[38247] <= 16'b1111111111011110;
        weights1[38248] <= 16'b0000000000010110;
        weights1[38249] <= 16'b0000000000010100;
        weights1[38250] <= 16'b0000000000010100;
        weights1[38251] <= 16'b0000000000101110;
        weights1[38252] <= 16'b0000000000100000;
        weights1[38253] <= 16'b0000000000110101;
        weights1[38254] <= 16'b0000000000110111;
        weights1[38255] <= 16'b0000000000000010;
        weights1[38256] <= 16'b0000000000011010;
        weights1[38257] <= 16'b0000000000011111;
        weights1[38258] <= 16'b1111111111111001;
        weights1[38259] <= 16'b0000000000011100;
        weights1[38260] <= 16'b0000000000011100;
        weights1[38261] <= 16'b0000000000001000;
        weights1[38262] <= 16'b0000000000000011;
        weights1[38263] <= 16'b0000000000101110;
        weights1[38264] <= 16'b0000000000011011;
        weights1[38265] <= 16'b0000000000011100;
        weights1[38266] <= 16'b0000000000011101;
        weights1[38267] <= 16'b0000000000110111;
        weights1[38268] <= 16'b0000000000001110;
        weights1[38269] <= 16'b0000000000011010;
        weights1[38270] <= 16'b1111111111011001;
        weights1[38271] <= 16'b1111111111100101;
        weights1[38272] <= 16'b1111111111010001;
        weights1[38273] <= 16'b1111111111001001;
        weights1[38274] <= 16'b1111111111001000;
        weights1[38275] <= 16'b1111111111010010;
        weights1[38276] <= 16'b0000000000010010;
        weights1[38277] <= 16'b0000000000000101;
        weights1[38278] <= 16'b0000000000001111;
        weights1[38279] <= 16'b0000000000010011;
        weights1[38280] <= 16'b0000000000010100;
        weights1[38281] <= 16'b0000000000011110;
        weights1[38282] <= 16'b0000000000100010;
        weights1[38283] <= 16'b0000000000010111;
        weights1[38284] <= 16'b0000000000011011;
        weights1[38285] <= 16'b0000000000010001;
        weights1[38286] <= 16'b0000000000011000;
        weights1[38287] <= 16'b0000000000010111;
        weights1[38288] <= 16'b0000000000100001;
        weights1[38289] <= 16'b0000000000011011;
        weights1[38290] <= 16'b0000000000011001;
        weights1[38291] <= 16'b0000000000011011;
        weights1[38292] <= 16'b0000000000000110;
        weights1[38293] <= 16'b1111111111110011;
        weights1[38294] <= 16'b0000000000000010;
        weights1[38295] <= 16'b1111111111111001;
        weights1[38296] <= 16'b1111111111101001;
        weights1[38297] <= 16'b1111111111001000;
        weights1[38298] <= 16'b1111111110100110;
        weights1[38299] <= 16'b1111111110110110;
        weights1[38300] <= 16'b1111111110110111;
        weights1[38301] <= 16'b1111111111001011;
        weights1[38302] <= 16'b1111111111000111;
        weights1[38303] <= 16'b1111111111011000;
        weights1[38304] <= 16'b0000000000000000;
        weights1[38305] <= 16'b1111111111111101;
        weights1[38306] <= 16'b1111111111111000;
        weights1[38307] <= 16'b1111111111100000;
        weights1[38308] <= 16'b0000000000000000;
        weights1[38309] <= 16'b1111111111111000;
        weights1[38310] <= 16'b1111111111111111;
        weights1[38311] <= 16'b0000000000000001;
        weights1[38312] <= 16'b0000000000001000;
        weights1[38313] <= 16'b0000000000001001;
        weights1[38314] <= 16'b1111111111101111;
        weights1[38315] <= 16'b1111111111110100;
        weights1[38316] <= 16'b1111111111111111;
        weights1[38317] <= 16'b1111111111101000;
        weights1[38318] <= 16'b0000000000001000;
        weights1[38319] <= 16'b1111111111010111;
        weights1[38320] <= 16'b1111111111101100;
        weights1[38321] <= 16'b1111111111101000;
        weights1[38322] <= 16'b1111111111010110;
        weights1[38323] <= 16'b1111111110001100;
        weights1[38324] <= 16'b1111111101101100;
        weights1[38325] <= 16'b1111111101111100;
        weights1[38326] <= 16'b1111111101111110;
        weights1[38327] <= 16'b1111111110011001;
        weights1[38328] <= 16'b1111111110110100;
        weights1[38329] <= 16'b1111111111001110;
        weights1[38330] <= 16'b1111111111011001;
        weights1[38331] <= 16'b1111111111011000;
        weights1[38332] <= 16'b1111111111111110;
        weights1[38333] <= 16'b1111111111110101;
        weights1[38334] <= 16'b1111111111100001;
        weights1[38335] <= 16'b1111111111010011;
        weights1[38336] <= 16'b1111111111000110;
        weights1[38337] <= 16'b1111111111001111;
        weights1[38338] <= 16'b1111111111010001;
        weights1[38339] <= 16'b1111111111011001;
        weights1[38340] <= 16'b1111111111011000;
        weights1[38341] <= 16'b1111111111010111;
        weights1[38342] <= 16'b1111111111010110;
        weights1[38343] <= 16'b1111111110111001;
        weights1[38344] <= 16'b1111111110101001;
        weights1[38345] <= 16'b1111111110101001;
        weights1[38346] <= 16'b1111111101101011;
        weights1[38347] <= 16'b1111111101110101;
        weights1[38348] <= 16'b1111111101011001;
        weights1[38349] <= 16'b1111111101010001;
        weights1[38350] <= 16'b1111111101001100;
        weights1[38351] <= 16'b1111111101101011;
        weights1[38352] <= 16'b1111111101110011;
        weights1[38353] <= 16'b1111111110000101;
        weights1[38354] <= 16'b1111111110011010;
        weights1[38355] <= 16'b1111111110101010;
        weights1[38356] <= 16'b1111111110110001;
        weights1[38357] <= 16'b1111111111010001;
        weights1[38358] <= 16'b1111111111011101;
        weights1[38359] <= 16'b1111111111100110;
        weights1[38360] <= 16'b1111111111111001;
        weights1[38361] <= 16'b1111111111110110;
        weights1[38362] <= 16'b1111111111011011;
        weights1[38363] <= 16'b1111111111010110;
        weights1[38364] <= 16'b1111111111001010;
        weights1[38365] <= 16'b1111111110110010;
        weights1[38366] <= 16'b1111111110101011;
        weights1[38367] <= 16'b1111111110100000;
        weights1[38368] <= 16'b1111111110010011;
        weights1[38369] <= 16'b1111111110000101;
        weights1[38370] <= 16'b1111111110000001;
        weights1[38371] <= 16'b1111111101101010;
        weights1[38372] <= 16'b1111111101110101;
        weights1[38373] <= 16'b1111111101101000;
        weights1[38374] <= 16'b1111111101110001;
        weights1[38375] <= 16'b1111111101101001;
        weights1[38376] <= 16'b1111111101101110;
        weights1[38377] <= 16'b1111111101110010;
        weights1[38378] <= 16'b1111111101111011;
        weights1[38379] <= 16'b1111111110000111;
        weights1[38380] <= 16'b1111111110100000;
        weights1[38381] <= 16'b1111111110110000;
        weights1[38382] <= 16'b1111111111000110;
        weights1[38383] <= 16'b1111111111000010;
        weights1[38384] <= 16'b1111111111000111;
        weights1[38385] <= 16'b1111111111011101;
        weights1[38386] <= 16'b1111111111100110;
        weights1[38387] <= 16'b1111111111110101;
        weights1[38388] <= 16'b1111111111111100;
        weights1[38389] <= 16'b1111111111111100;
        weights1[38390] <= 16'b1111111111110000;
        weights1[38391] <= 16'b1111111111101000;
        weights1[38392] <= 16'b1111111111011001;
        weights1[38393] <= 16'b1111111111001100;
        weights1[38394] <= 16'b1111111111001011;
        weights1[38395] <= 16'b1111111110111100;
        weights1[38396] <= 16'b1111111110111001;
        weights1[38397] <= 16'b1111111110101010;
        weights1[38398] <= 16'b1111111110100110;
        weights1[38399] <= 16'b1111111110100000;
        weights1[38400] <= 16'b1111111110100100;
        weights1[38401] <= 16'b1111111110100001;
        weights1[38402] <= 16'b1111111110011101;
        weights1[38403] <= 16'b1111111110100100;
        weights1[38404] <= 16'b1111111110011100;
        weights1[38405] <= 16'b1111111110100111;
        weights1[38406] <= 16'b1111111110101110;
        weights1[38407] <= 16'b1111111110110110;
        weights1[38408] <= 16'b1111111111000100;
        weights1[38409] <= 16'b1111111111001111;
        weights1[38410] <= 16'b1111111111011110;
        weights1[38411] <= 16'b1111111111100010;
        weights1[38412] <= 16'b1111111111011010;
        weights1[38413] <= 16'b1111111111101101;
        weights1[38414] <= 16'b1111111111110000;
        weights1[38415] <= 16'b1111111111111101;
        weights1[38416] <= 16'b0000000000000000;
        weights1[38417] <= 16'b0000000000000001;
        weights1[38418] <= 16'b0000000000000000;
        weights1[38419] <= 16'b0000000000000000;
        weights1[38420] <= 16'b1111111111111111;
        weights1[38421] <= 16'b1111111111111110;
        weights1[38422] <= 16'b1111111111111101;
        weights1[38423] <= 16'b1111111111111010;
        weights1[38424] <= 16'b1111111111111011;
        weights1[38425] <= 16'b1111111111111111;
        weights1[38426] <= 16'b1111111111111101;
        weights1[38427] <= 16'b1111111111111110;
        weights1[38428] <= 16'b1111111111111011;
        weights1[38429] <= 16'b1111111111110101;
        weights1[38430] <= 16'b1111111111110001;
        weights1[38431] <= 16'b1111111111111101;
        weights1[38432] <= 16'b1111111111111001;
        weights1[38433] <= 16'b0000000000001011;
        weights1[38434] <= 16'b0000000000000011;
        weights1[38435] <= 16'b1111111111111000;
        weights1[38436] <= 16'b1111111111110110;
        weights1[38437] <= 16'b1111111111111111;
        weights1[38438] <= 16'b1111111111111010;
        weights1[38439] <= 16'b1111111111111101;
        weights1[38440] <= 16'b1111111111111111;
        weights1[38441] <= 16'b0000000000000011;
        weights1[38442] <= 16'b0000000000000010;
        weights1[38443] <= 16'b0000000000000000;
        weights1[38444] <= 16'b0000000000000000;
        weights1[38445] <= 16'b0000000000000001;
        weights1[38446] <= 16'b0000000000000100;
        weights1[38447] <= 16'b0000000000000110;
        weights1[38448] <= 16'b0000000000000010;
        weights1[38449] <= 16'b0000000000000111;
        weights1[38450] <= 16'b0000000000001010;
        weights1[38451] <= 16'b0000000000000110;
        weights1[38452] <= 16'b0000000000001001;
        weights1[38453] <= 16'b0000000000001100;
        weights1[38454] <= 16'b0000000000000000;
        weights1[38455] <= 16'b1111111111101001;
        weights1[38456] <= 16'b1111111111110101;
        weights1[38457] <= 16'b1111111111110111;
        weights1[38458] <= 16'b1111111111100111;
        weights1[38459] <= 16'b0000000000001101;
        weights1[38460] <= 16'b0000000000001110;
        weights1[38461] <= 16'b0000000000001011;
        weights1[38462] <= 16'b1111111111111111;
        weights1[38463] <= 16'b1111111111111000;
        weights1[38464] <= 16'b1111111111111001;
        weights1[38465] <= 16'b0000000000000001;
        weights1[38466] <= 16'b0000000000000000;
        weights1[38467] <= 16'b0000000000000100;
        weights1[38468] <= 16'b0000000000000010;
        weights1[38469] <= 16'b0000000000000011;
        weights1[38470] <= 16'b0000000000000001;
        weights1[38471] <= 16'b1111111111111111;
        weights1[38472] <= 16'b0000000000000000;
        weights1[38473] <= 16'b0000000000000010;
        weights1[38474] <= 16'b0000000000001010;
        weights1[38475] <= 16'b0000000000001100;
        weights1[38476] <= 16'b0000000000001110;
        weights1[38477] <= 16'b0000000000010001;
        weights1[38478] <= 16'b0000000000010001;
        weights1[38479] <= 16'b0000000000010101;
        weights1[38480] <= 16'b0000000000001000;
        weights1[38481] <= 16'b0000000000001011;
        weights1[38482] <= 16'b1111111111111110;
        weights1[38483] <= 16'b1111111111101110;
        weights1[38484] <= 16'b0000000000000010;
        weights1[38485] <= 16'b0000000000000000;
        weights1[38486] <= 16'b1111111111110100;
        weights1[38487] <= 16'b1111111111101110;
        weights1[38488] <= 16'b1111111111110001;
        weights1[38489] <= 16'b1111111111110000;
        weights1[38490] <= 16'b1111111111110110;
        weights1[38491] <= 16'b0000000000000001;
        weights1[38492] <= 16'b1111111111111101;
        weights1[38493] <= 16'b1111111111111101;
        weights1[38494] <= 16'b1111111111111101;
        weights1[38495] <= 16'b0000000000000011;
        weights1[38496] <= 16'b0000000000000010;
        weights1[38497] <= 16'b0000000000000101;
        weights1[38498] <= 16'b0000000000000101;
        weights1[38499] <= 16'b0000000000000100;
        weights1[38500] <= 16'b0000000000000001;
        weights1[38501] <= 16'b0000000000000100;
        weights1[38502] <= 16'b0000000000001110;
        weights1[38503] <= 16'b0000000000010100;
        weights1[38504] <= 16'b0000000000011100;
        weights1[38505] <= 16'b0000000000100001;
        weights1[38506] <= 16'b0000000000011001;
        weights1[38507] <= 16'b0000000000001010;
        weights1[38508] <= 16'b0000000000011001;
        weights1[38509] <= 16'b0000000000010110;
        weights1[38510] <= 16'b0000000000010000;
        weights1[38511] <= 16'b0000000000000000;
        weights1[38512] <= 16'b1111111111101111;
        weights1[38513] <= 16'b1111111111111111;
        weights1[38514] <= 16'b1111111111111101;
        weights1[38515] <= 16'b1111111111110100;
        weights1[38516] <= 16'b1111111111110100;
        weights1[38517] <= 16'b1111111111100111;
        weights1[38518] <= 16'b1111111111011000;
        weights1[38519] <= 16'b1111111111100101;
        weights1[38520] <= 16'b1111111111011010;
        weights1[38521] <= 16'b1111111111110101;
        weights1[38522] <= 16'b1111111111111011;
        weights1[38523] <= 16'b0000000000000000;
        weights1[38524] <= 16'b0000000000000100;
        weights1[38525] <= 16'b0000000000000011;
        weights1[38526] <= 16'b0000000000001000;
        weights1[38527] <= 16'b0000000000000011;
        weights1[38528] <= 16'b0000000000000110;
        weights1[38529] <= 16'b0000000000001000;
        weights1[38530] <= 16'b0000000000010011;
        weights1[38531] <= 16'b0000000000011110;
        weights1[38532] <= 16'b0000000000011011;
        weights1[38533] <= 16'b0000000000011000;
        weights1[38534] <= 16'b0000000000011101;
        weights1[38535] <= 16'b0000000000011000;
        weights1[38536] <= 16'b0000000000001000;
        weights1[38537] <= 16'b0000000000011001;
        weights1[38538] <= 16'b1111111111111101;
        weights1[38539] <= 16'b0000000000001011;
        weights1[38540] <= 16'b1111111111110101;
        weights1[38541] <= 16'b1111111111111111;
        weights1[38542] <= 16'b1111111111111111;
        weights1[38543] <= 16'b1111111111111000;
        weights1[38544] <= 16'b0000000000010010;
        weights1[38545] <= 16'b0000000000000101;
        weights1[38546] <= 16'b0000000000010001;
        weights1[38547] <= 16'b1111111111111001;
        weights1[38548] <= 16'b1111111111110001;
        weights1[38549] <= 16'b1111111111101111;
        weights1[38550] <= 16'b1111111111111001;
        weights1[38551] <= 16'b0000000000000001;
        weights1[38552] <= 16'b0000000000001010;
        weights1[38553] <= 16'b0000000000000100;
        weights1[38554] <= 16'b0000000000001011;
        weights1[38555] <= 16'b0000000000001101;
        weights1[38556] <= 16'b0000000000000111;
        weights1[38557] <= 16'b0000000000010001;
        weights1[38558] <= 16'b0000000000010001;
        weights1[38559] <= 16'b0000000000011010;
        weights1[38560] <= 16'b0000000000010011;
        weights1[38561] <= 16'b0000000000001001;
        weights1[38562] <= 16'b0000000000001110;
        weights1[38563] <= 16'b0000000000010100;
        weights1[38564] <= 16'b0000000000000011;
        weights1[38565] <= 16'b0000000000010000;
        weights1[38566] <= 16'b1111111111111110;
        weights1[38567] <= 16'b0000000000001001;
        weights1[38568] <= 16'b1111111111101100;
        weights1[38569] <= 16'b0000000000001011;
        weights1[38570] <= 16'b1111111111100101;
        weights1[38571] <= 16'b1111111111110111;
        weights1[38572] <= 16'b1111111111110010;
        weights1[38573] <= 16'b1111111111110101;
        weights1[38574] <= 16'b1111111111111010;
        weights1[38575] <= 16'b1111111111111110;
        weights1[38576] <= 16'b1111111111110110;
        weights1[38577] <= 16'b0000000000000010;
        weights1[38578] <= 16'b0000000000001001;
        weights1[38579] <= 16'b0000000000000111;
        weights1[38580] <= 16'b0000000000001010;
        weights1[38581] <= 16'b0000000000000001;
        weights1[38582] <= 16'b0000000000001101;
        weights1[38583] <= 16'b0000000000000100;
        weights1[38584] <= 16'b0000000000001001;
        weights1[38585] <= 16'b0000000000001111;
        weights1[38586] <= 16'b0000000000010011;
        weights1[38587] <= 16'b0000000000010100;
        weights1[38588] <= 16'b0000000000001010;
        weights1[38589] <= 16'b0000000000010010;
        weights1[38590] <= 16'b1111111111111110;
        weights1[38591] <= 16'b0000000000010100;
        weights1[38592] <= 16'b1111111111111001;
        weights1[38593] <= 16'b1111111111111001;
        weights1[38594] <= 16'b0000000000001000;
        weights1[38595] <= 16'b1111111111111010;
        weights1[38596] <= 16'b1111111111110101;
        weights1[38597] <= 16'b1111111111110001;
        weights1[38598] <= 16'b0000000000000000;
        weights1[38599] <= 16'b1111111111110110;
        weights1[38600] <= 16'b1111111111111010;
        weights1[38601] <= 16'b0000000000000101;
        weights1[38602] <= 16'b0000000000001101;
        weights1[38603] <= 16'b1111111111101010;
        weights1[38604] <= 16'b0000000000011100;
        weights1[38605] <= 16'b0000000000011101;
        weights1[38606] <= 16'b0000000000000110;
        weights1[38607] <= 16'b0000000000000110;
        weights1[38608] <= 16'b0000000000001001;
        weights1[38609] <= 16'b0000000000001110;
        weights1[38610] <= 16'b0000000000001101;
        weights1[38611] <= 16'b1111111111111101;
        weights1[38612] <= 16'b0000000000001010;
        weights1[38613] <= 16'b0000000000010001;
        weights1[38614] <= 16'b0000000000001000;
        weights1[38615] <= 16'b0000000000001000;
        weights1[38616] <= 16'b0000000000000011;
        weights1[38617] <= 16'b0000000000000000;
        weights1[38618] <= 16'b1111111111111110;
        weights1[38619] <= 16'b1111111111111111;
        weights1[38620] <= 16'b0000000000000101;
        weights1[38621] <= 16'b0000000000000100;
        weights1[38622] <= 16'b1111111111110101;
        weights1[38623] <= 16'b1111111111111001;
        weights1[38624] <= 16'b1111111111101010;
        weights1[38625] <= 16'b0000000000010000;
        weights1[38626] <= 16'b1111111111111011;
        weights1[38627] <= 16'b1111111111110101;
        weights1[38628] <= 16'b0000000000001111;
        weights1[38629] <= 16'b0000000000000101;
        weights1[38630] <= 16'b0000000000000010;
        weights1[38631] <= 16'b0000000000001011;
        weights1[38632] <= 16'b0000000000011010;
        weights1[38633] <= 16'b0000000000000010;
        weights1[38634] <= 16'b0000000000001010;
        weights1[38635] <= 16'b1111111111111010;
        weights1[38636] <= 16'b1111111111110100;
        weights1[38637] <= 16'b1111111111101111;
        weights1[38638] <= 16'b0000000000001100;
        weights1[38639] <= 16'b1111111111110101;
        weights1[38640] <= 16'b0000000000001000;
        weights1[38641] <= 16'b0000000000000111;
        weights1[38642] <= 16'b0000000000000101;
        weights1[38643] <= 16'b0000000000001001;
        weights1[38644] <= 16'b0000000000000001;
        weights1[38645] <= 16'b0000000000001100;
        weights1[38646] <= 16'b1111111111111110;
        weights1[38647] <= 16'b1111111111111010;
        weights1[38648] <= 16'b1111111111101111;
        weights1[38649] <= 16'b1111111111100010;
        weights1[38650] <= 16'b1111111111010101;
        weights1[38651] <= 16'b1111111111101111;
        weights1[38652] <= 16'b1111111111111001;
        weights1[38653] <= 16'b1111111111111000;
        weights1[38654] <= 16'b1111111111110010;
        weights1[38655] <= 16'b0000000000100000;
        weights1[38656] <= 16'b1111111111110010;
        weights1[38657] <= 16'b0000000000001111;
        weights1[38658] <= 16'b1111111111110111;
        weights1[38659] <= 16'b0000000000000100;
        weights1[38660] <= 16'b1111111111111001;
        weights1[38661] <= 16'b1111111111111110;
        weights1[38662] <= 16'b0000000000011011;
        weights1[38663] <= 16'b1111111111111101;
        weights1[38664] <= 16'b1111111111010110;
        weights1[38665] <= 16'b0000000000001000;
        weights1[38666] <= 16'b1111111111111000;
        weights1[38667] <= 16'b1111111111110001;
        weights1[38668] <= 16'b0000000000000011;
        weights1[38669] <= 16'b0000000000000100;
        weights1[38670] <= 16'b0000000000000011;
        weights1[38671] <= 16'b0000000000000001;
        weights1[38672] <= 16'b1111111111110111;
        weights1[38673] <= 16'b1111111111110100;
        weights1[38674] <= 16'b1111111111110001;
        weights1[38675] <= 16'b1111111111100011;
        weights1[38676] <= 16'b1111111111001001;
        weights1[38677] <= 16'b1111111111000111;
        weights1[38678] <= 16'b1111111111000000;
        weights1[38679] <= 16'b1111111111100111;
        weights1[38680] <= 16'b1111111111101000;
        weights1[38681] <= 16'b1111111111101010;
        weights1[38682] <= 16'b0000000000000001;
        weights1[38683] <= 16'b0000000000000101;
        weights1[38684] <= 16'b0000000000001011;
        weights1[38685] <= 16'b0000000000000111;
        weights1[38686] <= 16'b0000000000000111;
        weights1[38687] <= 16'b0000000000000010;
        weights1[38688] <= 16'b1111111111111100;
        weights1[38689] <= 16'b0000000000000101;
        weights1[38690] <= 16'b1111111111111011;
        weights1[38691] <= 16'b1111111111100001;
        weights1[38692] <= 16'b0000000000001001;
        weights1[38693] <= 16'b1111111111111011;
        weights1[38694] <= 16'b1111111111111001;
        weights1[38695] <= 16'b1111111111111101;
        weights1[38696] <= 16'b0000000000000100;
        weights1[38697] <= 16'b1111111111111110;
        weights1[38698] <= 16'b0000000000000010;
        weights1[38699] <= 16'b0000000000000001;
        weights1[38700] <= 16'b1111111111111111;
        weights1[38701] <= 16'b1111111111110001;
        weights1[38702] <= 16'b1111111111101001;
        weights1[38703] <= 16'b1111111111001000;
        weights1[38704] <= 16'b1111111110110101;
        weights1[38705] <= 16'b1111111111001011;
        weights1[38706] <= 16'b1111111111000001;
        weights1[38707] <= 16'b1111111111101011;
        weights1[38708] <= 16'b1111111111100110;
        weights1[38709] <= 16'b1111111111101111;
        weights1[38710] <= 16'b0000000000000111;
        weights1[38711] <= 16'b0000000000001001;
        weights1[38712] <= 16'b1111111111110101;
        weights1[38713] <= 16'b1111111111111001;
        weights1[38714] <= 16'b0000000000000011;
        weights1[38715] <= 16'b0000000000000110;
        weights1[38716] <= 16'b0000000000010000;
        weights1[38717] <= 16'b0000000000001100;
        weights1[38718] <= 16'b1111111111111101;
        weights1[38719] <= 16'b0000000000000100;
        weights1[38720] <= 16'b1111111111111011;
        weights1[38721] <= 16'b0000000000000101;
        weights1[38722] <= 16'b0000000000001100;
        weights1[38723] <= 16'b0000000000001001;
        weights1[38724] <= 16'b0000000000000101;
        weights1[38725] <= 16'b1111111111111111;
        weights1[38726] <= 16'b0000000000000011;
        weights1[38727] <= 16'b1111111111111101;
        weights1[38728] <= 16'b1111111111110101;
        weights1[38729] <= 16'b1111111111101011;
        weights1[38730] <= 16'b1111111111011011;
        weights1[38731] <= 16'b1111111111010001;
        weights1[38732] <= 16'b1111111111000101;
        weights1[38733] <= 16'b1111111111001111;
        weights1[38734] <= 16'b1111111111100001;
        weights1[38735] <= 16'b0000000000000001;
        weights1[38736] <= 16'b0000000000001000;
        weights1[38737] <= 16'b0000000000000101;
        weights1[38738] <= 16'b0000000000000101;
        weights1[38739] <= 16'b0000000000000101;
        weights1[38740] <= 16'b0000000000000111;
        weights1[38741] <= 16'b1111111111101100;
        weights1[38742] <= 16'b0000000000000101;
        weights1[38743] <= 16'b1111111111110101;
        weights1[38744] <= 16'b1111111111110111;
        weights1[38745] <= 16'b0000000000001101;
        weights1[38746] <= 16'b0000000000001100;
        weights1[38747] <= 16'b0000000000011011;
        weights1[38748] <= 16'b0000000000000110;
        weights1[38749] <= 16'b0000000000001001;
        weights1[38750] <= 16'b0000000000011001;
        weights1[38751] <= 16'b0000000000001000;
        weights1[38752] <= 16'b0000000000000000;
        weights1[38753] <= 16'b1111111111111100;
        weights1[38754] <= 16'b0000000000000000;
        weights1[38755] <= 16'b1111111111110001;
        weights1[38756] <= 16'b1111111111011111;
        weights1[38757] <= 16'b1111111111010101;
        weights1[38758] <= 16'b1111111111001000;
        weights1[38759] <= 16'b1111111110110110;
        weights1[38760] <= 16'b1111111111000001;
        weights1[38761] <= 16'b1111111111010100;
        weights1[38762] <= 16'b1111111111110100;
        weights1[38763] <= 16'b1111111111111011;
        weights1[38764] <= 16'b0000000000000101;
        weights1[38765] <= 16'b1111111111111011;
        weights1[38766] <= 16'b0000000000001101;
        weights1[38767] <= 16'b0000000000001111;
        weights1[38768] <= 16'b1111111111110110;
        weights1[38769] <= 16'b1111111111101100;
        weights1[38770] <= 16'b0000000000001000;
        weights1[38771] <= 16'b0000000000000110;
        weights1[38772] <= 16'b0000000000010000;
        weights1[38773] <= 16'b0000000000100010;
        weights1[38774] <= 16'b0000000000001000;
        weights1[38775] <= 16'b0000000000010000;
        weights1[38776] <= 16'b0000000000000010;
        weights1[38777] <= 16'b1111111111111010;
        weights1[38778] <= 16'b0000000000000011;
        weights1[38779] <= 16'b0000000000001101;
        weights1[38780] <= 16'b0000000000000000;
        weights1[38781] <= 16'b1111111111111101;
        weights1[38782] <= 16'b1111111111110000;
        weights1[38783] <= 16'b1111111111100100;
        weights1[38784] <= 16'b1111111111010010;
        weights1[38785] <= 16'b1111111111001001;
        weights1[38786] <= 16'b1111111111000000;
        weights1[38787] <= 16'b1111111111010100;
        weights1[38788] <= 16'b1111111111000011;
        weights1[38789] <= 16'b1111111111000100;
        weights1[38790] <= 16'b0000000000001000;
        weights1[38791] <= 16'b0000000000000011;
        weights1[38792] <= 16'b0000000000011000;
        weights1[38793] <= 16'b0000000000011001;
        weights1[38794] <= 16'b0000000000001111;
        weights1[38795] <= 16'b1111111111101000;
        weights1[38796] <= 16'b1111111111010110;
        weights1[38797] <= 16'b1111111111010100;
        weights1[38798] <= 16'b1111111111110001;
        weights1[38799] <= 16'b0000000000000010;
        weights1[38800] <= 16'b0000000000001111;
        weights1[38801] <= 16'b1111111111111110;
        weights1[38802] <= 16'b1111111111110010;
        weights1[38803] <= 16'b0000000000000110;
        weights1[38804] <= 16'b0000000000010101;
        weights1[38805] <= 16'b0000000000000001;
        weights1[38806] <= 16'b0000000000000100;
        weights1[38807] <= 16'b0000000000001001;
        weights1[38808] <= 16'b1111111111111100;
        weights1[38809] <= 16'b0000000000000001;
        weights1[38810] <= 16'b1111111111101001;
        weights1[38811] <= 16'b1111111111011101;
        weights1[38812] <= 16'b1111111111001111;
        weights1[38813] <= 16'b1111111111000101;
        weights1[38814] <= 16'b1111111111000101;
        weights1[38815] <= 16'b1111111111010011;
        weights1[38816] <= 16'b1111111111010001;
        weights1[38817] <= 16'b1111111111101111;
        weights1[38818] <= 16'b0000000000001110;
        weights1[38819] <= 16'b0000000000100001;
        weights1[38820] <= 16'b0000000000011011;
        weights1[38821] <= 16'b0000000000010111;
        weights1[38822] <= 16'b0000000000000111;
        weights1[38823] <= 16'b1111111111101100;
        weights1[38824] <= 16'b1111111110111001;
        weights1[38825] <= 16'b1111111110100101;
        weights1[38826] <= 16'b1111111111000100;
        weights1[38827] <= 16'b0000000000010010;
        weights1[38828] <= 16'b1111111111101110;
        weights1[38829] <= 16'b0000000000000010;
        weights1[38830] <= 16'b0000000000000101;
        weights1[38831] <= 16'b0000000000000011;
        weights1[38832] <= 16'b1111111111111001;
        weights1[38833] <= 16'b0000000000000101;
        weights1[38834] <= 16'b0000000000000011;
        weights1[38835] <= 16'b1111111111111101;
        weights1[38836] <= 16'b1111111111111000;
        weights1[38837] <= 16'b1111111111111010;
        weights1[38838] <= 16'b1111111111100101;
        weights1[38839] <= 16'b1111111111100010;
        weights1[38840] <= 16'b1111111111011010;
        weights1[38841] <= 16'b1111111111010100;
        weights1[38842] <= 16'b1111111111001100;
        weights1[38843] <= 16'b1111111111100000;
        weights1[38844] <= 16'b1111111111101110;
        weights1[38845] <= 16'b1111111111101011;
        weights1[38846] <= 16'b0000000000011011;
        weights1[38847] <= 16'b0000000000001111;
        weights1[38848] <= 16'b0000000000010111;
        weights1[38849] <= 16'b0000000000010101;
        weights1[38850] <= 16'b0000000000000110;
        weights1[38851] <= 16'b0000000000010001;
        weights1[38852] <= 16'b1111111110110000;
        weights1[38853] <= 16'b1111111101111111;
        weights1[38854] <= 16'b1111111111000101;
        weights1[38855] <= 16'b1111111111110010;
        weights1[38856] <= 16'b1111111111111010;
        weights1[38857] <= 16'b1111111111111111;
        weights1[38858] <= 16'b1111111111110110;
        weights1[38859] <= 16'b1111111111111100;
        weights1[38860] <= 16'b0000000000000010;
        weights1[38861] <= 16'b0000000000001101;
        weights1[38862] <= 16'b1111111111111110;
        weights1[38863] <= 16'b0000000000001010;
        weights1[38864] <= 16'b1111111111111010;
        weights1[38865] <= 16'b1111111111110011;
        weights1[38866] <= 16'b1111111111101110;
        weights1[38867] <= 16'b1111111111101011;
        weights1[38868] <= 16'b1111111111100000;
        weights1[38869] <= 16'b1111111111100111;
        weights1[38870] <= 16'b1111111111100000;
        weights1[38871] <= 16'b1111111111101111;
        weights1[38872] <= 16'b1111111111100011;
        weights1[38873] <= 16'b0000000000001010;
        weights1[38874] <= 16'b0000000000010100;
        weights1[38875] <= 16'b0000000000010000;
        weights1[38876] <= 16'b0000000000111101;
        weights1[38877] <= 16'b0000000000101010;
        weights1[38878] <= 16'b1111111111111111;
        weights1[38879] <= 16'b1111111111100101;
        weights1[38880] <= 16'b1111111101110100;
        weights1[38881] <= 16'b1111111101111101;
        weights1[38882] <= 16'b1111111111110110;
        weights1[38883] <= 16'b1111111111101100;
        weights1[38884] <= 16'b1111111111100100;
        weights1[38885] <= 16'b1111111111101100;
        weights1[38886] <= 16'b1111111111101111;
        weights1[38887] <= 16'b1111111111100111;
        weights1[38888] <= 16'b0000000000000001;
        weights1[38889] <= 16'b1111111111110001;
        weights1[38890] <= 16'b1111111111110110;
        weights1[38891] <= 16'b0000000000001001;
        weights1[38892] <= 16'b1111111111110110;
        weights1[38893] <= 16'b1111111111110001;
        weights1[38894] <= 16'b1111111111110011;
        weights1[38895] <= 16'b1111111111110101;
        weights1[38896] <= 16'b1111111111101101;
        weights1[38897] <= 16'b1111111111100000;
        weights1[38898] <= 16'b1111111111111111;
        weights1[38899] <= 16'b1111111111110011;
        weights1[38900] <= 16'b1111111111110100;
        weights1[38901] <= 16'b1111111111111000;
        weights1[38902] <= 16'b0000000000010111;
        weights1[38903] <= 16'b0000000000011011;
        weights1[38904] <= 16'b0000000000101001;
        weights1[38905] <= 16'b1111111111101111;
        weights1[38906] <= 16'b1111111111110111;
        weights1[38907] <= 16'b1111111110111001;
        weights1[38908] <= 16'b1111111101000110;
        weights1[38909] <= 16'b1111111110101100;
        weights1[38910] <= 16'b1111111111100010;
        weights1[38911] <= 16'b1111111111110010;
        weights1[38912] <= 16'b1111111111100111;
        weights1[38913] <= 16'b1111111111101000;
        weights1[38914] <= 16'b1111111111110011;
        weights1[38915] <= 16'b1111111111110011;
        weights1[38916] <= 16'b1111111111111100;
        weights1[38917] <= 16'b1111111111110100;
        weights1[38918] <= 16'b1111111111111000;
        weights1[38919] <= 16'b0000000000000000;
        weights1[38920] <= 16'b1111111111110001;
        weights1[38921] <= 16'b1111111111111110;
        weights1[38922] <= 16'b1111111111111011;
        weights1[38923] <= 16'b1111111111111001;
        weights1[38924] <= 16'b0000000000000110;
        weights1[38925] <= 16'b1111111111111011;
        weights1[38926] <= 16'b0000000000000111;
        weights1[38927] <= 16'b1111111111111011;
        weights1[38928] <= 16'b1111111111111011;
        weights1[38929] <= 16'b1111111111111111;
        weights1[38930] <= 16'b0000000000011100;
        weights1[38931] <= 16'b0000000000000101;
        weights1[38932] <= 16'b0000000000000110;
        weights1[38933] <= 16'b1111111111110010;
        weights1[38934] <= 16'b1111111111110101;
        weights1[38935] <= 16'b1111111101111010;
        weights1[38936] <= 16'b1111111101100111;
        weights1[38937] <= 16'b1111111111100011;
        weights1[38938] <= 16'b1111111111111010;
        weights1[38939] <= 16'b1111111111100011;
        weights1[38940] <= 16'b1111111111111010;
        weights1[38941] <= 16'b1111111111110100;
        weights1[38942] <= 16'b1111111111111000;
        weights1[38943] <= 16'b1111111111111100;
        weights1[38944] <= 16'b1111111111111001;
        weights1[38945] <= 16'b1111111111110111;
        weights1[38946] <= 16'b1111111111110101;
        weights1[38947] <= 16'b0000000000000010;
        weights1[38948] <= 16'b1111111111111010;
        weights1[38949] <= 16'b1111111111111101;
        weights1[38950] <= 16'b0000000000001000;
        weights1[38951] <= 16'b0000000000001000;
        weights1[38952] <= 16'b0000000000000000;
        weights1[38953] <= 16'b0000000000010010;
        weights1[38954] <= 16'b0000000000001100;
        weights1[38955] <= 16'b1111111111110101;
        weights1[38956] <= 16'b1111111111110101;
        weights1[38957] <= 16'b0000000000001101;
        weights1[38958] <= 16'b1111111111111010;
        weights1[38959] <= 16'b1111111111111101;
        weights1[38960] <= 16'b1111111111111100;
        weights1[38961] <= 16'b1111111111100001;
        weights1[38962] <= 16'b1111111111000010;
        weights1[38963] <= 16'b1111111101000000;
        weights1[38964] <= 16'b1111111110101011;
        weights1[38965] <= 16'b1111111111100111;
        weights1[38966] <= 16'b1111111111110101;
        weights1[38967] <= 16'b1111111111110001;
        weights1[38968] <= 16'b1111111111111010;
        weights1[38969] <= 16'b1111111111111010;
        weights1[38970] <= 16'b0000000000000000;
        weights1[38971] <= 16'b1111111111110011;
        weights1[38972] <= 16'b1111111111101110;
        weights1[38973] <= 16'b0000000000000011;
        weights1[38974] <= 16'b1111111111111011;
        weights1[38975] <= 16'b1111111111111100;
        weights1[38976] <= 16'b1111111111111111;
        weights1[38977] <= 16'b0000000000000111;
        weights1[38978] <= 16'b0000000000010011;
        weights1[38979] <= 16'b0000000000001011;
        weights1[38980] <= 16'b0000000000000111;
        weights1[38981] <= 16'b0000000000000101;
        weights1[38982] <= 16'b0000000000000010;
        weights1[38983] <= 16'b1111111111111010;
        weights1[38984] <= 16'b1111111111111000;
        weights1[38985] <= 16'b1111111111110111;
        weights1[38986] <= 16'b1111111111111100;
        weights1[38987] <= 16'b0000000000001111;
        weights1[38988] <= 16'b1111111111101010;
        weights1[38989] <= 16'b1111111111100001;
        weights1[38990] <= 16'b1111111110101011;
        weights1[38991] <= 16'b1111111110100000;
        weights1[38992] <= 16'b1111111111110000;
        weights1[38993] <= 16'b0000000000000110;
        weights1[38994] <= 16'b0000000000000001;
        weights1[38995] <= 16'b0000000000001110;
        weights1[38996] <= 16'b0000000000000010;
        weights1[38997] <= 16'b1111111111110011;
        weights1[38998] <= 16'b0000000000000101;
        weights1[38999] <= 16'b1111111111111000;
        weights1[39000] <= 16'b1111111111110111;
        weights1[39001] <= 16'b1111111111111101;
        weights1[39002] <= 16'b1111111111111010;
        weights1[39003] <= 16'b0000000000000101;
        weights1[39004] <= 16'b0000000000000100;
        weights1[39005] <= 16'b0000000000000001;
        weights1[39006] <= 16'b0000000000010011;
        weights1[39007] <= 16'b0000000000010010;
        weights1[39008] <= 16'b0000000000010000;
        weights1[39009] <= 16'b1111111111100011;
        weights1[39010] <= 16'b1111111111110101;
        weights1[39011] <= 16'b1111111111110101;
        weights1[39012] <= 16'b0000000000011001;
        weights1[39013] <= 16'b1111111111111100;
        weights1[39014] <= 16'b1111111111111001;
        weights1[39015] <= 16'b1111111111101111;
        weights1[39016] <= 16'b1111111111111101;
        weights1[39017] <= 16'b1111111111011100;
        weights1[39018] <= 16'b1111111111101001;
        weights1[39019] <= 16'b1111111111101111;
        weights1[39020] <= 16'b0000000000000010;
        weights1[39021] <= 16'b0000000000000011;
        weights1[39022] <= 16'b1111111111111101;
        weights1[39023] <= 16'b0000000000000110;
        weights1[39024] <= 16'b0000000000001101;
        weights1[39025] <= 16'b0000000000001010;
        weights1[39026] <= 16'b0000000000000110;
        weights1[39027] <= 16'b1111111111110101;
        weights1[39028] <= 16'b0000000000000000;
        weights1[39029] <= 16'b1111111111111111;
        weights1[39030] <= 16'b0000000000000001;
        weights1[39031] <= 16'b0000000000001000;
        weights1[39032] <= 16'b0000000000000111;
        weights1[39033] <= 16'b0000000000000110;
        weights1[39034] <= 16'b0000000000010001;
        weights1[39035] <= 16'b0000000000000010;
        weights1[39036] <= 16'b0000000000000110;
        weights1[39037] <= 16'b1111111111110100;
        weights1[39038] <= 16'b0000000000000111;
        weights1[39039] <= 16'b1111111111110010;
        weights1[39040] <= 16'b0000000000001110;
        weights1[39041] <= 16'b1111111111111001;
        weights1[39042] <= 16'b1111111111111111;
        weights1[39043] <= 16'b1111111111110100;
        weights1[39044] <= 16'b0000000000000100;
        weights1[39045] <= 16'b0000000000001101;
        weights1[39046] <= 16'b0000000000010011;
        weights1[39047] <= 16'b1111111111110010;
        weights1[39048] <= 16'b0000000000000001;
        weights1[39049] <= 16'b1111111111111101;
        weights1[39050] <= 16'b1111111111111000;
        weights1[39051] <= 16'b0000000000001000;
        weights1[39052] <= 16'b0000000000010001;
        weights1[39053] <= 16'b1111111111111100;
        weights1[39054] <= 16'b1111111111111001;
        weights1[39055] <= 16'b0000000000000011;
        weights1[39056] <= 16'b0000000000000100;
        weights1[39057] <= 16'b0000000000001000;
        weights1[39058] <= 16'b0000000000001010;
        weights1[39059] <= 16'b0000000000001011;
        weights1[39060] <= 16'b0000000000000011;
        weights1[39061] <= 16'b0000000000001110;
        weights1[39062] <= 16'b0000000000000011;
        weights1[39063] <= 16'b0000000000000001;
        weights1[39064] <= 16'b0000000000010010;
        weights1[39065] <= 16'b0000000000010110;
        weights1[39066] <= 16'b0000000000000001;
        weights1[39067] <= 16'b0000000000010010;
        weights1[39068] <= 16'b1111111111111001;
        weights1[39069] <= 16'b0000000000000000;
        weights1[39070] <= 16'b1111111111100100;
        weights1[39071] <= 16'b0000000000000010;
        weights1[39072] <= 16'b1111111111110000;
        weights1[39073] <= 16'b0000000000011110;
        weights1[39074] <= 16'b0000000000011000;
        weights1[39075] <= 16'b0000000000011110;
        weights1[39076] <= 16'b1111111111111111;
        weights1[39077] <= 16'b0000000000001100;
        weights1[39078] <= 16'b0000000000001000;
        weights1[39079] <= 16'b1111111111111000;
        weights1[39080] <= 16'b0000000000010100;
        weights1[39081] <= 16'b0000000000001000;
        weights1[39082] <= 16'b0000000000000110;
        weights1[39083] <= 16'b0000000000010010;
        weights1[39084] <= 16'b0000000000000100;
        weights1[39085] <= 16'b0000000000010010;
        weights1[39086] <= 16'b0000000000001111;
        weights1[39087] <= 16'b0000000000000110;
        weights1[39088] <= 16'b0000000000000010;
        weights1[39089] <= 16'b0000000000000111;
        weights1[39090] <= 16'b0000000000000100;
        weights1[39091] <= 16'b1111111111111010;
        weights1[39092] <= 16'b0000000000001001;
        weights1[39093] <= 16'b0000000000000101;
        weights1[39094] <= 16'b1111111111111111;
        weights1[39095] <= 16'b0000000000011010;
        weights1[39096] <= 16'b0000000000001100;
        weights1[39097] <= 16'b1111111111111111;
        weights1[39098] <= 16'b0000000000000110;
        weights1[39099] <= 16'b1111111111111010;
        weights1[39100] <= 16'b0000000000001110;
        weights1[39101] <= 16'b0000000000011000;
        weights1[39102] <= 16'b0000000000101101;
        weights1[39103] <= 16'b0000000000011111;
        weights1[39104] <= 16'b0000000000100001;
        weights1[39105] <= 16'b0000000000100010;
        weights1[39106] <= 16'b0000000000001110;
        weights1[39107] <= 16'b0000000000001011;
        weights1[39108] <= 16'b0000000000000000;
        weights1[39109] <= 16'b1111111111111001;
        weights1[39110] <= 16'b0000000000001011;
        weights1[39111] <= 16'b0000000000001111;
        weights1[39112] <= 16'b0000000000001110;
        weights1[39113] <= 16'b0000000000001110;
        weights1[39114] <= 16'b0000000000000011;
        weights1[39115] <= 16'b0000000000000000;
        weights1[39116] <= 16'b0000000000000110;
        weights1[39117] <= 16'b0000000000001011;
        weights1[39118] <= 16'b0000000000000111;
        weights1[39119] <= 16'b0000000000000100;
        weights1[39120] <= 16'b0000000000010101;
        weights1[39121] <= 16'b1111111111111110;
        weights1[39122] <= 16'b0000000000000100;
        weights1[39123] <= 16'b0000000000001011;
        weights1[39124] <= 16'b1111111111111100;
        weights1[39125] <= 16'b1111111111110111;
        weights1[39126] <= 16'b0000000000100010;
        weights1[39127] <= 16'b0000000000010111;
        weights1[39128] <= 16'b0000000000011101;
        weights1[39129] <= 16'b0000000000101101;
        weights1[39130] <= 16'b0000000000100010;
        weights1[39131] <= 16'b0000000000101101;
        weights1[39132] <= 16'b0000000000110000;
        weights1[39133] <= 16'b0000000000101100;
        weights1[39134] <= 16'b0000000000100101;
        weights1[39135] <= 16'b0000000000010100;
        weights1[39136] <= 16'b0000000000011000;
        weights1[39137] <= 16'b0000000000000101;
        weights1[39138] <= 16'b0000000000010100;
        weights1[39139] <= 16'b0000000000000001;
        weights1[39140] <= 16'b0000000000001110;
        weights1[39141] <= 16'b0000000000000110;
        weights1[39142] <= 16'b0000000000000001;
        weights1[39143] <= 16'b1111111111111110;
        weights1[39144] <= 16'b0000000000000101;
        weights1[39145] <= 16'b0000000000001011;
        weights1[39146] <= 16'b0000000000001011;
        weights1[39147] <= 16'b0000000000001000;
        weights1[39148] <= 16'b0000000000001100;
        weights1[39149] <= 16'b0000000000000110;
        weights1[39150] <= 16'b0000000000000111;
        weights1[39151] <= 16'b0000000000001011;
        weights1[39152] <= 16'b1111111111111110;
        weights1[39153] <= 16'b1111111111111000;
        weights1[39154] <= 16'b1111111111111110;
        weights1[39155] <= 16'b0000000000010001;
        weights1[39156] <= 16'b0000000000010001;
        weights1[39157] <= 16'b0000000000011000;
        weights1[39158] <= 16'b0000000000010010;
        weights1[39159] <= 16'b0000000000010111;
        weights1[39160] <= 16'b0000000000101000;
        weights1[39161] <= 16'b0000000000011010;
        weights1[39162] <= 16'b0000000000011100;
        weights1[39163] <= 16'b0000000000001110;
        weights1[39164] <= 16'b0000000000010110;
        weights1[39165] <= 16'b0000000000000101;
        weights1[39166] <= 16'b0000000000010110;
        weights1[39167] <= 16'b0000000000000001;
        weights1[39168] <= 16'b0000000000000010;
        weights1[39169] <= 16'b1111111111111001;
        weights1[39170] <= 16'b1111111111111101;
        weights1[39171] <= 16'b1111111111111101;
        weights1[39172] <= 16'b0000000000000000;
        weights1[39173] <= 16'b0000000000000110;
        weights1[39174] <= 16'b0000000000001000;
        weights1[39175] <= 16'b0000000000001011;
        weights1[39176] <= 16'b0000000000000101;
        weights1[39177] <= 16'b0000000000000101;
        weights1[39178] <= 16'b1111111111111111;
        weights1[39179] <= 16'b1111111111111001;
        weights1[39180] <= 16'b0000000000000000;
        weights1[39181] <= 16'b1111111111111101;
        weights1[39182] <= 16'b0000000000000010;
        weights1[39183] <= 16'b0000000000010101;
        weights1[39184] <= 16'b0000000000100001;
        weights1[39185] <= 16'b0000000000011101;
        weights1[39186] <= 16'b0000000000100000;
        weights1[39187] <= 16'b0000000000010000;
        weights1[39188] <= 16'b0000000000010110;
        weights1[39189] <= 16'b0000000000011111;
        weights1[39190] <= 16'b0000000000001111;
        weights1[39191] <= 16'b0000000000001110;
        weights1[39192] <= 16'b0000000000011001;
        weights1[39193] <= 16'b0000000000001010;
        weights1[39194] <= 16'b0000000000001001;
        weights1[39195] <= 16'b1111111111110010;
        weights1[39196] <= 16'b1111111111111000;
        weights1[39197] <= 16'b1111111111110101;
        weights1[39198] <= 16'b1111111111111010;
        weights1[39199] <= 16'b1111111111111110;
        weights1[39200] <= 16'b0000000000000001;
        weights1[39201] <= 16'b0000000000000001;
        weights1[39202] <= 16'b0000000000000001;
        weights1[39203] <= 16'b1111111111111111;
        weights1[39204] <= 16'b1111111111111010;
        weights1[39205] <= 16'b1111111111101010;
        weights1[39206] <= 16'b1111111111100100;
        weights1[39207] <= 16'b1111111111101011;
        weights1[39208] <= 16'b1111111111100010;
        weights1[39209] <= 16'b1111111111011110;
        weights1[39210] <= 16'b1111111111011010;
        weights1[39211] <= 16'b1111111111101110;
        weights1[39212] <= 16'b1111111111110001;
        weights1[39213] <= 16'b1111111111100111;
        weights1[39214] <= 16'b0000000000000001;
        weights1[39215] <= 16'b1111111111111110;
        weights1[39216] <= 16'b0000000000000001;
        weights1[39217] <= 16'b0000000000010000;
        weights1[39218] <= 16'b0000000000010101;
        weights1[39219] <= 16'b0000000000100100;
        weights1[39220] <= 16'b0000000000100100;
        weights1[39221] <= 16'b0000000000100101;
        weights1[39222] <= 16'b0000000000001110;
        weights1[39223] <= 16'b0000000000100000;
        weights1[39224] <= 16'b0000000000011000;
        weights1[39225] <= 16'b0000000000011001;
        weights1[39226] <= 16'b0000000000001101;
        weights1[39227] <= 16'b0000000000000100;
        weights1[39228] <= 16'b0000000000000001;
        weights1[39229] <= 16'b0000000000000001;
        weights1[39230] <= 16'b0000000000000001;
        weights1[39231] <= 16'b1111111111111110;
        weights1[39232] <= 16'b1111111111110010;
        weights1[39233] <= 16'b1111111111101011;
        weights1[39234] <= 16'b1111111111100110;
        weights1[39235] <= 16'b1111111111101010;
        weights1[39236] <= 16'b1111111111100000;
        weights1[39237] <= 16'b1111111111011100;
        weights1[39238] <= 16'b1111111111100110;
        weights1[39239] <= 16'b1111111111111001;
        weights1[39240] <= 16'b1111111111111100;
        weights1[39241] <= 16'b1111111111110001;
        weights1[39242] <= 16'b0000000000000110;
        weights1[39243] <= 16'b1111111111111101;
        weights1[39244] <= 16'b1111111111111111;
        weights1[39245] <= 16'b0000000000001111;
        weights1[39246] <= 16'b0000000000011011;
        weights1[39247] <= 16'b0000000000011101;
        weights1[39248] <= 16'b0000000000011001;
        weights1[39249] <= 16'b0000000000100111;
        weights1[39250] <= 16'b0000000000100101;
        weights1[39251] <= 16'b0000000000100010;
        weights1[39252] <= 16'b0000000000101111;
        weights1[39253] <= 16'b0000000000100101;
        weights1[39254] <= 16'b0000000000011110;
        weights1[39255] <= 16'b0000000000001001;
        weights1[39256] <= 16'b1111111111111111;
        weights1[39257] <= 16'b0000000000000000;
        weights1[39258] <= 16'b1111111111111110;
        weights1[39259] <= 16'b1111111111111010;
        weights1[39260] <= 16'b1111111111101000;
        weights1[39261] <= 16'b1111111111110100;
        weights1[39262] <= 16'b1111111111110010;
        weights1[39263] <= 16'b1111111111110110;
        weights1[39264] <= 16'b1111111111100010;
        weights1[39265] <= 16'b0000000000001101;
        weights1[39266] <= 16'b0000000000001101;
        weights1[39267] <= 16'b0000000000001010;
        weights1[39268] <= 16'b0000000000000000;
        weights1[39269] <= 16'b0000000000001101;
        weights1[39270] <= 16'b0000000000010000;
        weights1[39271] <= 16'b0000000000011100;
        weights1[39272] <= 16'b0000000000010000;
        weights1[39273] <= 16'b0000000000011001;
        weights1[39274] <= 16'b0000000000011101;
        weights1[39275] <= 16'b0000000000011001;
        weights1[39276] <= 16'b0000000000011000;
        weights1[39277] <= 16'b0000000000100100;
        weights1[39278] <= 16'b0000000000101111;
        weights1[39279] <= 16'b0000000000010111;
        weights1[39280] <= 16'b0000000000100110;
        weights1[39281] <= 16'b0000000000100001;
        weights1[39282] <= 16'b0000000000011101;
        weights1[39283] <= 16'b0000000000010101;
        weights1[39284] <= 16'b1111111111111101;
        weights1[39285] <= 16'b1111111111111010;
        weights1[39286] <= 16'b1111111111110111;
        weights1[39287] <= 16'b1111111111101110;
        weights1[39288] <= 16'b1111111111101010;
        weights1[39289] <= 16'b1111111111110000;
        weights1[39290] <= 16'b1111111111101110;
        weights1[39291] <= 16'b1111111111110110;
        weights1[39292] <= 16'b1111111111111010;
        weights1[39293] <= 16'b0000000000000010;
        weights1[39294] <= 16'b0000000000010010;
        weights1[39295] <= 16'b0000000000000101;
        weights1[39296] <= 16'b0000000000001110;
        weights1[39297] <= 16'b0000000000011100;
        weights1[39298] <= 16'b1111111111110111;
        weights1[39299] <= 16'b0000000000011110;
        weights1[39300] <= 16'b0000000000011101;
        weights1[39301] <= 16'b0000000000001010;
        weights1[39302] <= 16'b0000000000011011;
        weights1[39303] <= 16'b0000000000010101;
        weights1[39304] <= 16'b0000000000100101;
        weights1[39305] <= 16'b0000000000011100;
        weights1[39306] <= 16'b0000000000100111;
        weights1[39307] <= 16'b0000000000100110;
        weights1[39308] <= 16'b0000000000101110;
        weights1[39309] <= 16'b0000000000011010;
        weights1[39310] <= 16'b0000000000011010;
        weights1[39311] <= 16'b0000000000001011;
        weights1[39312] <= 16'b1111111111111011;
        weights1[39313] <= 16'b1111111111110001;
        weights1[39314] <= 16'b1111111111110101;
        weights1[39315] <= 16'b1111111111110011;
        weights1[39316] <= 16'b1111111111100000;
        weights1[39317] <= 16'b0000000000000101;
        weights1[39318] <= 16'b0000000000000010;
        weights1[39319] <= 16'b0000000000001000;
        weights1[39320] <= 16'b1111111111110100;
        weights1[39321] <= 16'b0000000000000110;
        weights1[39322] <= 16'b0000000000100000;
        weights1[39323] <= 16'b0000000000010010;
        weights1[39324] <= 16'b0000000000001000;
        weights1[39325] <= 16'b0000000000001101;
        weights1[39326] <= 16'b0000000000100001;
        weights1[39327] <= 16'b0000000000101001;
        weights1[39328] <= 16'b0000000000001111;
        weights1[39329] <= 16'b0000000000010001;
        weights1[39330] <= 16'b0000000000010110;
        weights1[39331] <= 16'b0000000000010001;
        weights1[39332] <= 16'b0000000000110001;
        weights1[39333] <= 16'b0000000001000101;
        weights1[39334] <= 16'b0000000001001010;
        weights1[39335] <= 16'b0000000000111010;
        weights1[39336] <= 16'b0000000000110111;
        weights1[39337] <= 16'b0000000000010010;
        weights1[39338] <= 16'b1111111111111011;
        weights1[39339] <= 16'b1111111111110100;
        weights1[39340] <= 16'b1111111111111101;
        weights1[39341] <= 16'b1111111111101101;
        weights1[39342] <= 16'b1111111111101001;
        weights1[39343] <= 16'b1111111111101001;
        weights1[39344] <= 16'b1111111111110100;
        weights1[39345] <= 16'b1111111111111011;
        weights1[39346] <= 16'b1111111111111111;
        weights1[39347] <= 16'b1111111111111001;
        weights1[39348] <= 16'b0000000000000001;
        weights1[39349] <= 16'b0000000000000011;
        weights1[39350] <= 16'b0000000000000001;
        weights1[39351] <= 16'b0000000000001110;
        weights1[39352] <= 16'b0000000000001001;
        weights1[39353] <= 16'b0000000000011100;
        weights1[39354] <= 16'b0000000000001000;
        weights1[39355] <= 16'b0000000000010101;
        weights1[39356] <= 16'b0000000000010000;
        weights1[39357] <= 16'b0000000000111100;
        weights1[39358] <= 16'b0000000000101101;
        weights1[39359] <= 16'b0000000000110011;
        weights1[39360] <= 16'b0000000001011010;
        weights1[39361] <= 16'b0000000000111100;
        weights1[39362] <= 16'b0000000000101001;
        weights1[39363] <= 16'b0000000000010110;
        weights1[39364] <= 16'b0000000000001110;
        weights1[39365] <= 16'b1111111111100110;
        weights1[39366] <= 16'b1111111111010000;
        weights1[39367] <= 16'b1111111111011111;
        weights1[39368] <= 16'b1111111111111011;
        weights1[39369] <= 16'b1111111111110001;
        weights1[39370] <= 16'b0000000000000001;
        weights1[39371] <= 16'b1111111111101111;
        weights1[39372] <= 16'b1111111111111000;
        weights1[39373] <= 16'b1111111111111001;
        weights1[39374] <= 16'b0000000000000010;
        weights1[39375] <= 16'b1111111111111011;
        weights1[39376] <= 16'b0000000000001110;
        weights1[39377] <= 16'b0000000000011000;
        weights1[39378] <= 16'b0000000000001011;
        weights1[39379] <= 16'b0000000000001111;
        weights1[39380] <= 16'b0000000000010000;
        weights1[39381] <= 16'b0000000000000010;
        weights1[39382] <= 16'b0000000000011111;
        weights1[39383] <= 16'b0000000000100000;
        weights1[39384] <= 16'b0000000000111011;
        weights1[39385] <= 16'b0000000000100100;
        weights1[39386] <= 16'b0000000000110110;
        weights1[39387] <= 16'b0000000000111000;
        weights1[39388] <= 16'b1111111111110110;
        weights1[39389] <= 16'b1111111111100001;
        weights1[39390] <= 16'b1111111111001010;
        weights1[39391] <= 16'b1111111110011001;
        weights1[39392] <= 16'b1111111110100001;
        weights1[39393] <= 16'b1111111110011101;
        weights1[39394] <= 16'b1111111110101110;
        weights1[39395] <= 16'b1111111111000000;
        weights1[39396] <= 16'b1111111111111001;
        weights1[39397] <= 16'b1111111111110101;
        weights1[39398] <= 16'b1111111111110100;
        weights1[39399] <= 16'b1111111111111000;
        weights1[39400] <= 16'b0000000000000010;
        weights1[39401] <= 16'b0000000000000110;
        weights1[39402] <= 16'b0000000000001111;
        weights1[39403] <= 16'b0000000000000010;
        weights1[39404] <= 16'b0000000000000001;
        weights1[39405] <= 16'b0000000000000010;
        weights1[39406] <= 16'b0000000000010001;
        weights1[39407] <= 16'b0000000000001010;
        weights1[39408] <= 16'b0000000000010101;
        weights1[39409] <= 16'b1111111111110111;
        weights1[39410] <= 16'b0000000000000010;
        weights1[39411] <= 16'b1111111111111001;
        weights1[39412] <= 16'b1111111111100110;
        weights1[39413] <= 16'b1111111110111110;
        weights1[39414] <= 16'b1111111110001001;
        weights1[39415] <= 16'b1111111101011010;
        weights1[39416] <= 16'b1111111101001111;
        weights1[39417] <= 16'b1111111101001011;
        weights1[39418] <= 16'b1111111101000010;
        weights1[39419] <= 16'b1111111101100011;
        weights1[39420] <= 16'b1111111101111010;
        weights1[39421] <= 16'b1111111110001000;
        weights1[39422] <= 16'b1111111110010111;
        weights1[39423] <= 16'b1111111110011110;
        weights1[39424] <= 16'b1111111111110100;
        weights1[39425] <= 16'b1111111111110010;
        weights1[39426] <= 16'b1111111111111010;
        weights1[39427] <= 16'b1111111111111100;
        weights1[39428] <= 16'b1111111111111100;
        weights1[39429] <= 16'b0000000000000001;
        weights1[39430] <= 16'b0000000000000100;
        weights1[39431] <= 16'b1111111111111100;
        weights1[39432] <= 16'b0000000000001101;
        weights1[39433] <= 16'b0000000000000001;
        weights1[39434] <= 16'b0000000000000100;
        weights1[39435] <= 16'b1111111111101110;
        weights1[39436] <= 16'b1111111111101110;
        weights1[39437] <= 16'b1111111111001100;
        weights1[39438] <= 16'b1111111110010111;
        weights1[39439] <= 16'b1111111101100111;
        weights1[39440] <= 16'b1111111100110011;
        weights1[39441] <= 16'b1111111011110010;
        weights1[39442] <= 16'b1111111011101110;
        weights1[39443] <= 16'b1111111011111101;
        weights1[39444] <= 16'b1111111100101011;
        weights1[39445] <= 16'b1111111100110011;
        weights1[39446] <= 16'b1111111101010101;
        weights1[39447] <= 16'b1111111101100011;
        weights1[39448] <= 16'b1111111101101100;
        weights1[39449] <= 16'b1111111110000000;
        weights1[39450] <= 16'b1111111110000010;
        weights1[39451] <= 16'b1111111110001101;
        weights1[39452] <= 16'b1111111111101111;
        weights1[39453] <= 16'b0000000000000100;
        weights1[39454] <= 16'b0000000000001100;
        weights1[39455] <= 16'b1111111111111111;
        weights1[39456] <= 16'b0000000000001111;
        weights1[39457] <= 16'b0000000000001000;
        weights1[39458] <= 16'b0000000000001010;
        weights1[39459] <= 16'b1111111111111110;
        weights1[39460] <= 16'b0000000000000011;
        weights1[39461] <= 16'b1111111111111011;
        weights1[39462] <= 16'b1111111111111010;
        weights1[39463] <= 16'b1111111111110001;
        weights1[39464] <= 16'b1111111111110001;
        weights1[39465] <= 16'b1111111111010110;
        weights1[39466] <= 16'b1111111111011111;
        weights1[39467] <= 16'b1111111111101000;
        weights1[39468] <= 16'b1111111111100100;
        weights1[39469] <= 16'b1111111111011011;
        weights1[39470] <= 16'b1111111111000010;
        weights1[39471] <= 16'b1111111110101001;
        weights1[39472] <= 16'b1111111110000010;
        weights1[39473] <= 16'b1111111101010101;
        weights1[39474] <= 16'b1111111101011100;
        weights1[39475] <= 16'b1111111101100011;
        weights1[39476] <= 16'b1111111101110100;
        weights1[39477] <= 16'b1111111110000001;
        weights1[39478] <= 16'b1111111110100101;
        weights1[39479] <= 16'b1111111110100110;
        weights1[39480] <= 16'b1111111111110000;
        weights1[39481] <= 16'b1111111111111110;
        weights1[39482] <= 16'b0000000000000011;
        weights1[39483] <= 16'b0000000000001101;
        weights1[39484] <= 16'b1111111111111101;
        weights1[39485] <= 16'b0000000000000001;
        weights1[39486] <= 16'b1111111111111100;
        weights1[39487] <= 16'b0000000000000000;
        weights1[39488] <= 16'b0000000000000001;
        weights1[39489] <= 16'b0000000000000001;
        weights1[39490] <= 16'b1111111111111011;
        weights1[39491] <= 16'b1111111111110001;
        weights1[39492] <= 16'b1111111111111110;
        weights1[39493] <= 16'b1111111111110011;
        weights1[39494] <= 16'b0000000000000010;
        weights1[39495] <= 16'b0000000000000000;
        weights1[39496] <= 16'b1111111111111001;
        weights1[39497] <= 16'b0000000000001000;
        weights1[39498] <= 16'b1111111111110010;
        weights1[39499] <= 16'b1111111111111100;
        weights1[39500] <= 16'b1111111111100111;
        weights1[39501] <= 16'b1111111111101111;
        weights1[39502] <= 16'b1111111111011101;
        weights1[39503] <= 16'b1111111111011100;
        weights1[39504] <= 16'b1111111111001011;
        weights1[39505] <= 16'b1111111111101011;
        weights1[39506] <= 16'b1111111111010100;
        weights1[39507] <= 16'b1111111111001001;
        weights1[39508] <= 16'b1111111111110101;
        weights1[39509] <= 16'b1111111111111100;
        weights1[39510] <= 16'b0000000000001000;
        weights1[39511] <= 16'b0000000000001001;
        weights1[39512] <= 16'b0000000000000011;
        weights1[39513] <= 16'b0000000000001001;
        weights1[39514] <= 16'b0000000000000000;
        weights1[39515] <= 16'b0000000000000011;
        weights1[39516] <= 16'b1111111111111010;
        weights1[39517] <= 16'b0000000000000110;
        weights1[39518] <= 16'b1111111111111000;
        weights1[39519] <= 16'b0000000000000101;
        weights1[39520] <= 16'b0000000000000000;
        weights1[39521] <= 16'b0000000000000001;
        weights1[39522] <= 16'b1111111111111010;
        weights1[39523] <= 16'b1111111111110001;
        weights1[39524] <= 16'b0000000000010001;
        weights1[39525] <= 16'b0000000000001010;
        weights1[39526] <= 16'b0000000000010001;
        weights1[39527] <= 16'b0000000000011001;
        weights1[39528] <= 16'b0000000000100011;
        weights1[39529] <= 16'b0000000000000110;
        weights1[39530] <= 16'b0000000000010100;
        weights1[39531] <= 16'b0000000000001111;
        weights1[39532] <= 16'b0000000000100010;
        weights1[39533] <= 16'b0000000000010001;
        weights1[39534] <= 16'b0000000000001001;
        weights1[39535] <= 16'b0000000000000111;
        weights1[39536] <= 16'b1111111111111010;
        weights1[39537] <= 16'b0000000000000011;
        weights1[39538] <= 16'b1111111111111100;
        weights1[39539] <= 16'b0000000000001000;
        weights1[39540] <= 16'b0000000000001000;
        weights1[39541] <= 16'b0000000000001010;
        weights1[39542] <= 16'b0000000000010001;
        weights1[39543] <= 16'b0000000000000100;
        weights1[39544] <= 16'b1111111111110111;
        weights1[39545] <= 16'b1111111111110110;
        weights1[39546] <= 16'b1111111111111010;
        weights1[39547] <= 16'b0000000000001110;
        weights1[39548] <= 16'b1111111111101001;
        weights1[39549] <= 16'b1111111111111110;
        weights1[39550] <= 16'b1111111111111000;
        weights1[39551] <= 16'b1111111111101101;
        weights1[39552] <= 16'b0000000000000000;
        weights1[39553] <= 16'b1111111111110110;
        weights1[39554] <= 16'b0000000000010010;
        weights1[39555] <= 16'b0000000000010010;
        weights1[39556] <= 16'b0000000000011011;
        weights1[39557] <= 16'b0000000000110000;
        weights1[39558] <= 16'b0000000000010111;
        weights1[39559] <= 16'b0000000000010100;
        weights1[39560] <= 16'b0000000000100001;
        weights1[39561] <= 16'b0000000000001101;
        weights1[39562] <= 16'b0000000000110101;
        weights1[39563] <= 16'b0000000000110110;
        weights1[39564] <= 16'b1111111111111111;
        weights1[39565] <= 16'b1111111111111100;
        weights1[39566] <= 16'b0000000000000111;
        weights1[39567] <= 16'b1111111111111100;
        weights1[39568] <= 16'b0000000000000011;
        weights1[39569] <= 16'b1111111111111010;
        weights1[39570] <= 16'b1111111111111111;
        weights1[39571] <= 16'b0000000000000010;
        weights1[39572] <= 16'b0000000000000100;
        weights1[39573] <= 16'b1111111111111110;
        weights1[39574] <= 16'b0000000000000101;
        weights1[39575] <= 16'b1111111111111101;
        weights1[39576] <= 16'b1111111111110111;
        weights1[39577] <= 16'b0000000000000011;
        weights1[39578] <= 16'b0000000000000000;
        weights1[39579] <= 16'b0000000000001010;
        weights1[39580] <= 16'b0000000000001001;
        weights1[39581] <= 16'b0000000000010110;
        weights1[39582] <= 16'b0000000000001101;
        weights1[39583] <= 16'b0000000000011100;
        weights1[39584] <= 16'b0000000000010111;
        weights1[39585] <= 16'b0000000000010001;
        weights1[39586] <= 16'b0000000000010111;
        weights1[39587] <= 16'b0000000000010101;
        weights1[39588] <= 16'b0000000000101110;
        weights1[39589] <= 16'b0000000000001000;
        weights1[39590] <= 16'b0000000000001100;
        weights1[39591] <= 16'b0000000000110010;
        weights1[39592] <= 16'b1111111111110111;
        weights1[39593] <= 16'b0000000000000100;
        weights1[39594] <= 16'b0000000000000111;
        weights1[39595] <= 16'b0000000000001000;
        weights1[39596] <= 16'b1111111111111110;
        weights1[39597] <= 16'b0000000000010011;
        weights1[39598] <= 16'b1111111111110000;
        weights1[39599] <= 16'b0000000000001101;
        weights1[39600] <= 16'b1111111111110011;
        weights1[39601] <= 16'b1111111111111101;
        weights1[39602] <= 16'b1111111111111111;
        weights1[39603] <= 16'b1111111111111100;
        weights1[39604] <= 16'b1111111111111011;
        weights1[39605] <= 16'b1111111111111011;
        weights1[39606] <= 16'b0000000000000110;
        weights1[39607] <= 16'b0000000000000010;
        weights1[39608] <= 16'b1111111111110111;
        weights1[39609] <= 16'b0000000000001000;
        weights1[39610] <= 16'b0000000000010011;
        weights1[39611] <= 16'b0000000000000001;
        weights1[39612] <= 16'b0000000000001111;
        weights1[39613] <= 16'b0000000000000000;
        weights1[39614] <= 16'b0000000000000010;
        weights1[39615] <= 16'b1111111111110101;
        weights1[39616] <= 16'b0000000000001111;
        weights1[39617] <= 16'b0000000000000010;
        weights1[39618] <= 16'b0000000000101001;
        weights1[39619] <= 16'b0000000000100001;
        weights1[39620] <= 16'b0000000000000000;
        weights1[39621] <= 16'b1111111111111010;
        weights1[39622] <= 16'b0000000000001011;
        weights1[39623] <= 16'b1111111111110111;
        weights1[39624] <= 16'b0000000000000100;
        weights1[39625] <= 16'b0000000000010001;
        weights1[39626] <= 16'b0000000000000110;
        weights1[39627] <= 16'b0000000000001010;
        weights1[39628] <= 16'b0000000000000010;
        weights1[39629] <= 16'b1111111111111110;
        weights1[39630] <= 16'b1111111111111001;
        weights1[39631] <= 16'b1111111111100111;
        weights1[39632] <= 16'b1111111111110000;
        weights1[39633] <= 16'b1111111111110111;
        weights1[39634] <= 16'b1111111111111111;
        weights1[39635] <= 16'b0000000000000000;
        weights1[39636] <= 16'b0000000000000101;
        weights1[39637] <= 16'b1111111111111001;
        weights1[39638] <= 16'b0000000000000001;
        weights1[39639] <= 16'b1111111111110001;
        weights1[39640] <= 16'b1111111111110111;
        weights1[39641] <= 16'b1111111111110111;
        weights1[39642] <= 16'b0000000000000101;
        weights1[39643] <= 16'b1111111111011010;
        weights1[39644] <= 16'b1111111111111001;
        weights1[39645] <= 16'b0000000000000011;
        weights1[39646] <= 16'b0000000000001110;
        weights1[39647] <= 16'b0000000000001100;
        weights1[39648] <= 16'b1111111111110001;
        weights1[39649] <= 16'b1111111111111101;
        weights1[39650] <= 16'b0000000000001010;
        weights1[39651] <= 16'b0000000000001001;
        weights1[39652] <= 16'b1111111111111110;
        weights1[39653] <= 16'b1111111111110101;
        weights1[39654] <= 16'b0000000000000100;
        weights1[39655] <= 16'b1111111111111110;
        weights1[39656] <= 16'b0000000000000011;
        weights1[39657] <= 16'b1111111111111110;
        weights1[39658] <= 16'b1111111111111110;
        weights1[39659] <= 16'b1111111111111011;
        weights1[39660] <= 16'b0000000000001011;
        weights1[39661] <= 16'b1111111111111101;
        weights1[39662] <= 16'b1111111111111100;
        weights1[39663] <= 16'b1111111111111001;
        weights1[39664] <= 16'b1111111111110000;
        weights1[39665] <= 16'b0000000000001110;
        weights1[39666] <= 16'b1111111111111101;
        weights1[39667] <= 16'b1111111111111001;
        weights1[39668] <= 16'b1111111111110001;
        weights1[39669] <= 16'b1111111111111010;
        weights1[39670] <= 16'b0000000000000000;
        weights1[39671] <= 16'b1111111111100101;
        weights1[39672] <= 16'b1111111111101111;
        weights1[39673] <= 16'b1111111111110001;
        weights1[39674] <= 16'b1111111111101001;
        weights1[39675] <= 16'b0000000000011010;
        weights1[39676] <= 16'b1111111111111010;
        weights1[39677] <= 16'b0000000000000001;
        weights1[39678] <= 16'b1111111111110111;
        weights1[39679] <= 16'b1111111111110101;
        weights1[39680] <= 16'b1111111111101111;
        weights1[39681] <= 16'b1111111111111101;
        weights1[39682] <= 16'b0000000000001010;
        weights1[39683] <= 16'b0000000000000101;
        weights1[39684] <= 16'b0000000000000001;
        weights1[39685] <= 16'b0000000000001010;
        weights1[39686] <= 16'b0000000000000001;
        weights1[39687] <= 16'b0000000000000010;
        weights1[39688] <= 16'b1111111111110110;
        weights1[39689] <= 16'b1111111111111000;
        weights1[39690] <= 16'b0000000000000110;
        weights1[39691] <= 16'b1111111111110101;
        weights1[39692] <= 16'b1111111111101110;
        weights1[39693] <= 16'b1111111111110011;
        weights1[39694] <= 16'b1111111111101111;
        weights1[39695] <= 16'b0000000000001100;
        weights1[39696] <= 16'b0000000000000010;
        weights1[39697] <= 16'b0000000000010001;
        weights1[39698] <= 16'b1111111111110011;
        weights1[39699] <= 16'b0000000000000010;
        weights1[39700] <= 16'b0000000000000101;
        weights1[39701] <= 16'b1111111111100111;
        weights1[39702] <= 16'b0000000000000001;
        weights1[39703] <= 16'b0000000000001000;
        weights1[39704] <= 16'b0000000000001000;
        weights1[39705] <= 16'b0000000000001010;
        weights1[39706] <= 16'b0000000000000110;
        weights1[39707] <= 16'b0000000000000011;
        weights1[39708] <= 16'b0000000000001011;
        weights1[39709] <= 16'b0000000000001010;
        weights1[39710] <= 16'b1111111111111010;
        weights1[39711] <= 16'b1111111111110110;
        weights1[39712] <= 16'b0000000000000100;
        weights1[39713] <= 16'b1111111111110110;
        weights1[39714] <= 16'b1111111111111010;
        weights1[39715] <= 16'b1111111111111111;
        weights1[39716] <= 16'b1111111111111000;
        weights1[39717] <= 16'b1111111111111100;
        weights1[39718] <= 16'b1111111111111000;
        weights1[39719] <= 16'b1111111111111100;
        weights1[39720] <= 16'b1111111111110111;
        weights1[39721] <= 16'b1111111111110100;
        weights1[39722] <= 16'b0000000000001101;
        weights1[39723] <= 16'b0000000000000011;
        weights1[39724] <= 16'b1111111111111010;
        weights1[39725] <= 16'b0000000000000101;
        weights1[39726] <= 16'b1111111111111100;
        weights1[39727] <= 16'b1111111111111111;
        weights1[39728] <= 16'b1111111111111101;
        weights1[39729] <= 16'b1111111111111001;
        weights1[39730] <= 16'b1111111111111111;
        weights1[39731] <= 16'b1111111111111111;
        weights1[39732] <= 16'b1111111111110110;
        weights1[39733] <= 16'b0000000000001101;
        weights1[39734] <= 16'b1111111111111100;
        weights1[39735] <= 16'b1111111111111111;
        weights1[39736] <= 16'b1111111111110011;
        weights1[39737] <= 16'b1111111111111101;
        weights1[39738] <= 16'b1111111111111110;
        weights1[39739] <= 16'b0000000000000010;
        weights1[39740] <= 16'b1111111111111000;
        weights1[39741] <= 16'b1111111111111111;
        weights1[39742] <= 16'b0000000000000000;
        weights1[39743] <= 16'b0000000000000101;
        weights1[39744] <= 16'b0000000000001101;
        weights1[39745] <= 16'b0000000000000010;
        weights1[39746] <= 16'b0000000000000100;
        weights1[39747] <= 16'b0000000000000011;
        weights1[39748] <= 16'b1111111111111001;
        weights1[39749] <= 16'b0000000000000111;
        weights1[39750] <= 16'b1111111111101111;
        weights1[39751] <= 16'b1111111111110100;
        weights1[39752] <= 16'b0000000000000011;
        weights1[39753] <= 16'b1111111111101011;
        weights1[39754] <= 16'b0000000000000000;
        weights1[39755] <= 16'b1111111111110010;
        weights1[39756] <= 16'b0000000000001111;
        weights1[39757] <= 16'b1111111111111100;
        weights1[39758] <= 16'b1111111111111110;
        weights1[39759] <= 16'b0000000000000101;
        weights1[39760] <= 16'b1111111111110101;
        weights1[39761] <= 16'b1111111111101100;
        weights1[39762] <= 16'b0000000000000100;
        weights1[39763] <= 16'b0000000000000011;
        weights1[39764] <= 16'b1111111111110101;
        weights1[39765] <= 16'b1111111111111110;
        weights1[39766] <= 16'b1111111111111011;
        weights1[39767] <= 16'b0000000000000001;
        weights1[39768] <= 16'b0000000000001000;
        weights1[39769] <= 16'b0000000000010011;
        weights1[39770] <= 16'b1111111111101101;
        weights1[39771] <= 16'b0000000000000011;
        weights1[39772] <= 16'b0000000000001100;
        weights1[39773] <= 16'b1111111111110110;
        weights1[39774] <= 16'b0000000000000110;
        weights1[39775] <= 16'b0000000000000101;
        weights1[39776] <= 16'b0000000000000110;
        weights1[39777] <= 16'b1111111111111111;
        weights1[39778] <= 16'b1111111111111111;
        weights1[39779] <= 16'b0000000000001010;
        weights1[39780] <= 16'b1111111111110110;
        weights1[39781] <= 16'b1111111111111110;
        weights1[39782] <= 16'b0000000000011100;
        weights1[39783] <= 16'b0000000000011100;
        weights1[39784] <= 16'b1111111111110001;
        weights1[39785] <= 16'b0000000000000010;
        weights1[39786] <= 16'b1111111111110111;
        weights1[39787] <= 16'b1111111111110110;
        weights1[39788] <= 16'b1111111111111010;
        weights1[39789] <= 16'b1111111111111111;
        weights1[39790] <= 16'b0000000000000110;
        weights1[39791] <= 16'b0000000000001000;
        weights1[39792] <= 16'b1111111111111011;
        weights1[39793] <= 16'b0000000000000111;
        weights1[39794] <= 16'b0000000000010000;
        weights1[39795] <= 16'b1111111111101010;
        weights1[39796] <= 16'b1111111111111010;
        weights1[39797] <= 16'b0000000000000000;
        weights1[39798] <= 16'b1111111111111001;
        weights1[39799] <= 16'b0000000000000001;
        weights1[39800] <= 16'b0000000000000000;
        weights1[39801] <= 16'b0000000000000111;
        weights1[39802] <= 16'b0000000000000001;
        weights1[39803] <= 16'b1111111111111100;
        weights1[39804] <= 16'b1111111111111001;
        weights1[39805] <= 16'b0000000000000010;
        weights1[39806] <= 16'b1111111111111100;
        weights1[39807] <= 16'b1111111111111100;
        weights1[39808] <= 16'b0000000000010111;
        weights1[39809] <= 16'b1111111111111000;
        weights1[39810] <= 16'b1111111111110001;
        weights1[39811] <= 16'b1111111111110101;
        weights1[39812] <= 16'b1111111111101110;
        weights1[39813] <= 16'b0000000000001010;
        weights1[39814] <= 16'b1111111111100001;
        weights1[39815] <= 16'b1111111111110011;
        weights1[39816] <= 16'b1111111111111000;
        weights1[39817] <= 16'b0000000000000101;
        weights1[39818] <= 16'b0000000000000001;
        weights1[39819] <= 16'b1111111111111001;
        weights1[39820] <= 16'b1111111111111111;
        weights1[39821] <= 16'b1111111111111010;
        weights1[39822] <= 16'b1111111111111010;
        weights1[39823] <= 16'b1111111111110111;
        weights1[39824] <= 16'b0000000000001100;
        weights1[39825] <= 16'b1111111111111010;
        weights1[39826] <= 16'b1111111111111101;
        weights1[39827] <= 16'b1111111111111010;
        weights1[39828] <= 16'b1111111111110110;
        weights1[39829] <= 16'b1111111111110100;
        weights1[39830] <= 16'b1111111111111001;
        weights1[39831] <= 16'b0000000000000100;
        weights1[39832] <= 16'b0000000000000100;
        weights1[39833] <= 16'b0000000000000101;
        weights1[39834] <= 16'b1111111111111011;
        weights1[39835] <= 16'b0000000000010001;
        weights1[39836] <= 16'b1111111111110101;
        weights1[39837] <= 16'b1111111111111101;
        weights1[39838] <= 16'b1111111111111100;
        weights1[39839] <= 16'b1111111111111111;
        weights1[39840] <= 16'b1111111111111111;
        weights1[39841] <= 16'b0000000000000101;
        weights1[39842] <= 16'b1111111111110010;
        weights1[39843] <= 16'b0000000000000100;
        weights1[39844] <= 16'b0000000000000011;
        weights1[39845] <= 16'b1111111111111110;
        weights1[39846] <= 16'b1111111111111111;
        weights1[39847] <= 16'b0000000000001101;
        weights1[39848] <= 16'b0000000000000011;
        weights1[39849] <= 16'b0000000000000000;
        weights1[39850] <= 16'b0000000000000001;
        weights1[39851] <= 16'b1111111111111101;
        weights1[39852] <= 16'b1111111111110011;
        weights1[39853] <= 16'b0000000000000110;
        weights1[39854] <= 16'b0000000000000001;
        weights1[39855] <= 16'b0000000000011101;
        weights1[39856] <= 16'b0000000000001100;
        weights1[39857] <= 16'b1111111111111001;
        weights1[39858] <= 16'b1111111111111101;
        weights1[39859] <= 16'b0000000000000001;
        weights1[39860] <= 16'b1111111111101100;
        weights1[39861] <= 16'b1111111111110000;
        weights1[39862] <= 16'b1111111111101011;
        weights1[39863] <= 16'b0000000000000011;
        weights1[39864] <= 16'b0000000000001001;
        weights1[39865] <= 16'b1111111111110001;
        weights1[39866] <= 16'b1111111111101101;
        weights1[39867] <= 16'b0000000000000010;
        weights1[39868] <= 16'b1111111111101000;
        weights1[39869] <= 16'b1111111111111011;
        weights1[39870] <= 16'b1111111111110100;
        weights1[39871] <= 16'b1111111111110111;
        weights1[39872] <= 16'b1111111111111111;
        weights1[39873] <= 16'b0000000000000111;
        weights1[39874] <= 16'b0000000000001010;
        weights1[39875] <= 16'b0000000000001001;
        weights1[39876] <= 16'b1111111111110111;
        weights1[39877] <= 16'b0000000000000010;
        weights1[39878] <= 16'b1111111111110011;
        weights1[39879] <= 16'b1111111111110111;
        weights1[39880] <= 16'b0000000000001000;
        weights1[39881] <= 16'b1111111111101100;
        weights1[39882] <= 16'b1111111111111011;
        weights1[39883] <= 16'b1111111111110110;
        weights1[39884] <= 16'b0000000000001010;
        weights1[39885] <= 16'b1111111111110110;
        weights1[39886] <= 16'b1111111111111101;
        weights1[39887] <= 16'b0000000000000100;
        weights1[39888] <= 16'b0000000000000110;
        weights1[39889] <= 16'b0000000000001001;
        weights1[39890] <= 16'b1111111111101000;
        weights1[39891] <= 16'b0000000000010011;
        weights1[39892] <= 16'b1111111111110010;
        weights1[39893] <= 16'b1111111111110101;
        weights1[39894] <= 16'b1111111111110000;
        weights1[39895] <= 16'b1111111111110111;
        weights1[39896] <= 16'b1111111111100101;
        weights1[39897] <= 16'b1111111111101100;
        weights1[39898] <= 16'b1111111111110011;
        weights1[39899] <= 16'b1111111111111011;
        weights1[39900] <= 16'b1111111111111011;
        weights1[39901] <= 16'b0000000000000011;
        weights1[39902] <= 16'b1111111111110101;
        weights1[39903] <= 16'b0000000000001011;
        weights1[39904] <= 16'b1111111111111001;
        weights1[39905] <= 16'b0000000000010101;
        weights1[39906] <= 16'b1111111111111000;
        weights1[39907] <= 16'b1111111111111111;
        weights1[39908] <= 16'b1111111111111011;
        weights1[39909] <= 16'b1111111111101101;
        weights1[39910] <= 16'b1111111111111000;
        weights1[39911] <= 16'b1111111111110011;
        weights1[39912] <= 16'b1111111111101100;
        weights1[39913] <= 16'b1111111111110011;
        weights1[39914] <= 16'b1111111111110000;
        weights1[39915] <= 16'b0000000000000000;
        weights1[39916] <= 16'b0000000000000000;
        weights1[39917] <= 16'b0000000000000001;
        weights1[39918] <= 16'b0000000000000111;
        weights1[39919] <= 16'b1111111111111110;
        weights1[39920] <= 16'b0000000000000010;
        weights1[39921] <= 16'b1111111111110000;
        weights1[39922] <= 16'b1111111111101100;
        weights1[39923] <= 16'b1111111111110110;
        weights1[39924] <= 16'b1111111111101110;
        weights1[39925] <= 16'b1111111111110101;
        weights1[39926] <= 16'b1111111111110101;
        weights1[39927] <= 16'b1111111111111100;
        weights1[39928] <= 16'b1111111111111101;
        weights1[39929] <= 16'b1111111111111101;
        weights1[39930] <= 16'b1111111111111110;
        weights1[39931] <= 16'b1111111111111111;
        weights1[39932] <= 16'b1111111111111101;
        weights1[39933] <= 16'b0000000000000100;
        weights1[39934] <= 16'b1111111111111111;
        weights1[39935] <= 16'b1111111111111010;
        weights1[39936] <= 16'b0000000000001110;
        weights1[39937] <= 16'b0000000000000111;
        weights1[39938] <= 16'b0000000000000101;
        weights1[39939] <= 16'b1111111111111101;
        weights1[39940] <= 16'b0000000000000111;
        weights1[39941] <= 16'b0000000000001111;
        weights1[39942] <= 16'b1111111111101111;
        weights1[39943] <= 16'b1111111111111100;
        weights1[39944] <= 16'b1111111111101111;
        weights1[39945] <= 16'b1111111111101100;
        weights1[39946] <= 16'b1111111111111001;
        weights1[39947] <= 16'b1111111111101001;
        weights1[39948] <= 16'b1111111111110100;
        weights1[39949] <= 16'b1111111111101001;
        weights1[39950] <= 16'b1111111111101010;
        weights1[39951] <= 16'b1111111111110100;
        weights1[39952] <= 16'b1111111111111011;
        weights1[39953] <= 16'b1111111111111111;
        weights1[39954] <= 16'b1111111111111110;
        weights1[39955] <= 16'b0000000000000001;
        weights1[39956] <= 16'b1111111111111110;
        weights1[39957] <= 16'b1111111111111101;
        weights1[39958] <= 16'b0000000000000111;
        weights1[39959] <= 16'b0000000000001001;
        weights1[39960] <= 16'b0000000000000001;
        weights1[39961] <= 16'b0000000000001011;
        weights1[39962] <= 16'b1111111111111110;
        weights1[39963] <= 16'b0000000000000001;
        weights1[39964] <= 16'b0000000000000011;
        weights1[39965] <= 16'b0000000000000001;
        weights1[39966] <= 16'b1111111111101010;
        weights1[39967] <= 16'b1111111111011101;
        weights1[39968] <= 16'b1111111111100000;
        weights1[39969] <= 16'b1111111111011101;
        weights1[39970] <= 16'b1111111111011010;
        weights1[39971] <= 16'b1111111111011101;
        weights1[39972] <= 16'b1111111111100010;
        weights1[39973] <= 16'b1111111111011110;
        weights1[39974] <= 16'b1111111111011111;
        weights1[39975] <= 16'b1111111111100010;
        weights1[39976] <= 16'b1111111111101110;
        weights1[39977] <= 16'b1111111111101011;
        weights1[39978] <= 16'b1111111111110111;
        weights1[39979] <= 16'b1111111111111010;
        weights1[39980] <= 16'b0000000000000000;
        weights1[39981] <= 16'b0000000000000001;
        weights1[39982] <= 16'b0000000000000001;
        weights1[39983] <= 16'b0000000000000100;
        weights1[39984] <= 16'b0000000000000000;
        weights1[39985] <= 16'b0000000000000001;
        weights1[39986] <= 16'b0000000000000001;
        weights1[39987] <= 16'b1111111111111110;
        weights1[39988] <= 16'b0000000000000001;
        weights1[39989] <= 16'b1111111111110111;
        weights1[39990] <= 16'b1111111111110111;
        weights1[39991] <= 16'b1111111111110100;
        weights1[39992] <= 16'b1111111111101110;
        weights1[39993] <= 16'b1111111111110100;
        weights1[39994] <= 16'b1111111111110010;
        weights1[39995] <= 16'b1111111111111000;
        weights1[39996] <= 16'b1111111111111011;
        weights1[39997] <= 16'b1111111111111011;
        weights1[39998] <= 16'b1111111111110111;
        weights1[39999] <= 16'b1111111111110001;
        weights1[40000] <= 16'b1111111111111011;
        weights1[40001] <= 16'b1111111111110100;
        weights1[40002] <= 16'b1111111111111011;
        weights1[40003] <= 16'b1111111111111000;
        weights1[40004] <= 16'b1111111111111001;
        weights1[40005] <= 16'b1111111111111110;
        weights1[40006] <= 16'b1111111111111010;
        weights1[40007] <= 16'b0000000000000000;
        weights1[40008] <= 16'b0000000000000100;
        weights1[40009] <= 16'b0000000000000100;
        weights1[40010] <= 16'b0000000000000011;
        weights1[40011] <= 16'b0000000000000010;
        weights1[40012] <= 16'b0000000000000000;
        weights1[40013] <= 16'b0000000000000001;
        weights1[40014] <= 16'b1111111111111100;
        weights1[40015] <= 16'b1111111111111101;
        weights1[40016] <= 16'b1111111111110101;
        weights1[40017] <= 16'b1111111111111010;
        weights1[40018] <= 16'b1111111111110101;
        weights1[40019] <= 16'b1111111111110100;
        weights1[40020] <= 16'b1111111111110001;
        weights1[40021] <= 16'b1111111111101110;
        weights1[40022] <= 16'b1111111111111001;
        weights1[40023] <= 16'b1111111111111100;
        weights1[40024] <= 16'b1111111111111101;
        weights1[40025] <= 16'b1111111111111010;
        weights1[40026] <= 16'b1111111111110111;
        weights1[40027] <= 16'b1111111111101110;
        weights1[40028] <= 16'b1111111111110011;
        weights1[40029] <= 16'b1111111111111011;
        weights1[40030] <= 16'b1111111111111010;
        weights1[40031] <= 16'b1111111111110110;
        weights1[40032] <= 16'b1111111111110100;
        weights1[40033] <= 16'b1111111111101111;
        weights1[40034] <= 16'b1111111111110010;
        weights1[40035] <= 16'b1111111111111001;
        weights1[40036] <= 16'b1111111111111111;
        weights1[40037] <= 16'b1111111111111111;
        weights1[40038] <= 16'b0000000000000011;
        weights1[40039] <= 16'b0000000000000010;
        weights1[40040] <= 16'b0000000000000000;
        weights1[40041] <= 16'b1111111111111101;
        weights1[40042] <= 16'b1111111111111001;
        weights1[40043] <= 16'b1111111111111001;
        weights1[40044] <= 16'b0000000000000001;
        weights1[40045] <= 16'b1111111111111101;
        weights1[40046] <= 16'b1111111111110110;
        weights1[40047] <= 16'b1111111111111000;
        weights1[40048] <= 16'b1111111111111110;
        weights1[40049] <= 16'b0000000000000011;
        weights1[40050] <= 16'b1111111111110111;
        weights1[40051] <= 16'b1111111111110111;
        weights1[40052] <= 16'b1111111111111101;
        weights1[40053] <= 16'b1111111111110100;
        weights1[40054] <= 16'b1111111111101110;
        weights1[40055] <= 16'b1111111111101100;
        weights1[40056] <= 16'b1111111111101001;
        weights1[40057] <= 16'b1111111111110000;
        weights1[40058] <= 16'b1111111111110100;
        weights1[40059] <= 16'b1111111111110100;
        weights1[40060] <= 16'b1111111111101110;
        weights1[40061] <= 16'b1111111111101101;
        weights1[40062] <= 16'b1111111111110000;
        weights1[40063] <= 16'b1111111111110111;
        weights1[40064] <= 16'b1111111111110100;
        weights1[40065] <= 16'b1111111111111001;
        weights1[40066] <= 16'b1111111111111111;
        weights1[40067] <= 16'b0000000000000010;
        weights1[40068] <= 16'b1111111111111101;
        weights1[40069] <= 16'b1111111111110110;
        weights1[40070] <= 16'b1111111111110011;
        weights1[40071] <= 16'b1111111111110111;
        weights1[40072] <= 16'b1111111111111110;
        weights1[40073] <= 16'b0000000000000010;
        weights1[40074] <= 16'b0000000000000000;
        weights1[40075] <= 16'b1111111111111010;
        weights1[40076] <= 16'b0000000000000100;
        weights1[40077] <= 16'b0000000000000100;
        weights1[40078] <= 16'b1111111111110110;
        weights1[40079] <= 16'b1111111111111010;
        weights1[40080] <= 16'b0000000000000001;
        weights1[40081] <= 16'b0000000000000111;
        weights1[40082] <= 16'b0000000000000000;
        weights1[40083] <= 16'b1111111111110011;
        weights1[40084] <= 16'b1111111111110001;
        weights1[40085] <= 16'b1111111111100011;
        weights1[40086] <= 16'b1111111111101101;
        weights1[40087] <= 16'b1111111111111001;
        weights1[40088] <= 16'b0000000000000010;
        weights1[40089] <= 16'b1111111111110000;
        weights1[40090] <= 16'b1111111111111011;
        weights1[40091] <= 16'b1111111111111001;
        weights1[40092] <= 16'b1111111111110101;
        weights1[40093] <= 16'b1111111111111011;
        weights1[40094] <= 16'b0000000000000100;
        weights1[40095] <= 16'b1111111111111111;
        weights1[40096] <= 16'b1111111111111010;
        weights1[40097] <= 16'b1111111111110011;
        weights1[40098] <= 16'b1111111111110000;
        weights1[40099] <= 16'b1111111111110000;
        weights1[40100] <= 16'b0000000000000000;
        weights1[40101] <= 16'b0000000000000111;
        weights1[40102] <= 16'b0000000000000100;
        weights1[40103] <= 16'b0000000000000110;
        weights1[40104] <= 16'b0000000000001101;
        weights1[40105] <= 16'b0000000000000110;
        weights1[40106] <= 16'b1111111111111010;
        weights1[40107] <= 16'b1111111111110100;
        weights1[40108] <= 16'b1111111111111001;
        weights1[40109] <= 16'b1111111111111000;
        weights1[40110] <= 16'b1111111111110101;
        weights1[40111] <= 16'b1111111111101111;
        weights1[40112] <= 16'b0000000000000001;
        weights1[40113] <= 16'b1111111111111011;
        weights1[40114] <= 16'b1111111111111011;
        weights1[40115] <= 16'b1111111111111111;
        weights1[40116] <= 16'b0000000000000000;
        weights1[40117] <= 16'b1111111111111101;
        weights1[40118] <= 16'b0000000000000011;
        weights1[40119] <= 16'b0000000000000101;
        weights1[40120] <= 16'b1111111111111110;
        weights1[40121] <= 16'b1111111111111100;
        weights1[40122] <= 16'b1111111111111110;
        weights1[40123] <= 16'b0000000000000001;
        weights1[40124] <= 16'b1111111111111001;
        weights1[40125] <= 16'b1111111111110100;
        weights1[40126] <= 16'b1111111111101111;
        weights1[40127] <= 16'b1111111111110010;
        weights1[40128] <= 16'b1111111111111101;
        weights1[40129] <= 16'b1111111111111110;
        weights1[40130] <= 16'b0000000000010010;
        weights1[40131] <= 16'b0000000000010011;
        weights1[40132] <= 16'b0000000000010100;
        weights1[40133] <= 16'b1111111111111110;
        weights1[40134] <= 16'b1111111111110101;
        weights1[40135] <= 16'b1111111111110111;
        weights1[40136] <= 16'b1111111111110111;
        weights1[40137] <= 16'b1111111111111011;
        weights1[40138] <= 16'b0000000000000000;
        weights1[40139] <= 16'b0000000000001001;
        weights1[40140] <= 16'b0000000000000000;
        weights1[40141] <= 16'b0000000000000101;
        weights1[40142] <= 16'b0000000000001000;
        weights1[40143] <= 16'b0000000000001011;
        weights1[40144] <= 16'b0000000000001001;
        weights1[40145] <= 16'b1111111111111110;
        weights1[40146] <= 16'b1111111111111010;
        weights1[40147] <= 16'b0000000000000000;
        weights1[40148] <= 16'b0000000000001000;
        weights1[40149] <= 16'b0000000000000001;
        weights1[40150] <= 16'b0000000000000111;
        weights1[40151] <= 16'b0000000000000010;
        weights1[40152] <= 16'b1111111111111001;
        weights1[40153] <= 16'b1111111111111010;
        weights1[40154] <= 16'b1111111111110111;
        weights1[40155] <= 16'b1111111111110111;
        weights1[40156] <= 16'b1111111111111100;
        weights1[40157] <= 16'b0000000000010001;
        weights1[40158] <= 16'b0000000000011010;
        weights1[40159] <= 16'b0000000000011010;
        weights1[40160] <= 16'b0000000000010011;
        weights1[40161] <= 16'b0000000000000100;
        weights1[40162] <= 16'b1111111111110101;
        weights1[40163] <= 16'b0000000000000000;
        weights1[40164] <= 16'b0000000000000011;
        weights1[40165] <= 16'b0000000000000010;
        weights1[40166] <= 16'b1111111111110111;
        weights1[40167] <= 16'b1111111111111110;
        weights1[40168] <= 16'b0000000000000111;
        weights1[40169] <= 16'b0000000000000111;
        weights1[40170] <= 16'b0000000000010000;
        weights1[40171] <= 16'b0000000000010010;
        weights1[40172] <= 16'b0000000000010110;
        weights1[40173] <= 16'b0000000000010110;
        weights1[40174] <= 16'b0000000000011000;
        weights1[40175] <= 16'b0000000000001100;
        weights1[40176] <= 16'b0000000000001001;
        weights1[40177] <= 16'b0000000000001011;
        weights1[40178] <= 16'b0000000000001100;
        weights1[40179] <= 16'b0000000000000001;
        weights1[40180] <= 16'b1111111111111100;
        weights1[40181] <= 16'b1111111111111101;
        weights1[40182] <= 16'b1111111111111000;
        weights1[40183] <= 16'b1111111111111111;
        weights1[40184] <= 16'b0000000000001010;
        weights1[40185] <= 16'b0000000000001100;
        weights1[40186] <= 16'b0000000000011110;
        weights1[40187] <= 16'b0000000000100111;
        weights1[40188] <= 16'b0000000000010010;
        weights1[40189] <= 16'b0000000000001110;
        weights1[40190] <= 16'b0000000000001011;
        weights1[40191] <= 16'b0000000000001010;
        weights1[40192] <= 16'b0000000000000110;
        weights1[40193] <= 16'b0000000000001001;
        weights1[40194] <= 16'b0000000000000110;
        weights1[40195] <= 16'b0000000000001001;
        weights1[40196] <= 16'b0000000000001100;
        weights1[40197] <= 16'b0000000000001001;
        weights1[40198] <= 16'b0000000000001111;
        weights1[40199] <= 16'b0000000000011001;
        weights1[40200] <= 16'b0000000000010111;
        weights1[40201] <= 16'b0000000000010100;
        weights1[40202] <= 16'b0000000000011000;
        weights1[40203] <= 16'b0000000000011010;
        weights1[40204] <= 16'b0000000000010011;
        weights1[40205] <= 16'b0000000000010010;
        weights1[40206] <= 16'b0000000000001111;
        weights1[40207] <= 16'b0000000000001100;
        weights1[40208] <= 16'b1111111111111000;
        weights1[40209] <= 16'b1111111111111001;
        weights1[40210] <= 16'b1111111111111100;
        weights1[40211] <= 16'b0000000000000101;
        weights1[40212] <= 16'b0000000000000011;
        weights1[40213] <= 16'b0000000000010100;
        weights1[40214] <= 16'b0000000000011100;
        weights1[40215] <= 16'b0000000000011000;
        weights1[40216] <= 16'b0000000000011001;
        weights1[40217] <= 16'b0000000000100010;
        weights1[40218] <= 16'b0000000000001011;
        weights1[40219] <= 16'b1111111111110110;
        weights1[40220] <= 16'b0000000000000001;
        weights1[40221] <= 16'b0000000000011000;
        weights1[40222] <= 16'b0000000000010001;
        weights1[40223] <= 16'b0000000000001100;
        weights1[40224] <= 16'b0000000000001100;
        weights1[40225] <= 16'b0000000000001010;
        weights1[40226] <= 16'b0000000000011000;
        weights1[40227] <= 16'b0000000000010100;
        weights1[40228] <= 16'b0000000000010011;
        weights1[40229] <= 16'b0000000000010010;
        weights1[40230] <= 16'b0000000000011001;
        weights1[40231] <= 16'b0000000000010101;
        weights1[40232] <= 16'b0000000000011110;
        weights1[40233] <= 16'b0000000000010001;
        weights1[40234] <= 16'b0000000000001111;
        weights1[40235] <= 16'b0000000000011001;
        weights1[40236] <= 16'b1111111111111001;
        weights1[40237] <= 16'b1111111111111010;
        weights1[40238] <= 16'b0000000000000010;
        weights1[40239] <= 16'b0000000000010001;
        weights1[40240] <= 16'b0000000000000100;
        weights1[40241] <= 16'b0000000000010111;
        weights1[40242] <= 16'b0000000000100110;
        weights1[40243] <= 16'b0000000000100110;
        weights1[40244] <= 16'b0000000000010100;
        weights1[40245] <= 16'b0000000000001100;
        weights1[40246] <= 16'b0000000000000010;
        weights1[40247] <= 16'b0000000000000001;
        weights1[40248] <= 16'b0000000000001001;
        weights1[40249] <= 16'b0000000000001101;
        weights1[40250] <= 16'b0000000000001111;
        weights1[40251] <= 16'b0000000000001001;
        weights1[40252] <= 16'b0000000000000101;
        weights1[40253] <= 16'b0000000000001011;
        weights1[40254] <= 16'b0000000000010001;
        weights1[40255] <= 16'b0000000000011001;
        weights1[40256] <= 16'b0000000000011000;
        weights1[40257] <= 16'b0000000000011001;
        weights1[40258] <= 16'b0000000000011011;
        weights1[40259] <= 16'b0000000000010110;
        weights1[40260] <= 16'b0000000000011001;
        weights1[40261] <= 16'b0000000000001010;
        weights1[40262] <= 16'b0000000000001100;
        weights1[40263] <= 16'b0000000000010110;
        weights1[40264] <= 16'b1111111111111110;
        weights1[40265] <= 16'b0000000000000101;
        weights1[40266] <= 16'b0000000000001101;
        weights1[40267] <= 16'b0000000000000101;
        weights1[40268] <= 16'b0000000000000110;
        weights1[40269] <= 16'b0000000000011101;
        weights1[40270] <= 16'b0000000000100100;
        weights1[40271] <= 16'b0000000000011011;
        weights1[40272] <= 16'b0000000000010110;
        weights1[40273] <= 16'b0000000000000100;
        weights1[40274] <= 16'b1111111111110110;
        weights1[40275] <= 16'b0000000000000101;
        weights1[40276] <= 16'b0000000000001011;
        weights1[40277] <= 16'b0000000000010111;
        weights1[40278] <= 16'b0000000000010010;
        weights1[40279] <= 16'b1111111111111111;
        weights1[40280] <= 16'b0000000000000001;
        weights1[40281] <= 16'b0000000000001011;
        weights1[40282] <= 16'b0000000000000111;
        weights1[40283] <= 16'b0000000000011000;
        weights1[40284] <= 16'b0000000000011011;
        weights1[40285] <= 16'b0000000000011001;
        weights1[40286] <= 16'b0000000000010100;
        weights1[40287] <= 16'b0000000000010001;
        weights1[40288] <= 16'b0000000000010111;
        weights1[40289] <= 16'b0000000000000100;
        weights1[40290] <= 16'b0000000000010100;
        weights1[40291] <= 16'b0000000000001111;
        weights1[40292] <= 16'b1111111111111111;
        weights1[40293] <= 16'b0000000000000001;
        weights1[40294] <= 16'b0000000000000010;
        weights1[40295] <= 16'b0000000000000101;
        weights1[40296] <= 16'b0000000000001011;
        weights1[40297] <= 16'b0000000000001011;
        weights1[40298] <= 16'b0000000000010011;
        weights1[40299] <= 16'b0000000000100101;
        weights1[40300] <= 16'b0000000000011010;
        weights1[40301] <= 16'b0000000000000101;
        weights1[40302] <= 16'b1111111111111110;
        weights1[40303] <= 16'b0000000000000000;
        weights1[40304] <= 16'b0000000000000111;
        weights1[40305] <= 16'b0000000000000011;
        weights1[40306] <= 16'b1111111111111100;
        weights1[40307] <= 16'b1111111111111010;
        weights1[40308] <= 16'b1111111111111001;
        weights1[40309] <= 16'b1111111111111011;
        weights1[40310] <= 16'b1111111111110000;
        weights1[40311] <= 16'b1111111111111101;
        weights1[40312] <= 16'b0000000000001010;
        weights1[40313] <= 16'b0000000000011001;
        weights1[40314] <= 16'b0000000000011010;
        weights1[40315] <= 16'b0000000000011011;
        weights1[40316] <= 16'b0000000000001101;
        weights1[40317] <= 16'b0000000000000100;
        weights1[40318] <= 16'b0000000000001010;
        weights1[40319] <= 16'b0000000000001101;
        weights1[40320] <= 16'b1111111111111110;
        weights1[40321] <= 16'b0000000000000110;
        weights1[40322] <= 16'b0000000000001011;
        weights1[40323] <= 16'b0000000000001111;
        weights1[40324] <= 16'b0000000000001011;
        weights1[40325] <= 16'b0000000000001011;
        weights1[40326] <= 16'b0000000000011111;
        weights1[40327] <= 16'b0000000000011010;
        weights1[40328] <= 16'b0000000000001111;
        weights1[40329] <= 16'b1111111111110101;
        weights1[40330] <= 16'b1111111111110011;
        weights1[40331] <= 16'b0000000000000000;
        weights1[40332] <= 16'b0000000000000010;
        weights1[40333] <= 16'b0000000000001101;
        weights1[40334] <= 16'b1111111111111100;
        weights1[40335] <= 16'b1111111111110000;
        weights1[40336] <= 16'b1111111111100111;
        weights1[40337] <= 16'b1111111111101010;
        weights1[40338] <= 16'b1111111111101110;
        weights1[40339] <= 16'b1111111111110010;
        weights1[40340] <= 16'b0000000000001100;
        weights1[40341] <= 16'b0000000000010001;
        weights1[40342] <= 16'b0000000000100000;
        weights1[40343] <= 16'b0000000000100101;
        weights1[40344] <= 16'b0000000000011111;
        weights1[40345] <= 16'b0000000000001101;
        weights1[40346] <= 16'b0000000000001100;
        weights1[40347] <= 16'b0000000000001010;
        weights1[40348] <= 16'b0000000000000010;
        weights1[40349] <= 16'b0000000000000011;
        weights1[40350] <= 16'b0000000000000110;
        weights1[40351] <= 16'b0000000000010100;
        weights1[40352] <= 16'b0000000000011001;
        weights1[40353] <= 16'b0000000000010111;
        weights1[40354] <= 16'b0000000000100100;
        weights1[40355] <= 16'b0000000000010011;
        weights1[40356] <= 16'b0000000000001110;
        weights1[40357] <= 16'b0000000000000001;
        weights1[40358] <= 16'b1111111111110000;
        weights1[40359] <= 16'b1111111111110110;
        weights1[40360] <= 16'b0000000000000000;
        weights1[40361] <= 16'b0000000000000001;
        weights1[40362] <= 16'b1111111111101010;
        weights1[40363] <= 16'b1111111111101010;
        weights1[40364] <= 16'b1111111111101000;
        weights1[40365] <= 16'b1111111111011111;
        weights1[40366] <= 16'b1111111111011101;
        weights1[40367] <= 16'b1111111111101111;
        weights1[40368] <= 16'b1111111111111101;
        weights1[40369] <= 16'b0000000000010100;
        weights1[40370] <= 16'b0000000000010101;
        weights1[40371] <= 16'b0000000000100000;
        weights1[40372] <= 16'b0000000000011011;
        weights1[40373] <= 16'b0000000000011010;
        weights1[40374] <= 16'b0000000000001010;
        weights1[40375] <= 16'b0000000000001101;
        weights1[40376] <= 16'b1111111111111111;
        weights1[40377] <= 16'b0000000000000011;
        weights1[40378] <= 16'b1111111111111011;
        weights1[40379] <= 16'b0000000000001100;
        weights1[40380] <= 16'b0000000000010011;
        weights1[40381] <= 16'b0000000000011101;
        weights1[40382] <= 16'b0000000000011010;
        weights1[40383] <= 16'b0000000000010100;
        weights1[40384] <= 16'b0000000000000100;
        weights1[40385] <= 16'b0000000000000010;
        weights1[40386] <= 16'b1111111111110000;
        weights1[40387] <= 16'b1111111111100101;
        weights1[40388] <= 16'b1111111111110000;
        weights1[40389] <= 16'b1111111111101101;
        weights1[40390] <= 16'b1111111111101111;
        weights1[40391] <= 16'b1111111111101100;
        weights1[40392] <= 16'b1111111111101011;
        weights1[40393] <= 16'b1111111111101111;
        weights1[40394] <= 16'b1111111111101100;
        weights1[40395] <= 16'b1111111111101010;
        weights1[40396] <= 16'b1111111111101011;
        weights1[40397] <= 16'b0000000000000100;
        weights1[40398] <= 16'b0000000000100011;
        weights1[40399] <= 16'b0000000000100010;
        weights1[40400] <= 16'b0000000000100001;
        weights1[40401] <= 16'b0000000000010011;
        weights1[40402] <= 16'b0000000000010110;
        weights1[40403] <= 16'b0000000000010001;
        weights1[40404] <= 16'b1111111111111001;
        weights1[40405] <= 16'b1111111111111001;
        weights1[40406] <= 16'b0000000000000110;
        weights1[40407] <= 16'b0000000000000100;
        weights1[40408] <= 16'b0000000000001010;
        weights1[40409] <= 16'b0000000000011100;
        weights1[40410] <= 16'b0000000000011111;
        weights1[40411] <= 16'b0000000000011000;
        weights1[40412] <= 16'b0000000000000111;
        weights1[40413] <= 16'b1111111111101110;
        weights1[40414] <= 16'b1111111111101111;
        weights1[40415] <= 16'b1111111111101001;
        weights1[40416] <= 16'b1111111111101101;
        weights1[40417] <= 16'b1111111111110010;
        weights1[40418] <= 16'b1111111111110011;
        weights1[40419] <= 16'b1111111111110001;
        weights1[40420] <= 16'b1111111111110011;
        weights1[40421] <= 16'b1111111111100001;
        weights1[40422] <= 16'b1111111111101001;
        weights1[40423] <= 16'b1111111111100111;
        weights1[40424] <= 16'b1111111111100101;
        weights1[40425] <= 16'b0000000000000000;
        weights1[40426] <= 16'b0000000000001110;
        weights1[40427] <= 16'b0000000000011001;
        weights1[40428] <= 16'b0000000000011010;
        weights1[40429] <= 16'b0000000000011001;
        weights1[40430] <= 16'b0000000000001110;
        weights1[40431] <= 16'b0000000000001101;
        weights1[40432] <= 16'b1111111111110110;
        weights1[40433] <= 16'b1111111111110111;
        weights1[40434] <= 16'b1111111111111111;
        weights1[40435] <= 16'b1111111111110011;
        weights1[40436] <= 16'b1111111111111111;
        weights1[40437] <= 16'b0000000000010000;
        weights1[40438] <= 16'b0000000000010001;
        weights1[40439] <= 16'b0000000000001110;
        weights1[40440] <= 16'b1111111111111110;
        weights1[40441] <= 16'b1111111111110001;
        weights1[40442] <= 16'b1111111111101111;
        weights1[40443] <= 16'b1111111111110100;
        weights1[40444] <= 16'b1111111111110111;
        weights1[40445] <= 16'b1111111111111100;
        weights1[40446] <= 16'b1111111111111101;
        weights1[40447] <= 16'b0000000000000000;
        weights1[40448] <= 16'b1111111111101111;
        weights1[40449] <= 16'b1111111111101011;
        weights1[40450] <= 16'b1111111111101000;
        weights1[40451] <= 16'b1111111111010111;
        weights1[40452] <= 16'b1111111111101100;
        weights1[40453] <= 16'b1111111111111110;
        weights1[40454] <= 16'b0000000000001000;
        weights1[40455] <= 16'b0000000000010011;
        weights1[40456] <= 16'b0000000000011001;
        weights1[40457] <= 16'b0000000000001010;
        weights1[40458] <= 16'b0000000000000110;
        weights1[40459] <= 16'b0000000000001011;
        weights1[40460] <= 16'b1111111111111100;
        weights1[40461] <= 16'b1111111111110100;
        weights1[40462] <= 16'b1111111111110111;
        weights1[40463] <= 16'b1111111111110010;
        weights1[40464] <= 16'b1111111111111011;
        weights1[40465] <= 16'b0000000000000111;
        weights1[40466] <= 16'b0000000000001010;
        weights1[40467] <= 16'b0000000000010001;
        weights1[40468] <= 16'b0000000000001000;
        weights1[40469] <= 16'b0000000000001000;
        weights1[40470] <= 16'b0000000000000000;
        weights1[40471] <= 16'b0000000000000000;
        weights1[40472] <= 16'b1111111111101111;
        weights1[40473] <= 16'b1111111111110101;
        weights1[40474] <= 16'b0000000000000100;
        weights1[40475] <= 16'b0000000000001100;
        weights1[40476] <= 16'b1111111111111010;
        weights1[40477] <= 16'b1111111111100001;
        weights1[40478] <= 16'b1111111111100101;
        weights1[40479] <= 16'b1111111111100001;
        weights1[40480] <= 16'b1111111111101011;
        weights1[40481] <= 16'b1111111111110111;
        weights1[40482] <= 16'b0000000000010001;
        weights1[40483] <= 16'b0000000000010011;
        weights1[40484] <= 16'b0000000000100001;
        weights1[40485] <= 16'b1111111111111110;
        weights1[40486] <= 16'b0000000000000010;
        weights1[40487] <= 16'b0000000000001000;
        weights1[40488] <= 16'b1111111111110101;
        weights1[40489] <= 16'b1111111111110100;
        weights1[40490] <= 16'b1111111111111011;
        weights1[40491] <= 16'b1111111111110000;
        weights1[40492] <= 16'b1111111111110000;
        weights1[40493] <= 16'b1111111111111100;
        weights1[40494] <= 16'b0000000000001100;
        weights1[40495] <= 16'b0000000000001010;
        weights1[40496] <= 16'b0000000000001110;
        weights1[40497] <= 16'b0000000000001101;
        weights1[40498] <= 16'b0000000000000011;
        weights1[40499] <= 16'b1111111111111011;
        weights1[40500] <= 16'b0000000000000001;
        weights1[40501] <= 16'b0000000000001000;
        weights1[40502] <= 16'b0000000000001011;
        weights1[40503] <= 16'b0000000000000001;
        weights1[40504] <= 16'b0000000000000100;
        weights1[40505] <= 16'b1111111111100111;
        weights1[40506] <= 16'b1111111111011000;
        weights1[40507] <= 16'b1111111111010111;
        weights1[40508] <= 16'b1111111111101000;
        weights1[40509] <= 16'b1111111111111001;
        weights1[40510] <= 16'b0000000000001011;
        weights1[40511] <= 16'b0000000000011000;
        weights1[40512] <= 16'b0000000000010101;
        weights1[40513] <= 16'b0000000000000101;
        weights1[40514] <= 16'b0000000000001001;
        weights1[40515] <= 16'b0000000000000011;
        weights1[40516] <= 16'b1111111111110100;
        weights1[40517] <= 16'b1111111111101100;
        weights1[40518] <= 16'b1111111111110011;
        weights1[40519] <= 16'b1111111111101111;
        weights1[40520] <= 16'b1111111111101101;
        weights1[40521] <= 16'b0000000000000001;
        weights1[40522] <= 16'b0000000000001110;
        weights1[40523] <= 16'b0000000000011001;
        weights1[40524] <= 16'b0000000000010111;
        weights1[40525] <= 16'b0000000000001001;
        weights1[40526] <= 16'b1111111111111100;
        weights1[40527] <= 16'b1111111111111000;
        weights1[40528] <= 16'b1111111111111000;
        weights1[40529] <= 16'b0000000000001010;
        weights1[40530] <= 16'b0000000000010010;
        weights1[40531] <= 16'b0000000000010010;
        weights1[40532] <= 16'b0000000000001011;
        weights1[40533] <= 16'b1111111111101000;
        weights1[40534] <= 16'b1111111111011001;
        weights1[40535] <= 16'b1111111111100100;
        weights1[40536] <= 16'b1111111111110100;
        weights1[40537] <= 16'b1111111111110101;
        weights1[40538] <= 16'b0000000000000110;
        weights1[40539] <= 16'b0000000000001110;
        weights1[40540] <= 16'b0000000000010001;
        weights1[40541] <= 16'b0000000000000110;
        weights1[40542] <= 16'b0000000000000010;
        weights1[40543] <= 16'b1111111111110110;
        weights1[40544] <= 16'b1111111111110100;
        weights1[40545] <= 16'b1111111111110001;
        weights1[40546] <= 16'b1111111111110110;
        weights1[40547] <= 16'b1111111111101111;
        weights1[40548] <= 16'b1111111111110001;
        weights1[40549] <= 16'b0000000000000001;
        weights1[40550] <= 16'b0000000000001001;
        weights1[40551] <= 16'b0000000000010100;
        weights1[40552] <= 16'b0000000000001100;
        weights1[40553] <= 16'b0000000000001010;
        weights1[40554] <= 16'b1111111111111100;
        weights1[40555] <= 16'b1111111111110111;
        weights1[40556] <= 16'b1111111111111001;
        weights1[40557] <= 16'b0000000000001001;
        weights1[40558] <= 16'b0000000000001000;
        weights1[40559] <= 16'b0000000000010010;
        weights1[40560] <= 16'b1111111111111011;
        weights1[40561] <= 16'b1111111111011011;
        weights1[40562] <= 16'b1111111111101000;
        weights1[40563] <= 16'b1111111111100111;
        weights1[40564] <= 16'b1111111111110100;
        weights1[40565] <= 16'b1111111111110111;
        weights1[40566] <= 16'b0000000000000000;
        weights1[40567] <= 16'b0000000000001101;
        weights1[40568] <= 16'b0000000000010001;
        weights1[40569] <= 16'b0000000000000110;
        weights1[40570] <= 16'b1111111111111101;
        weights1[40571] <= 16'b1111111111111010;
        weights1[40572] <= 16'b1111111111110101;
        weights1[40573] <= 16'b1111111111111000;
        weights1[40574] <= 16'b1111111111110110;
        weights1[40575] <= 16'b1111111111111101;
        weights1[40576] <= 16'b1111111111110111;
        weights1[40577] <= 16'b1111111111110001;
        weights1[40578] <= 16'b1111111111110001;
        weights1[40579] <= 16'b0000000000001000;
        weights1[40580] <= 16'b0000000000001110;
        weights1[40581] <= 16'b0000000000011001;
        weights1[40582] <= 16'b0000000000000010;
        weights1[40583] <= 16'b1111111111110101;
        weights1[40584] <= 16'b0000000000000110;
        weights1[40585] <= 16'b0000000000000101;
        weights1[40586] <= 16'b0000000000000000;
        weights1[40587] <= 16'b0000000000001010;
        weights1[40588] <= 16'b1111111111100111;
        weights1[40589] <= 16'b1111111111010100;
        weights1[40590] <= 16'b1111111111011011;
        weights1[40591] <= 16'b1111111111110110;
        weights1[40592] <= 16'b0000000000000001;
        weights1[40593] <= 16'b1111111111111011;
        weights1[40594] <= 16'b1111111111111000;
        weights1[40595] <= 16'b0000000000000100;
        weights1[40596] <= 16'b0000000000001000;
        weights1[40597] <= 16'b1111111111111111;
        weights1[40598] <= 16'b1111111111110101;
        weights1[40599] <= 16'b1111111111110111;
        weights1[40600] <= 16'b0000000000000010;
        weights1[40601] <= 16'b1111111111111001;
        weights1[40602] <= 16'b1111111111110110;
        weights1[40603] <= 16'b1111111111101111;
        weights1[40604] <= 16'b1111111111100111;
        weights1[40605] <= 16'b1111111111101111;
        weights1[40606] <= 16'b1111111111111100;
        weights1[40607] <= 16'b0000000000001000;
        weights1[40608] <= 16'b0000000000001110;
        weights1[40609] <= 16'b0000000000010011;
        weights1[40610] <= 16'b0000000000010111;
        weights1[40611] <= 16'b0000000000001001;
        weights1[40612] <= 16'b0000000000000011;
        weights1[40613] <= 16'b0000000000000111;
        weights1[40614] <= 16'b0000000000000000;
        weights1[40615] <= 16'b1111111111110001;
        weights1[40616] <= 16'b1111111111101111;
        weights1[40617] <= 16'b1111111111100110;
        weights1[40618] <= 16'b1111111111101111;
        weights1[40619] <= 16'b1111111111111100;
        weights1[40620] <= 16'b1111111111111001;
        weights1[40621] <= 16'b1111111111110100;
        weights1[40622] <= 16'b1111111111111000;
        weights1[40623] <= 16'b1111111111110111;
        weights1[40624] <= 16'b1111111111111000;
        weights1[40625] <= 16'b1111111111111011;
        weights1[40626] <= 16'b1111111111110100;
        weights1[40627] <= 16'b1111111111111001;
        weights1[40628] <= 16'b0000000000000001;
        weights1[40629] <= 16'b1111111111111011;
        weights1[40630] <= 16'b1111111111110100;
        weights1[40631] <= 16'b1111111111111000;
        weights1[40632] <= 16'b1111111111101110;
        weights1[40633] <= 16'b1111111111101111;
        weights1[40634] <= 16'b1111111111101100;
        weights1[40635] <= 16'b1111111111101110;
        weights1[40636] <= 16'b1111111111110001;
        weights1[40637] <= 16'b0000000000000010;
        weights1[40638] <= 16'b0000000000001011;
        weights1[40639] <= 16'b0000000000010100;
        weights1[40640] <= 16'b0000000000001100;
        weights1[40641] <= 16'b1111111111111111;
        weights1[40642] <= 16'b1111111111110010;
        weights1[40643] <= 16'b1111111111110010;
        weights1[40644] <= 16'b1111111111111000;
        weights1[40645] <= 16'b1111111111110010;
        weights1[40646] <= 16'b1111111111110000;
        weights1[40647] <= 16'b0000000000000011;
        weights1[40648] <= 16'b1111111111111001;
        weights1[40649] <= 16'b1111111111110101;
        weights1[40650] <= 16'b1111111111101100;
        weights1[40651] <= 16'b1111111111101000;
        weights1[40652] <= 16'b1111111111101101;
        weights1[40653] <= 16'b1111111111110100;
        weights1[40654] <= 16'b1111111111110111;
        weights1[40655] <= 16'b1111111111111011;
        weights1[40656] <= 16'b1111111111111100;
        weights1[40657] <= 16'b0000000000000001;
        weights1[40658] <= 16'b1111111111110111;
        weights1[40659] <= 16'b1111111111111100;
        weights1[40660] <= 16'b1111111111110110;
        weights1[40661] <= 16'b1111111111110010;
        weights1[40662] <= 16'b1111111111100110;
        weights1[40663] <= 16'b1111111111011001;
        weights1[40664] <= 16'b1111111111100110;
        weights1[40665] <= 16'b1111111111101011;
        weights1[40666] <= 16'b1111111111111110;
        weights1[40667] <= 16'b0000000000000111;
        weights1[40668] <= 16'b0000000000000100;
        weights1[40669] <= 16'b1111111111111010;
        weights1[40670] <= 16'b1111111111110111;
        weights1[40671] <= 16'b1111111111110110;
        weights1[40672] <= 16'b1111111111111011;
        weights1[40673] <= 16'b1111111111101100;
        weights1[40674] <= 16'b1111111111110010;
        weights1[40675] <= 16'b1111111111111101;
        weights1[40676] <= 16'b1111111111110011;
        weights1[40677] <= 16'b1111111111100011;
        weights1[40678] <= 16'b1111111111101001;
        weights1[40679] <= 16'b1111111111101011;
        weights1[40680] <= 16'b1111111111110010;
        weights1[40681] <= 16'b1111111111101011;
        weights1[40682] <= 16'b1111111111111111;
        weights1[40683] <= 16'b1111111111111011;
        weights1[40684] <= 16'b1111111111111110;
        weights1[40685] <= 16'b1111111111111110;
        weights1[40686] <= 16'b1111111111111110;
        weights1[40687] <= 16'b1111111111111011;
        weights1[40688] <= 16'b1111111111111001;
        weights1[40689] <= 16'b1111111111110100;
        weights1[40690] <= 16'b1111111111110000;
        weights1[40691] <= 16'b1111111111111000;
        weights1[40692] <= 16'b1111111111110001;
        weights1[40693] <= 16'b1111111111101000;
        weights1[40694] <= 16'b1111111111101001;
        weights1[40695] <= 16'b1111111111101010;
        weights1[40696] <= 16'b1111111111101001;
        weights1[40697] <= 16'b1111111111100111;
        weights1[40698] <= 16'b1111111111110011;
        weights1[40699] <= 16'b1111111111111011;
        weights1[40700] <= 16'b1111111111111101;
        weights1[40701] <= 16'b1111111111110110;
        weights1[40702] <= 16'b1111111111110101;
        weights1[40703] <= 16'b1111111111110110;
        weights1[40704] <= 16'b1111111111101000;
        weights1[40705] <= 16'b1111111111101101;
        weights1[40706] <= 16'b1111111111101101;
        weights1[40707] <= 16'b1111111111110000;
        weights1[40708] <= 16'b1111111111100101;
        weights1[40709] <= 16'b1111111111110000;
        weights1[40710] <= 16'b1111111111111011;
        weights1[40711] <= 16'b1111111111111100;
        weights1[40712] <= 16'b0000000000000000;
        weights1[40713] <= 16'b1111111111111011;
        weights1[40714] <= 16'b1111111111111000;
        weights1[40715] <= 16'b1111111111110111;
        weights1[40716] <= 16'b1111111111111011;
        weights1[40717] <= 16'b0000000000000011;
        weights1[40718] <= 16'b1111111111111111;
        weights1[40719] <= 16'b0000000000000010;
        weights1[40720] <= 16'b0000000000000100;
        weights1[40721] <= 16'b1111111111111100;
        weights1[40722] <= 16'b1111111111110001;
        weights1[40723] <= 16'b1111111111111100;
        weights1[40724] <= 16'b1111111111111000;
        weights1[40725] <= 16'b1111111111111010;
        weights1[40726] <= 16'b1111111111110111;
        weights1[40727] <= 16'b1111111111111111;
        weights1[40728] <= 16'b0000000000000011;
        weights1[40729] <= 16'b1111111111111100;
        weights1[40730] <= 16'b1111111111110100;
        weights1[40731] <= 16'b1111111111110011;
        weights1[40732] <= 16'b1111111111100111;
        weights1[40733] <= 16'b1111111111100111;
        weights1[40734] <= 16'b1111111111101110;
        weights1[40735] <= 16'b1111111111101101;
        weights1[40736] <= 16'b1111111111101110;
        weights1[40737] <= 16'b1111111111110100;
        weights1[40738] <= 16'b1111111111111001;
        weights1[40739] <= 16'b1111111111111101;
        weights1[40740] <= 16'b1111111111111110;
        weights1[40741] <= 16'b1111111111111010;
        weights1[40742] <= 16'b1111111111111001;
        weights1[40743] <= 16'b1111111111110101;
        weights1[40744] <= 16'b1111111111110000;
        weights1[40745] <= 16'b1111111111110110;
        weights1[40746] <= 16'b1111111111111010;
        weights1[40747] <= 16'b1111111111111111;
        weights1[40748] <= 16'b1111111111111000;
        weights1[40749] <= 16'b0000000000000000;
        weights1[40750] <= 16'b1111111111111011;
        weights1[40751] <= 16'b0000000000000111;
        weights1[40752] <= 16'b0000000000000000;
        weights1[40753] <= 16'b0000000000000010;
        weights1[40754] <= 16'b0000000000000010;
        weights1[40755] <= 16'b0000000000001111;
        weights1[40756] <= 16'b0000000000001001;
        weights1[40757] <= 16'b1111111111111011;
        weights1[40758] <= 16'b1111111111111000;
        weights1[40759] <= 16'b1111111111110010;
        weights1[40760] <= 16'b1111111111101000;
        weights1[40761] <= 16'b1111111111101010;
        weights1[40762] <= 16'b1111111111101101;
        weights1[40763] <= 16'b1111111111110000;
        weights1[40764] <= 16'b1111111111110101;
        weights1[40765] <= 16'b1111111111111100;
        weights1[40766] <= 16'b1111111111111101;
        weights1[40767] <= 16'b1111111111111110;
        weights1[40768] <= 16'b1111111111111111;
        weights1[40769] <= 16'b1111111111111111;
        weights1[40770] <= 16'b1111111111111111;
        weights1[40771] <= 16'b1111111111111111;
        weights1[40772] <= 16'b0000000000000001;
        weights1[40773] <= 16'b0000000000000011;
        weights1[40774] <= 16'b0000000000000010;
        weights1[40775] <= 16'b0000000000000100;
        weights1[40776] <= 16'b0000000000010011;
        weights1[40777] <= 16'b0000000000011010;
        weights1[40778] <= 16'b0000000000100101;
        weights1[40779] <= 16'b0000000000110101;
        weights1[40780] <= 16'b0000000000111000;
        weights1[40781] <= 16'b0000000001000100;
        weights1[40782] <= 16'b0000000001001111;
        weights1[40783] <= 16'b0000000001001001;
        weights1[40784] <= 16'b0000000000110010;
        weights1[40785] <= 16'b0000000000101100;
        weights1[40786] <= 16'b0000000000100010;
        weights1[40787] <= 16'b0000000000100111;
        weights1[40788] <= 16'b0000000000100001;
        weights1[40789] <= 16'b0000000000010111;
        weights1[40790] <= 16'b0000000000010000;
        weights1[40791] <= 16'b0000000000010010;
        weights1[40792] <= 16'b0000000000001100;
        weights1[40793] <= 16'b0000000000000111;
        weights1[40794] <= 16'b0000000000000101;
        weights1[40795] <= 16'b0000000000000001;
        weights1[40796] <= 16'b0000000000000000;
        weights1[40797] <= 16'b1111111111111111;
        weights1[40798] <= 16'b1111111111111111;
        weights1[40799] <= 16'b1111111111111111;
        weights1[40800] <= 16'b1111111111111111;
        weights1[40801] <= 16'b1111111111111001;
        weights1[40802] <= 16'b1111111111111011;
        weights1[40803] <= 16'b0000000000000111;
        weights1[40804] <= 16'b0000000000010111;
        weights1[40805] <= 16'b0000000000011000;
        weights1[40806] <= 16'b0000000000100010;
        weights1[40807] <= 16'b0000000000101010;
        weights1[40808] <= 16'b0000000001000011;
        weights1[40809] <= 16'b0000000001010000;
        weights1[40810] <= 16'b0000000001000110;
        weights1[40811] <= 16'b0000000000111011;
        weights1[40812] <= 16'b0000000000110010;
        weights1[40813] <= 16'b0000000000111111;
        weights1[40814] <= 16'b0000000000100010;
        weights1[40815] <= 16'b0000000000011011;
        weights1[40816] <= 16'b0000000000011100;
        weights1[40817] <= 16'b0000000000011110;
        weights1[40818] <= 16'b0000000000011010;
        weights1[40819] <= 16'b0000000000011011;
        weights1[40820] <= 16'b0000000000001111;
        weights1[40821] <= 16'b0000000000001110;
        weights1[40822] <= 16'b0000000000001010;
        weights1[40823] <= 16'b0000000000000100;
        weights1[40824] <= 16'b1111111111111111;
        weights1[40825] <= 16'b1111111111111111;
        weights1[40826] <= 16'b1111111111111110;
        weights1[40827] <= 16'b1111111111111011;
        weights1[40828] <= 16'b1111111111111011;
        weights1[40829] <= 16'b1111111111110101;
        weights1[40830] <= 16'b1111111111110101;
        weights1[40831] <= 16'b1111111111111111;
        weights1[40832] <= 16'b0000000000000011;
        weights1[40833] <= 16'b1111111111111110;
        weights1[40834] <= 16'b0000000000001001;
        weights1[40835] <= 16'b0000000000001110;
        weights1[40836] <= 16'b0000000000010110;
        weights1[40837] <= 16'b0000000000111010;
        weights1[40838] <= 16'b0000000000101111;
        weights1[40839] <= 16'b0000000000111011;
        weights1[40840] <= 16'b0000000000111111;
        weights1[40841] <= 16'b0000000000110101;
        weights1[40842] <= 16'b0000000000100010;
        weights1[40843] <= 16'b0000000000101000;
        weights1[40844] <= 16'b0000000000011110;
        weights1[40845] <= 16'b0000000000110011;
        weights1[40846] <= 16'b0000000000010011;
        weights1[40847] <= 16'b0000000000011011;
        weights1[40848] <= 16'b0000000000010001;
        weights1[40849] <= 16'b0000000000001000;
        weights1[40850] <= 16'b0000000000001000;
        weights1[40851] <= 16'b0000000000001001;
        weights1[40852] <= 16'b1111111111111101;
        weights1[40853] <= 16'b1111111111111101;
        weights1[40854] <= 16'b1111111111111100;
        weights1[40855] <= 16'b1111111111110101;
        weights1[40856] <= 16'b1111111111101111;
        weights1[40857] <= 16'b1111111111101100;
        weights1[40858] <= 16'b1111111111100001;
        weights1[40859] <= 16'b1111111111100101;
        weights1[40860] <= 16'b1111111111101110;
        weights1[40861] <= 16'b1111111111101000;
        weights1[40862] <= 16'b1111111111100010;
        weights1[40863] <= 16'b1111111111101010;
        weights1[40864] <= 16'b1111111111110000;
        weights1[40865] <= 16'b0000000000000101;
        weights1[40866] <= 16'b0000000000010100;
        weights1[40867] <= 16'b0000000000011011;
        weights1[40868] <= 16'b0000000000101011;
        weights1[40869] <= 16'b0000000000100101;
        weights1[40870] <= 16'b0000000000110101;
        weights1[40871] <= 16'b0000000000101000;
        weights1[40872] <= 16'b0000000000100101;
        weights1[40873] <= 16'b0000000000100111;
        weights1[40874] <= 16'b0000000000001110;
        weights1[40875] <= 16'b0000000000010111;
        weights1[40876] <= 16'b0000000000001000;
        weights1[40877] <= 16'b0000000000001001;
        weights1[40878] <= 16'b0000000000001100;
        weights1[40879] <= 16'b0000000000000110;
        weights1[40880] <= 16'b1111111111111011;
        weights1[40881] <= 16'b1111111111111101;
        weights1[40882] <= 16'b1111111111110000;
        weights1[40883] <= 16'b1111111111110001;
        weights1[40884] <= 16'b1111111111100011;
        weights1[40885] <= 16'b1111111111011101;
        weights1[40886] <= 16'b1111111111010001;
        weights1[40887] <= 16'b1111111111010000;
        weights1[40888] <= 16'b1111111111001110;
        weights1[40889] <= 16'b1111111110111011;
        weights1[40890] <= 16'b1111111110110011;
        weights1[40891] <= 16'b1111111110111101;
        weights1[40892] <= 16'b1111111111001001;
        weights1[40893] <= 16'b1111111111001111;
        weights1[40894] <= 16'b1111111111010110;
        weights1[40895] <= 16'b1111111111110001;
        weights1[40896] <= 16'b1111111111111001;
        weights1[40897] <= 16'b0000000000000111;
        weights1[40898] <= 16'b0000000000001111;
        weights1[40899] <= 16'b0000000000010100;
        weights1[40900] <= 16'b0000000000011010;
        weights1[40901] <= 16'b0000000000001011;
        weights1[40902] <= 16'b0000000000011011;
        weights1[40903] <= 16'b0000000000010110;
        weights1[40904] <= 16'b0000000000011010;
        weights1[40905] <= 16'b1111111111111001;
        weights1[40906] <= 16'b1111111111111111;
        weights1[40907] <= 16'b0000000000001000;
        weights1[40908] <= 16'b1111111111111100;
        weights1[40909] <= 16'b1111111111110001;
        weights1[40910] <= 16'b1111111111100001;
        weights1[40911] <= 16'b1111111111011000;
        weights1[40912] <= 16'b1111111111001100;
        weights1[40913] <= 16'b1111111111001100;
        weights1[40914] <= 16'b1111111110111000;
        weights1[40915] <= 16'b1111111110100111;
        weights1[40916] <= 16'b1111111110101010;
        weights1[40917] <= 16'b1111111110100100;
        weights1[40918] <= 16'b1111111110100101;
        weights1[40919] <= 16'b1111111110101000;
        weights1[40920] <= 16'b1111111110110000;
        weights1[40921] <= 16'b1111111110101110;
        weights1[40922] <= 16'b1111111110110111;
        weights1[40923] <= 16'b1111111110111011;
        weights1[40924] <= 16'b1111111111001111;
        weights1[40925] <= 16'b1111111111011010;
        weights1[40926] <= 16'b1111111111010111;
        weights1[40927] <= 16'b1111111111101010;
        weights1[40928] <= 16'b0000000000000011;
        weights1[40929] <= 16'b1111111111101100;
        weights1[40930] <= 16'b0000000000000011;
        weights1[40931] <= 16'b0000000000001111;
        weights1[40932] <= 16'b0000000000010010;
        weights1[40933] <= 16'b0000000000000111;
        weights1[40934] <= 16'b0000000000001100;
        weights1[40935] <= 16'b0000000000000111;
        weights1[40936] <= 16'b1111111111111000;
        weights1[40937] <= 16'b1111111111101110;
        weights1[40938] <= 16'b1111111111101001;
        weights1[40939] <= 16'b1111111111010110;
        weights1[40940] <= 16'b1111111111000101;
        weights1[40941] <= 16'b1111111110111110;
        weights1[40942] <= 16'b1111111110011011;
        weights1[40943] <= 16'b1111111110000110;
        weights1[40944] <= 16'b1111111110010010;
        weights1[40945] <= 16'b1111111110000011;
        weights1[40946] <= 16'b1111111110000110;
        weights1[40947] <= 16'b1111111110001010;
        weights1[40948] <= 16'b1111111110010111;
        weights1[40949] <= 16'b1111111110011011;
        weights1[40950] <= 16'b1111111110100000;
        weights1[40951] <= 16'b1111111110101000;
        weights1[40952] <= 16'b1111111110110011;
        weights1[40953] <= 16'b1111111110110111;
        weights1[40954] <= 16'b1111111111001101;
        weights1[40955] <= 16'b1111111111010111;
        weights1[40956] <= 16'b1111111111100010;
        weights1[40957] <= 16'b1111111111110110;
        weights1[40958] <= 16'b1111111111101000;
        weights1[40959] <= 16'b0000000000001000;
        weights1[40960] <= 16'b0000000000001011;
        weights1[40961] <= 16'b0000000000000001;
        weights1[40962] <= 16'b0000000000001000;
        weights1[40963] <= 16'b0000000000001010;
        weights1[40964] <= 16'b1111111111111000;
        weights1[40965] <= 16'b1111111111101111;
        weights1[40966] <= 16'b1111111111101101;
        weights1[40967] <= 16'b1111111111100001;
        weights1[40968] <= 16'b1111111111011100;
        weights1[40969] <= 16'b1111111111011111;
        weights1[40970] <= 16'b1111111111001001;
        weights1[40971] <= 16'b1111111110111110;
        weights1[40972] <= 16'b1111111111000100;
        weights1[40973] <= 16'b1111111110101111;
        weights1[40974] <= 16'b1111111110100110;
        weights1[40975] <= 16'b1111111110010011;
        weights1[40976] <= 16'b1111111110011000;
        weights1[40977] <= 16'b1111111110011100;
        weights1[40978] <= 16'b1111111110110110;
        weights1[40979] <= 16'b1111111110110111;
        weights1[40980] <= 16'b1111111110101010;
        weights1[40981] <= 16'b1111111110100111;
        weights1[40982] <= 16'b1111111111001100;
        weights1[40983] <= 16'b1111111111100000;
        weights1[40984] <= 16'b1111111111101100;
        weights1[40985] <= 16'b1111111111011000;
        weights1[40986] <= 16'b1111111111110100;
        weights1[40987] <= 16'b0000000000010010;
        weights1[40988] <= 16'b0000000000001100;
        weights1[40989] <= 16'b1111111111111111;
        weights1[40990] <= 16'b0000000000000110;
        weights1[40991] <= 16'b1111111111111110;
        weights1[40992] <= 16'b1111111111111011;
        weights1[40993] <= 16'b1111111111111000;
        weights1[40994] <= 16'b1111111111110110;
        weights1[40995] <= 16'b1111111111110111;
        weights1[40996] <= 16'b1111111111111111;
        weights1[40997] <= 16'b0000000000000001;
        weights1[40998] <= 16'b0000000000001011;
        weights1[40999] <= 16'b1111111111110000;
        weights1[41000] <= 16'b1111111111011101;
        weights1[41001] <= 16'b1111111111110010;
        weights1[41002] <= 16'b1111111110111111;
        weights1[41003] <= 16'b1111111111000111;
        weights1[41004] <= 16'b1111111110101101;
        weights1[41005] <= 16'b1111111111000011;
        weights1[41006] <= 16'b1111111111001110;
        weights1[41007] <= 16'b1111111111000001;
        weights1[41008] <= 16'b1111111111011011;
        weights1[41009] <= 16'b1111111111101001;
        weights1[41010] <= 16'b1111111111100111;
        weights1[41011] <= 16'b1111111111100000;
        weights1[41012] <= 16'b1111111111111101;
        weights1[41013] <= 16'b0000000000000011;
        weights1[41014] <= 16'b1111111111101110;
        weights1[41015] <= 16'b1111111111111100;
        weights1[41016] <= 16'b1111111111111100;
        weights1[41017] <= 16'b0000000000000111;
        weights1[41018] <= 16'b1111111111101001;
        weights1[41019] <= 16'b1111111111110110;
        weights1[41020] <= 16'b0000000000000110;
        weights1[41021] <= 16'b1111111111111011;
        weights1[41022] <= 16'b0000000000001010;
        weights1[41023] <= 16'b0000000000011001;
        weights1[41024] <= 16'b0000000000101011;
        weights1[41025] <= 16'b0000000000011100;
        weights1[41026] <= 16'b0000000000100000;
        weights1[41027] <= 16'b0000000000011000;
        weights1[41028] <= 16'b0000000000001000;
        weights1[41029] <= 16'b1111111111110111;
        weights1[41030] <= 16'b1111111111110111;
        weights1[41031] <= 16'b1111111111100101;
        weights1[41032] <= 16'b1111111111101111;
        weights1[41033] <= 16'b1111111111011111;
        weights1[41034] <= 16'b1111111111110011;
        weights1[41035] <= 16'b1111111111111010;
        weights1[41036] <= 16'b0000000000001111;
        weights1[41037] <= 16'b0000000000001001;
        weights1[41038] <= 16'b0000000000000010;
        weights1[41039] <= 16'b1111111111110000;
        weights1[41040] <= 16'b1111111111110101;
        weights1[41041] <= 16'b0000000000000100;
        weights1[41042] <= 16'b1111111111111011;
        weights1[41043] <= 16'b1111111111111000;
        weights1[41044] <= 16'b1111111111111100;
        weights1[41045] <= 16'b1111111111110000;
        weights1[41046] <= 16'b1111111111110110;
        weights1[41047] <= 16'b1111111111111110;
        weights1[41048] <= 16'b0000000000001111;
        weights1[41049] <= 16'b0000000000010001;
        weights1[41050] <= 16'b0000000000100110;
        weights1[41051] <= 16'b0000000000101100;
        weights1[41052] <= 16'b0000000000101000;
        weights1[41053] <= 16'b0000000000100101;
        weights1[41054] <= 16'b0000000000011110;
        weights1[41055] <= 16'b0000000000101110;
        weights1[41056] <= 16'b0000000000101010;
        weights1[41057] <= 16'b0000000000100100;
        weights1[41058] <= 16'b0000000000001111;
        weights1[41059] <= 16'b0000000000011001;
        weights1[41060] <= 16'b0000000000011011;
        weights1[41061] <= 16'b1111111111111000;
        weights1[41062] <= 16'b0000000000000000;
        weights1[41063] <= 16'b1111111111110010;
        weights1[41064] <= 16'b1111111111110110;
        weights1[41065] <= 16'b1111111111111100;
        weights1[41066] <= 16'b0000000000000001;
        weights1[41067] <= 16'b0000000000001100;
        weights1[41068] <= 16'b0000000000001100;
        weights1[41069] <= 16'b1111111111111110;
        weights1[41070] <= 16'b0000000000010101;
        weights1[41071] <= 16'b0000000000001011;
        weights1[41072] <= 16'b1111111111111011;
        weights1[41073] <= 16'b1111111111111100;
        weights1[41074] <= 16'b0000000000000101;
        weights1[41075] <= 16'b1111111111111000;
        weights1[41076] <= 16'b0000000000010101;
        weights1[41077] <= 16'b0000000000011110;
        weights1[41078] <= 16'b0000000000101010;
        weights1[41079] <= 16'b0000000000100000;
        weights1[41080] <= 16'b0000000000100001;
        weights1[41081] <= 16'b0000000000010111;
        weights1[41082] <= 16'b0000000000011101;
        weights1[41083] <= 16'b0000000000001011;
        weights1[41084] <= 16'b0000000000101010;
        weights1[41085] <= 16'b0000000000011100;
        weights1[41086] <= 16'b0000000000100100;
        weights1[41087] <= 16'b0000000000011101;
        weights1[41088] <= 16'b0000000000011101;
        weights1[41089] <= 16'b0000000000001111;
        weights1[41090] <= 16'b0000000000100011;
        weights1[41091] <= 16'b0000000000011001;
        weights1[41092] <= 16'b0000000000010011;
        weights1[41093] <= 16'b0000000000000010;
        weights1[41094] <= 16'b0000000000011010;
        weights1[41095] <= 16'b1111111111111101;
        weights1[41096] <= 16'b0000000000001001;
        weights1[41097] <= 16'b0000000000010000;
        weights1[41098] <= 16'b0000000000000001;
        weights1[41099] <= 16'b0000000000000001;
        weights1[41100] <= 16'b1111111111100101;
        weights1[41101] <= 16'b0000000000000111;
        weights1[41102] <= 16'b0000000000001010;
        weights1[41103] <= 16'b1111111111101111;
        weights1[41104] <= 16'b0000000000011010;
        weights1[41105] <= 16'b0000000000010111;
        weights1[41106] <= 16'b0000000000011100;
        weights1[41107] <= 16'b0000000000001111;
        weights1[41108] <= 16'b1111111111110011;
        weights1[41109] <= 16'b0000000000000110;
        weights1[41110] <= 16'b0000000000001001;
        weights1[41111] <= 16'b0000000000011110;
        weights1[41112] <= 16'b0000000000110011;
        weights1[41113] <= 16'b0000000000010010;
        weights1[41114] <= 16'b0000000000010100;
        weights1[41115] <= 16'b0000000000101101;
        weights1[41116] <= 16'b0000000000100110;
        weights1[41117] <= 16'b0000000000110011;
        weights1[41118] <= 16'b0000000000101111;
        weights1[41119] <= 16'b0000000000011011;
        weights1[41120] <= 16'b0000000000101000;
        weights1[41121] <= 16'b0000000000010110;
        weights1[41122] <= 16'b0000000000010111;
        weights1[41123] <= 16'b0000000000011000;
        weights1[41124] <= 16'b0000000000010001;
        weights1[41125] <= 16'b0000000000000011;
        weights1[41126] <= 16'b1111111111111100;
        weights1[41127] <= 16'b1111111111111101;
        weights1[41128] <= 16'b0000000000000110;
        weights1[41129] <= 16'b0000000000001000;
        weights1[41130] <= 16'b1111111111111101;
        weights1[41131] <= 16'b1111111111111100;
        weights1[41132] <= 16'b0000000000011001;
        weights1[41133] <= 16'b0000000000010111;
        weights1[41134] <= 16'b0000000000001000;
        weights1[41135] <= 16'b1111111111111000;
        weights1[41136] <= 16'b1111111111111110;
        weights1[41137] <= 16'b0000000000010100;
        weights1[41138] <= 16'b1111111111110111;
        weights1[41139] <= 16'b1111111111110110;
        weights1[41140] <= 16'b0000000000001010;
        weights1[41141] <= 16'b0000000000011010;
        weights1[41142] <= 16'b0000000000011111;
        weights1[41143] <= 16'b0000000000011111;
        weights1[41144] <= 16'b0000000000101110;
        weights1[41145] <= 16'b0000000000011111;
        weights1[41146] <= 16'b0000000000011000;
        weights1[41147] <= 16'b0000000000101100;
        weights1[41148] <= 16'b0000000000011001;
        weights1[41149] <= 16'b0000000000100100;
        weights1[41150] <= 16'b0000000000110000;
        weights1[41151] <= 16'b0000000000001010;
        weights1[41152] <= 16'b0000000000010000;
        weights1[41153] <= 16'b0000000000010110;
        weights1[41154] <= 16'b0000000000000101;
        weights1[41155] <= 16'b0000000000000011;
        weights1[41156] <= 16'b0000000000000100;
        weights1[41157] <= 16'b0000000000001100;
        weights1[41158] <= 16'b0000000000010000;
        weights1[41159] <= 16'b1111111111110010;
        weights1[41160] <= 16'b0000000000010011;
        weights1[41161] <= 16'b0000000000001100;
        weights1[41162] <= 16'b0000000000000001;
        weights1[41163] <= 16'b1111111111111111;
        weights1[41164] <= 16'b0000000000000001;
        weights1[41165] <= 16'b1111111111011111;
        weights1[41166] <= 16'b1111111111110001;
        weights1[41167] <= 16'b1111111111110010;
        weights1[41168] <= 16'b0000000000000011;
        weights1[41169] <= 16'b1111111111111001;
        weights1[41170] <= 16'b0000000000000000;
        weights1[41171] <= 16'b1111111111111111;
        weights1[41172] <= 16'b0000000000001011;
        weights1[41173] <= 16'b0000000000000010;
        weights1[41174] <= 16'b0000000000000111;
        weights1[41175] <= 16'b0000000000001100;
        weights1[41176] <= 16'b0000000000010000;
        weights1[41177] <= 16'b0000000000000010;
        weights1[41178] <= 16'b0000000000001011;
        weights1[41179] <= 16'b0000000000011011;
        weights1[41180] <= 16'b0000000000001110;
        weights1[41181] <= 16'b1111111111111000;
        weights1[41182] <= 16'b0000000000010011;
        weights1[41183] <= 16'b0000000000011001;
        weights1[41184] <= 16'b1111111111111100;
        weights1[41185] <= 16'b0000000000000111;
        weights1[41186] <= 16'b0000000000001000;
        weights1[41187] <= 16'b1111111111111111;
        weights1[41188] <= 16'b0000000000010110;
        weights1[41189] <= 16'b0000000000010011;
        weights1[41190] <= 16'b0000000000000000;
        weights1[41191] <= 16'b1111111111110011;
        weights1[41192] <= 16'b1111111111100011;
        weights1[41193] <= 16'b1111111111110000;
        weights1[41194] <= 16'b0000000000000101;
        weights1[41195] <= 16'b1111111111111000;
        weights1[41196] <= 16'b1111111111110111;
        weights1[41197] <= 16'b1111111111111110;
        weights1[41198] <= 16'b1111111111111110;
        weights1[41199] <= 16'b1111111111110000;
        weights1[41200] <= 16'b1111111111100000;
        weights1[41201] <= 16'b1111111111100111;
        weights1[41202] <= 16'b1111111111100111;
        weights1[41203] <= 16'b1111111111011001;
        weights1[41204] <= 16'b1111111111011011;
        weights1[41205] <= 16'b1111111111110011;
        weights1[41206] <= 16'b1111111111111000;
        weights1[41207] <= 16'b1111111111110110;
        weights1[41208] <= 16'b0000000000000110;
        weights1[41209] <= 16'b1111111111110111;
        weights1[41210] <= 16'b1111111111111111;
        weights1[41211] <= 16'b1111111111110111;
        weights1[41212] <= 16'b0000000000001011;
        weights1[41213] <= 16'b0000000000001010;
        weights1[41214] <= 16'b1111111111111110;
        weights1[41215] <= 16'b0000000000010001;
        weights1[41216] <= 16'b0000000000001010;
        weights1[41217] <= 16'b0000000000000111;
        weights1[41218] <= 16'b0000000000000100;
        weights1[41219] <= 16'b0000000000000001;
        weights1[41220] <= 16'b1111111111111110;
        weights1[41221] <= 16'b1111111111111010;
        weights1[41222] <= 16'b1111111111110100;
        weights1[41223] <= 16'b1111111111111111;
        weights1[41224] <= 16'b0000000000000111;
        weights1[41225] <= 16'b1111111111101100;
        weights1[41226] <= 16'b1111111111011110;
        weights1[41227] <= 16'b1111111111110111;
        weights1[41228] <= 16'b1111111111011001;
        weights1[41229] <= 16'b1111111111010111;
        weights1[41230] <= 16'b1111111111010011;
        weights1[41231] <= 16'b1111111111010000;
        weights1[41232] <= 16'b1111111111011010;
        weights1[41233] <= 16'b1111111111011110;
        weights1[41234] <= 16'b1111111111101000;
        weights1[41235] <= 16'b1111111111110111;
        weights1[41236] <= 16'b1111111111110100;
        weights1[41237] <= 16'b1111111111110010;
        weights1[41238] <= 16'b1111111111111001;
        weights1[41239] <= 16'b1111111111110000;
        weights1[41240] <= 16'b1111111111111001;
        weights1[41241] <= 16'b0000000000000001;
        weights1[41242] <= 16'b0000000000000011;
        weights1[41243] <= 16'b0000000000011000;
        weights1[41244] <= 16'b0000000000000100;
        weights1[41245] <= 16'b0000000000000110;
        weights1[41246] <= 16'b1111111111110100;
        weights1[41247] <= 16'b1111111111111010;
        weights1[41248] <= 16'b0000000000001101;
        weights1[41249] <= 16'b1111111111111001;
        weights1[41250] <= 16'b0000000000011001;
        weights1[41251] <= 16'b1111111111111010;
        weights1[41252] <= 16'b1111111111101010;
        weights1[41253] <= 16'b1111111111100100;
        weights1[41254] <= 16'b1111111111011110;
        weights1[41255] <= 16'b1111111111011100;
        weights1[41256] <= 16'b1111111111010101;
        weights1[41257] <= 16'b1111111111010101;
        weights1[41258] <= 16'b1111111111100000;
        weights1[41259] <= 16'b1111111111010111;
        weights1[41260] <= 16'b1111111111011000;
        weights1[41261] <= 16'b1111111111010111;
        weights1[41262] <= 16'b1111111111100000;
        weights1[41263] <= 16'b1111111111001011;
        weights1[41264] <= 16'b1111111111101010;
        weights1[41265] <= 16'b1111111111110010;
        weights1[41266] <= 16'b0000000000001000;
        weights1[41267] <= 16'b1111111111101101;
        weights1[41268] <= 16'b0000000000010010;
        weights1[41269] <= 16'b0000000000000001;
        weights1[41270] <= 16'b0000000000000010;
        weights1[41271] <= 16'b0000000000010111;
        weights1[41272] <= 16'b1111111111111110;
        weights1[41273] <= 16'b1111111111111001;
        weights1[41274] <= 16'b1111111111101110;
        weights1[41275] <= 16'b1111111111110011;
        weights1[41276] <= 16'b1111111111111010;
        weights1[41277] <= 16'b1111111111110101;
        weights1[41278] <= 16'b0000000000000000;
        weights1[41279] <= 16'b1111111111100001;
        weights1[41280] <= 16'b1111111111100110;
        weights1[41281] <= 16'b1111111111010111;
        weights1[41282] <= 16'b1111111111010011;
        weights1[41283] <= 16'b1111111111010111;
        weights1[41284] <= 16'b1111111111011011;
        weights1[41285] <= 16'b1111111111011011;
        weights1[41286] <= 16'b1111111111101011;
        weights1[41287] <= 16'b1111111111010011;
        weights1[41288] <= 16'b1111111111100010;
        weights1[41289] <= 16'b1111111111101011;
        weights1[41290] <= 16'b1111111111100100;
        weights1[41291] <= 16'b1111111111011100;
        weights1[41292] <= 16'b1111111111110010;
        weights1[41293] <= 16'b0000000000001000;
        weights1[41294] <= 16'b1111111111101101;
        weights1[41295] <= 16'b0000000000001000;
        weights1[41296] <= 16'b0000000000010010;
        weights1[41297] <= 16'b0000000000000100;
        weights1[41298] <= 16'b0000000000011001;
        weights1[41299] <= 16'b0000000000010000;
        weights1[41300] <= 16'b0000000000000001;
        weights1[41301] <= 16'b1111111111110111;
        weights1[41302] <= 16'b1111111111111010;
        weights1[41303] <= 16'b1111111111111000;
        weights1[41304] <= 16'b1111111111101010;
        weights1[41305] <= 16'b1111111111101111;
        weights1[41306] <= 16'b1111111111101000;
        weights1[41307] <= 16'b1111111111011000;
        weights1[41308] <= 16'b1111111111100000;
        weights1[41309] <= 16'b1111111111011101;
        weights1[41310] <= 16'b1111111111001101;
        weights1[41311] <= 16'b1111111111001101;
        weights1[41312] <= 16'b1111111111011100;
        weights1[41313] <= 16'b1111111111100101;
        weights1[41314] <= 16'b1111111111010111;
        weights1[41315] <= 16'b1111111111101000;
        weights1[41316] <= 16'b1111111111101111;
        weights1[41317] <= 16'b0000000000000000;
        weights1[41318] <= 16'b1111111111011101;
        weights1[41319] <= 16'b1111111111111100;
        weights1[41320] <= 16'b1111111111111111;
        weights1[41321] <= 16'b1111111111111111;
        weights1[41322] <= 16'b0000000000001000;
        weights1[41323] <= 16'b0000000000001111;
        weights1[41324] <= 16'b0000000000001000;
        weights1[41325] <= 16'b0000000000000110;
        weights1[41326] <= 16'b0000000000010101;
        weights1[41327] <= 16'b0000000000011100;
        weights1[41328] <= 16'b0000000000000110;
        weights1[41329] <= 16'b0000000000001001;
        weights1[41330] <= 16'b1111111111111100;
        weights1[41331] <= 16'b1111111111110100;
        weights1[41332] <= 16'b1111111111100011;
        weights1[41333] <= 16'b1111111111101100;
        weights1[41334] <= 16'b1111111111110011;
        weights1[41335] <= 16'b1111111111110010;
        weights1[41336] <= 16'b1111111111011111;
        weights1[41337] <= 16'b1111111111101010;
        weights1[41338] <= 16'b1111111111100111;
        weights1[41339] <= 16'b1111111111100011;
        weights1[41340] <= 16'b1111111111100011;
        weights1[41341] <= 16'b1111111111011110;
        weights1[41342] <= 16'b1111111111101001;
        weights1[41343] <= 16'b0000000000000000;
        weights1[41344] <= 16'b1111111111101010;
        weights1[41345] <= 16'b1111111111101010;
        weights1[41346] <= 16'b1111111111111100;
        weights1[41347] <= 16'b0000000000000011;
        weights1[41348] <= 16'b0000000000010011;
        weights1[41349] <= 16'b0000000000000000;
        weights1[41350] <= 16'b0000000000010010;
        weights1[41351] <= 16'b0000000000001010;
        weights1[41352] <= 16'b0000000000000111;
        weights1[41353] <= 16'b0000000000001000;
        weights1[41354] <= 16'b0000000000010101;
        weights1[41355] <= 16'b0000000000010000;
        weights1[41356] <= 16'b0000000000000111;
        weights1[41357] <= 16'b1111111111111110;
        weights1[41358] <= 16'b1111111111111001;
        weights1[41359] <= 16'b1111111111111000;
        weights1[41360] <= 16'b1111111111111100;
        weights1[41361] <= 16'b0000000000001011;
        weights1[41362] <= 16'b1111111111111010;
        weights1[41363] <= 16'b1111111111110011;
        weights1[41364] <= 16'b1111111111110111;
        weights1[41365] <= 16'b1111111111101110;
        weights1[41366] <= 16'b1111111111011110;
        weights1[41367] <= 16'b1111111111100110;
        weights1[41368] <= 16'b1111111111100011;
        weights1[41369] <= 16'b1111111111101010;
        weights1[41370] <= 16'b1111111111110110;
        weights1[41371] <= 16'b1111111111101000;
        weights1[41372] <= 16'b1111111111110010;
        weights1[41373] <= 16'b0000000000000101;
        weights1[41374] <= 16'b1111111111111100;
        weights1[41375] <= 16'b1111111111111111;
        weights1[41376] <= 16'b0000000000100010;
        weights1[41377] <= 16'b0000000000001000;
        weights1[41378] <= 16'b0000000000001101;
        weights1[41379] <= 16'b0000000000010110;
        weights1[41380] <= 16'b1111111111111100;
        weights1[41381] <= 16'b0000000000000111;
        weights1[41382] <= 16'b0000000000001101;
        weights1[41383] <= 16'b0000000000010010;
        weights1[41384] <= 16'b0000000000001000;
        weights1[41385] <= 16'b0000000000000000;
        weights1[41386] <= 16'b0000000000001010;
        weights1[41387] <= 16'b0000000000000011;
        weights1[41388] <= 16'b0000000000001010;
        weights1[41389] <= 16'b0000000000001111;
        weights1[41390] <= 16'b1111111111111010;
        weights1[41391] <= 16'b0000000000000110;
        weights1[41392] <= 16'b0000000000001011;
        weights1[41393] <= 16'b0000000000010100;
        weights1[41394] <= 16'b1111111111111001;
        weights1[41395] <= 16'b0000000000010101;
        weights1[41396] <= 16'b0000000000001010;
        weights1[41397] <= 16'b0000000000001001;
        weights1[41398] <= 16'b0000000000000010;
        weights1[41399] <= 16'b0000000000000111;
        weights1[41400] <= 16'b0000000000000101;
        weights1[41401] <= 16'b0000000000000000;
        weights1[41402] <= 16'b0000000000001000;
        weights1[41403] <= 16'b0000000000000101;
        weights1[41404] <= 16'b1111111111110111;
        weights1[41405] <= 16'b0000000000000011;
        weights1[41406] <= 16'b0000000000010000;
        weights1[41407] <= 16'b0000000000001011;
        weights1[41408] <= 16'b0000000000001011;
        weights1[41409] <= 16'b0000000000010101;
        weights1[41410] <= 16'b0000000000000100;
        weights1[41411] <= 16'b0000000000001001;
        weights1[41412] <= 16'b0000000000000101;
        weights1[41413] <= 16'b0000000000000101;
        weights1[41414] <= 16'b0000000000010000;
        weights1[41415] <= 16'b0000000000001000;
        weights1[41416] <= 16'b0000000000001001;
        weights1[41417] <= 16'b0000000000010100;
        weights1[41418] <= 16'b0000000000000101;
        weights1[41419] <= 16'b0000000000000111;
        weights1[41420] <= 16'b0000000000011000;
        weights1[41421] <= 16'b0000000000010011;
        weights1[41422] <= 16'b0000000000011011;
        weights1[41423] <= 16'b0000000000011100;
        weights1[41424] <= 16'b0000000000001010;
        weights1[41425] <= 16'b0000000000010111;
        weights1[41426] <= 16'b0000000000010011;
        weights1[41427] <= 16'b0000000000010011;
        weights1[41428] <= 16'b0000000000010001;
        weights1[41429] <= 16'b0000000000010001;
        weights1[41430] <= 16'b0000000000011101;
        weights1[41431] <= 16'b0000000000001111;
        weights1[41432] <= 16'b1111111111111011;
        weights1[41433] <= 16'b0000000000000011;
        weights1[41434] <= 16'b1111111111110010;
        weights1[41435] <= 16'b0000000000000001;
        weights1[41436] <= 16'b0000000000000000;
        weights1[41437] <= 16'b1111111111111100;
        weights1[41438] <= 16'b1111111111111110;
        weights1[41439] <= 16'b1111111111111110;
        weights1[41440] <= 16'b0000000000001010;
        weights1[41441] <= 16'b0000000000001010;
        weights1[41442] <= 16'b0000000000001011;
        weights1[41443] <= 16'b0000000000001110;
        weights1[41444] <= 16'b0000000000010101;
        weights1[41445] <= 16'b0000000000001111;
        weights1[41446] <= 16'b0000000000101100;
        weights1[41447] <= 16'b0000000000010110;
        weights1[41448] <= 16'b0000000000101101;
        weights1[41449] <= 16'b0000000000011011;
        weights1[41450] <= 16'b0000000000100111;
        weights1[41451] <= 16'b0000000000011110;
        weights1[41452] <= 16'b0000000000100111;
        weights1[41453] <= 16'b0000000000011111;
        weights1[41454] <= 16'b0000000000010001;
        weights1[41455] <= 16'b0000000000001111;
        weights1[41456] <= 16'b0000000000001100;
        weights1[41457] <= 16'b0000000000001010;
        weights1[41458] <= 16'b0000000000001000;
        weights1[41459] <= 16'b0000000000000011;
        weights1[41460] <= 16'b1111111111111010;
        weights1[41461] <= 16'b1111111111111010;
        weights1[41462] <= 16'b1111111111101101;
        weights1[41463] <= 16'b1111111111011010;
        weights1[41464] <= 16'b1111111111110111;
        weights1[41465] <= 16'b1111111111111010;
        weights1[41466] <= 16'b1111111111111011;
        weights1[41467] <= 16'b1111111111111101;
        weights1[41468] <= 16'b0000000000001001;
        weights1[41469] <= 16'b0000000000010000;
        weights1[41470] <= 16'b0000000000001010;
        weights1[41471] <= 16'b0000000000000101;
        weights1[41472] <= 16'b0000000000010100;
        weights1[41473] <= 16'b0000000000010110;
        weights1[41474] <= 16'b0000000000100110;
        weights1[41475] <= 16'b0000000000000110;
        weights1[41476] <= 16'b0000000000010101;
        weights1[41477] <= 16'b0000000000001110;
        weights1[41478] <= 16'b0000000000011010;
        weights1[41479] <= 16'b0000000000001011;
        weights1[41480] <= 16'b0000000000000111;
        weights1[41481] <= 16'b0000000000010010;
        weights1[41482] <= 16'b0000000000011100;
        weights1[41483] <= 16'b0000000000000000;
        weights1[41484] <= 16'b0000000000010101;
        weights1[41485] <= 16'b1111111111111100;
        weights1[41486] <= 16'b0000000000000100;
        weights1[41487] <= 16'b0000000000010110;
        weights1[41488] <= 16'b1111111111111001;
        weights1[41489] <= 16'b0000000000001101;
        weights1[41490] <= 16'b1111111111111010;
        weights1[41491] <= 16'b1111111111111100;
        weights1[41492] <= 16'b1111111111111101;
        weights1[41493] <= 16'b1111111111101000;
        weights1[41494] <= 16'b1111111111110110;
        weights1[41495] <= 16'b1111111111111100;
        weights1[41496] <= 16'b0000000000001001;
        weights1[41497] <= 16'b0000000000001110;
        weights1[41498] <= 16'b0000000000001001;
        weights1[41499] <= 16'b0000000000001010;
        weights1[41500] <= 16'b0000000000010100;
        weights1[41501] <= 16'b0000000000010010;
        weights1[41502] <= 16'b0000000000011111;
        weights1[41503] <= 16'b0000000000000110;
        weights1[41504] <= 16'b0000000000000110;
        weights1[41505] <= 16'b0000000000001011;
        weights1[41506] <= 16'b1111111111110100;
        weights1[41507] <= 16'b0000000000001000;
        weights1[41508] <= 16'b0000000000001000;
        weights1[41509] <= 16'b1111111111111011;
        weights1[41510] <= 16'b1111111111111010;
        weights1[41511] <= 16'b0000000000001010;
        weights1[41512] <= 16'b0000000000000000;
        weights1[41513] <= 16'b1111111111111101;
        weights1[41514] <= 16'b0000000000001001;
        weights1[41515] <= 16'b0000000000011010;
        weights1[41516] <= 16'b1111111111111010;
        weights1[41517] <= 16'b0000000000000100;
        weights1[41518] <= 16'b0000000000001010;
        weights1[41519] <= 16'b0000000000001101;
        weights1[41520] <= 16'b1111111111111011;
        weights1[41521] <= 16'b1111111111110001;
        weights1[41522] <= 16'b1111111111110111;
        weights1[41523] <= 16'b1111111111111101;
        weights1[41524] <= 16'b0000000000000010;
        weights1[41525] <= 16'b0000000000001100;
        weights1[41526] <= 16'b1111111111111111;
        weights1[41527] <= 16'b1111111111111100;
        weights1[41528] <= 16'b0000000000000010;
        weights1[41529] <= 16'b0000000000010101;
        weights1[41530] <= 16'b0000000000011010;
        weights1[41531] <= 16'b1111111111111111;
        weights1[41532] <= 16'b0000000000010000;
        weights1[41533] <= 16'b0000000000000000;
        weights1[41534] <= 16'b0000000000001110;
        weights1[41535] <= 16'b0000000000001100;
        weights1[41536] <= 16'b1111111111111110;
        weights1[41537] <= 16'b0000000000001010;
        weights1[41538] <= 16'b0000000000001101;
        weights1[41539] <= 16'b0000000000000010;
        weights1[41540] <= 16'b0000000000001111;
        weights1[41541] <= 16'b0000000000010001;
        weights1[41542] <= 16'b1111111111111000;
        weights1[41543] <= 16'b1111111111111001;
        weights1[41544] <= 16'b0000000000000101;
        weights1[41545] <= 16'b0000000000000110;
        weights1[41546] <= 16'b0000000000000101;
        weights1[41547] <= 16'b1111111111111111;
        weights1[41548] <= 16'b1111111111111101;
        weights1[41549] <= 16'b1111111111111010;
        weights1[41550] <= 16'b1111111111111101;
        weights1[41551] <= 16'b0000000000000000;
        weights1[41552] <= 16'b0000000000000001;
        weights1[41553] <= 16'b0000000000000001;
        weights1[41554] <= 16'b1111111111111100;
        weights1[41555] <= 16'b1111111111110100;
        weights1[41556] <= 16'b1111111111110011;
        weights1[41557] <= 16'b1111111111101001;
        weights1[41558] <= 16'b1111111111100101;
        weights1[41559] <= 16'b1111111111011010;
        weights1[41560] <= 16'b1111111111010000;
        weights1[41561] <= 16'b1111111111010001;
        weights1[41562] <= 16'b1111111111010000;
        weights1[41563] <= 16'b1111111111010110;
        weights1[41564] <= 16'b1111111111001110;
        weights1[41565] <= 16'b1111111111010000;
        weights1[41566] <= 16'b1111111111100010;
        weights1[41567] <= 16'b1111111111010111;
        weights1[41568] <= 16'b1111111111010100;
        weights1[41569] <= 16'b1111111111011110;
        weights1[41570] <= 16'b1111111111101100;
        weights1[41571] <= 16'b1111111111100010;
        weights1[41572] <= 16'b1111111111101000;
        weights1[41573] <= 16'b1111111111110011;
        weights1[41574] <= 16'b1111111111111001;
        weights1[41575] <= 16'b1111111111111000;
        weights1[41576] <= 16'b1111111111111011;
        weights1[41577] <= 16'b1111111111111011;
        weights1[41578] <= 16'b1111111111111101;
        weights1[41579] <= 16'b1111111111111101;
        weights1[41580] <= 16'b0000000000000000;
        weights1[41581] <= 16'b1111111111111111;
        weights1[41582] <= 16'b1111111111111010;
        weights1[41583] <= 16'b1111111111110000;
        weights1[41584] <= 16'b1111111111100110;
        weights1[41585] <= 16'b1111111111011111;
        weights1[41586] <= 16'b1111111111010110;
        weights1[41587] <= 16'b1111111111001101;
        weights1[41588] <= 16'b1111111111001010;
        weights1[41589] <= 16'b1111111111000011;
        weights1[41590] <= 16'b1111111110111111;
        weights1[41591] <= 16'b1111111110111101;
        weights1[41592] <= 16'b1111111110111101;
        weights1[41593] <= 16'b1111111110111101;
        weights1[41594] <= 16'b1111111111001110;
        weights1[41595] <= 16'b1111111111010011;
        weights1[41596] <= 16'b1111111111010011;
        weights1[41597] <= 16'b1111111111001111;
        weights1[41598] <= 16'b1111111111100001;
        weights1[41599] <= 16'b1111111111100100;
        weights1[41600] <= 16'b1111111111100101;
        weights1[41601] <= 16'b1111111111101010;
        weights1[41602] <= 16'b1111111111101001;
        weights1[41603] <= 16'b1111111111100111;
        weights1[41604] <= 16'b1111111111101111;
        weights1[41605] <= 16'b1111111111111100;
        weights1[41606] <= 16'b1111111111111111;
        weights1[41607] <= 16'b1111111111111011;
        weights1[41608] <= 16'b1111111111111100;
        weights1[41609] <= 16'b1111111111111110;
        weights1[41610] <= 16'b1111111111111000;
        weights1[41611] <= 16'b1111111111101010;
        weights1[41612] <= 16'b1111111111010101;
        weights1[41613] <= 16'b1111111111010010;
        weights1[41614] <= 16'b1111111110111110;
        weights1[41615] <= 16'b1111111110111000;
        weights1[41616] <= 16'b1111111111000011;
        weights1[41617] <= 16'b1111111110110100;
        weights1[41618] <= 16'b1111111110101101;
        weights1[41619] <= 16'b1111111110110110;
        weights1[41620] <= 16'b1111111110111101;
        weights1[41621] <= 16'b1111111111001001;
        weights1[41622] <= 16'b1111111111001100;
        weights1[41623] <= 16'b1111111111001011;
        weights1[41624] <= 16'b1111111110111101;
        weights1[41625] <= 16'b1111111110111100;
        weights1[41626] <= 16'b1111111111010111;
        weights1[41627] <= 16'b1111111111011011;
        weights1[41628] <= 16'b1111111111011101;
        weights1[41629] <= 16'b1111111111100000;
        weights1[41630] <= 16'b1111111111100001;
        weights1[41631] <= 16'b1111111111101000;
        weights1[41632] <= 16'b1111111111011101;
        weights1[41633] <= 16'b1111111111101110;
        weights1[41634] <= 16'b1111111111110010;
        weights1[41635] <= 16'b1111111111111000;
        weights1[41636] <= 16'b1111111111111100;
        weights1[41637] <= 16'b1111111111111010;
        weights1[41638] <= 16'b1111111111110010;
        weights1[41639] <= 16'b1111111111100011;
        weights1[41640] <= 16'b1111111111010100;
        weights1[41641] <= 16'b1111111111001000;
        weights1[41642] <= 16'b1111111111000010;
        weights1[41643] <= 16'b1111111110110110;
        weights1[41644] <= 16'b1111111110111010;
        weights1[41645] <= 16'b1111111110111010;
        weights1[41646] <= 16'b1111111111000100;
        weights1[41647] <= 16'b1111111111001101;
        weights1[41648] <= 16'b1111111111010000;
        weights1[41649] <= 16'b1111111110110111;
        weights1[41650] <= 16'b1111111111011000;
        weights1[41651] <= 16'b1111111111001011;
        weights1[41652] <= 16'b1111111111001001;
        weights1[41653] <= 16'b1111111111011100;
        weights1[41654] <= 16'b1111111111010100;
        weights1[41655] <= 16'b1111111110111111;
        weights1[41656] <= 16'b1111111111001111;
        weights1[41657] <= 16'b1111111111010000;
        weights1[41658] <= 16'b1111111111001101;
        weights1[41659] <= 16'b1111111111011010;
        weights1[41660] <= 16'b1111111111011101;
        weights1[41661] <= 16'b1111111111100111;
        weights1[41662] <= 16'b1111111111110000;
        weights1[41663] <= 16'b1111111111110100;
        weights1[41664] <= 16'b1111111111111110;
        weights1[41665] <= 16'b1111111111110111;
        weights1[41666] <= 16'b1111111111110011;
        weights1[41667] <= 16'b1111111111101001;
        weights1[41668] <= 16'b1111111111010101;
        weights1[41669] <= 16'b1111111111000101;
        weights1[41670] <= 16'b1111111111011011;
        weights1[41671] <= 16'b1111111111000111;
        weights1[41672] <= 16'b1111111111010111;
        weights1[41673] <= 16'b1111111111001011;
        weights1[41674] <= 16'b1111111110111010;
        weights1[41675] <= 16'b1111111111010001;
        weights1[41676] <= 16'b1111111111010111;
        weights1[41677] <= 16'b1111111111011000;
        weights1[41678] <= 16'b1111111111001101;
        weights1[41679] <= 16'b1111111111100101;
        weights1[41680] <= 16'b1111111111111001;
        weights1[41681] <= 16'b1111111111011001;
        weights1[41682] <= 16'b1111111111010011;
        weights1[41683] <= 16'b1111111111010000;
        weights1[41684] <= 16'b1111111111010100;
        weights1[41685] <= 16'b1111111111100111;
        weights1[41686] <= 16'b1111111111100000;
        weights1[41687] <= 16'b1111111111011110;
        weights1[41688] <= 16'b1111111111101110;
        weights1[41689] <= 16'b1111111111101000;
        weights1[41690] <= 16'b1111111111111011;
        weights1[41691] <= 16'b1111111111111110;
        weights1[41692] <= 16'b1111111111111111;
        weights1[41693] <= 16'b1111111111111001;
        weights1[41694] <= 16'b1111111111110110;
        weights1[41695] <= 16'b1111111111100101;
        weights1[41696] <= 16'b1111111111011011;
        weights1[41697] <= 16'b1111111111010100;
        weights1[41698] <= 16'b1111111111011111;
        weights1[41699] <= 16'b1111111111010001;
        weights1[41700] <= 16'b1111111111111101;
        weights1[41701] <= 16'b1111111111111100;
        weights1[41702] <= 16'b1111111111100001;
        weights1[41703] <= 16'b1111111111111100;
        weights1[41704] <= 16'b0000000000000001;
        weights1[41705] <= 16'b1111111111001100;
        weights1[41706] <= 16'b1111111111010101;
        weights1[41707] <= 16'b1111111111001110;
        weights1[41708] <= 16'b1111111111010101;
        weights1[41709] <= 16'b1111111111100010;
        weights1[41710] <= 16'b1111111111001000;
        weights1[41711] <= 16'b1111111111000110;
        weights1[41712] <= 16'b1111111111000101;
        weights1[41713] <= 16'b1111111111001010;
        weights1[41714] <= 16'b1111111111101000;
        weights1[41715] <= 16'b1111111111110101;
        weights1[41716] <= 16'b1111111111111001;
        weights1[41717] <= 16'b1111111111101110;
        weights1[41718] <= 16'b1111111111111001;
        weights1[41719] <= 16'b0000000000000001;
        weights1[41720] <= 16'b0000000000000000;
        weights1[41721] <= 16'b0000000000000001;
        weights1[41722] <= 16'b1111111111111010;
        weights1[41723] <= 16'b1111111111110011;
        weights1[41724] <= 16'b1111111111101000;
        weights1[41725] <= 16'b1111111111100001;
        weights1[41726] <= 16'b1111111111100111;
        weights1[41727] <= 16'b1111111111111101;
        weights1[41728] <= 16'b0000000000000010;
        weights1[41729] <= 16'b0000000000000001;
        weights1[41730] <= 16'b1111111111111101;
        weights1[41731] <= 16'b1111111111011110;
        weights1[41732] <= 16'b1111111111111101;
        weights1[41733] <= 16'b1111111111110011;
        weights1[41734] <= 16'b0000000000001111;
        weights1[41735] <= 16'b1111111111111000;
        weights1[41736] <= 16'b1111111111100010;
        weights1[41737] <= 16'b0000000000010101;
        weights1[41738] <= 16'b1111111111101101;
        weights1[41739] <= 16'b1111111111110011;
        weights1[41740] <= 16'b1111111111100101;
        weights1[41741] <= 16'b0000000000000100;
        weights1[41742] <= 16'b0000000000000001;
        weights1[41743] <= 16'b0000000000000010;
        weights1[41744] <= 16'b1111111111111101;
        weights1[41745] <= 16'b0000000000001011;
        weights1[41746] <= 16'b1111111111101100;
        weights1[41747] <= 16'b1111111111111111;
        weights1[41748] <= 16'b0000000000000010;
        weights1[41749] <= 16'b0000000000000000;
        weights1[41750] <= 16'b1111111111111101;
        weights1[41751] <= 16'b1111111111110011;
        weights1[41752] <= 16'b1111111111100100;
        weights1[41753] <= 16'b1111111111110000;
        weights1[41754] <= 16'b1111111111100000;
        weights1[41755] <= 16'b0000000000001000;
        weights1[41756] <= 16'b1111111111110101;
        weights1[41757] <= 16'b0000000000000111;
        weights1[41758] <= 16'b0000000000011010;
        weights1[41759] <= 16'b0000000000010111;
        weights1[41760] <= 16'b0000000000001101;
        weights1[41761] <= 16'b0000000000011001;
        weights1[41762] <= 16'b0000000000000101;
        weights1[41763] <= 16'b0000000000000010;
        weights1[41764] <= 16'b0000000000100100;
        weights1[41765] <= 16'b0000000000010010;
        weights1[41766] <= 16'b0000000000010110;
        weights1[41767] <= 16'b0000000000100001;
        weights1[41768] <= 16'b0000000000001000;
        weights1[41769] <= 16'b0000000000010000;
        weights1[41770] <= 16'b0000000000010001;
        weights1[41771] <= 16'b1111111111110101;
        weights1[41772] <= 16'b0000000000000101;
        weights1[41773] <= 16'b1111111111110100;
        weights1[41774] <= 16'b1111111111101111;
        weights1[41775] <= 16'b1111111111111110;
        weights1[41776] <= 16'b0000000000000000;
        weights1[41777] <= 16'b0000000000000100;
        weights1[41778] <= 16'b0000000000000101;
        weights1[41779] <= 16'b1111111111111101;
        weights1[41780] <= 16'b1111111111101111;
        weights1[41781] <= 16'b0000000000000011;
        weights1[41782] <= 16'b0000000000000000;
        weights1[41783] <= 16'b1111111111110001;
        weights1[41784] <= 16'b0000000000001010;
        weights1[41785] <= 16'b0000000000000000;
        weights1[41786] <= 16'b1111111111100111;
        weights1[41787] <= 16'b0000000000000101;
        weights1[41788] <= 16'b0000000000010110;
        weights1[41789] <= 16'b0000000000001100;
        weights1[41790] <= 16'b0000000000000010;
        weights1[41791] <= 16'b0000000000001100;
        weights1[41792] <= 16'b0000000000000101;
        weights1[41793] <= 16'b0000000000010011;
        weights1[41794] <= 16'b1111111111110101;
        weights1[41795] <= 16'b0000000000001001;
        weights1[41796] <= 16'b1111111111100011;
        weights1[41797] <= 16'b0000000000001110;
        weights1[41798] <= 16'b1111111111111001;
        weights1[41799] <= 16'b1111111111110010;
        weights1[41800] <= 16'b1111111111111000;
        weights1[41801] <= 16'b0000000000000100;
        weights1[41802] <= 16'b1111111111101100;
        weights1[41803] <= 16'b1111111111111011;
        weights1[41804] <= 16'b0000000000000010;
        weights1[41805] <= 16'b0000000000000101;
        weights1[41806] <= 16'b0000000000010100;
        weights1[41807] <= 16'b0000000000001110;
        weights1[41808] <= 16'b1111111111110110;
        weights1[41809] <= 16'b1111111111101010;
        weights1[41810] <= 16'b0000000000001000;
        weights1[41811] <= 16'b1111111111101101;
        weights1[41812] <= 16'b1111111111101110;
        weights1[41813] <= 16'b1111111111101100;
        weights1[41814] <= 16'b1111111111101111;
        weights1[41815] <= 16'b1111111111111100;
        weights1[41816] <= 16'b1111111111111110;
        weights1[41817] <= 16'b0000000000001010;
        weights1[41818] <= 16'b0000000000001011;
        weights1[41819] <= 16'b0000000000001011;
        weights1[41820] <= 16'b0000000000000110;
        weights1[41821] <= 16'b0000000000011000;
        weights1[41822] <= 16'b0000000000001100;
        weights1[41823] <= 16'b0000000000001000;
        weights1[41824] <= 16'b1111111111101100;
        weights1[41825] <= 16'b1111111111111011;
        weights1[41826] <= 16'b1111111111111000;
        weights1[41827] <= 16'b1111111111110001;
        weights1[41828] <= 16'b1111111111111111;
        weights1[41829] <= 16'b0000000000001010;
        weights1[41830] <= 16'b1111111111111001;
        weights1[41831] <= 16'b0000000000000010;
        weights1[41832] <= 16'b0000000000000111;
        weights1[41833] <= 16'b0000000000001000;
        weights1[41834] <= 16'b0000000000001010;
        weights1[41835] <= 16'b0000000000001110;
        weights1[41836] <= 16'b0000000000010011;
        weights1[41837] <= 16'b0000000000001011;
        weights1[41838] <= 16'b0000000000011111;
        weights1[41839] <= 16'b0000000000000110;
        weights1[41840] <= 16'b0000000000001000;
        weights1[41841] <= 16'b0000000000000101;
        weights1[41842] <= 16'b0000000000010011;
        weights1[41843] <= 16'b1111111111101001;
        weights1[41844] <= 16'b1111111111111101;
        weights1[41845] <= 16'b1111111111111101;
        weights1[41846] <= 16'b1111111111110110;
        weights1[41847] <= 16'b1111111111111000;
        weights1[41848] <= 16'b0000000000001101;
        weights1[41849] <= 16'b0000000000000000;
        weights1[41850] <= 16'b1111111111110000;
        weights1[41851] <= 16'b1111111111111010;
        weights1[41852] <= 16'b0000000000001011;
        weights1[41853] <= 16'b0000000000001000;
        weights1[41854] <= 16'b1111111111111110;
        weights1[41855] <= 16'b1111111111101101;
        weights1[41856] <= 16'b1111111111110111;
        weights1[41857] <= 16'b0000000000001111;
        weights1[41858] <= 16'b0000000000000001;
        weights1[41859] <= 16'b0000000000000110;
        weights1[41860] <= 16'b0000000000001111;
        weights1[41861] <= 16'b0000000000010000;
        weights1[41862] <= 16'b0000000000110000;
        weights1[41863] <= 16'b0000000000101100;
        weights1[41864] <= 16'b0000000000011110;
        weights1[41865] <= 16'b0000000000010010;
        weights1[41866] <= 16'b0000000000000101;
        weights1[41867] <= 16'b0000000000000110;
        weights1[41868] <= 16'b0000000000011100;
        weights1[41869] <= 16'b0000000000010011;
        weights1[41870] <= 16'b0000000000001110;
        weights1[41871] <= 16'b0000000000001000;
        weights1[41872] <= 16'b0000000000000101;
        weights1[41873] <= 16'b1111111111101100;
        weights1[41874] <= 16'b1111111111110111;
        weights1[41875] <= 16'b1111111111111001;
        weights1[41876] <= 16'b1111111111111101;
        weights1[41877] <= 16'b1111111111111110;
        weights1[41878] <= 16'b0000000000001001;
        weights1[41879] <= 16'b1111111111110000;
        weights1[41880] <= 16'b0000000000001010;
        weights1[41881] <= 16'b1111111111111100;
        weights1[41882] <= 16'b1111111111101100;
        weights1[41883] <= 16'b1111111111011000;
        weights1[41884] <= 16'b0000000000000110;
        weights1[41885] <= 16'b0000000000000110;
        weights1[41886] <= 16'b0000000000001101;
        weights1[41887] <= 16'b0000000000011100;
        weights1[41888] <= 16'b0000000000001101;
        weights1[41889] <= 16'b0000000000001011;
        weights1[41890] <= 16'b0000000000101111;
        weights1[41891] <= 16'b0000000000100111;
        weights1[41892] <= 16'b0000000000101011;
        weights1[41893] <= 16'b0000000000100001;
        weights1[41894] <= 16'b0000000000100000;
        weights1[41895] <= 16'b0000000000100100;
        weights1[41896] <= 16'b0000000000000011;
        weights1[41897] <= 16'b0000000000100111;
        weights1[41898] <= 16'b0000000000001100;
        weights1[41899] <= 16'b0000000000001011;
        weights1[41900] <= 16'b1111111111111101;
        weights1[41901] <= 16'b0000000000001001;
        weights1[41902] <= 16'b1111111111111111;
        weights1[41903] <= 16'b1111111111110011;
        weights1[41904] <= 16'b0000000000000010;
        weights1[41905] <= 16'b0000000000001001;
        weights1[41906] <= 16'b1111111111111100;
        weights1[41907] <= 16'b1111111111111000;
        weights1[41908] <= 16'b1111111111101011;
        weights1[41909] <= 16'b1111111111111111;
        weights1[41910] <= 16'b1111111111110000;
        weights1[41911] <= 16'b1111111111110011;
        weights1[41912] <= 16'b1111111111101111;
        weights1[41913] <= 16'b1111111111111011;
        weights1[41914] <= 16'b0000000000010010;
        weights1[41915] <= 16'b0000000000001000;
        weights1[41916] <= 16'b0000000000001110;
        weights1[41917] <= 16'b0000000000011100;
        weights1[41918] <= 16'b0000000000101100;
        weights1[41919] <= 16'b0000000000100001;
        weights1[41920] <= 16'b0000000000100111;
        weights1[41921] <= 16'b0000000001000001;
        weights1[41922] <= 16'b0000000000010100;
        weights1[41923] <= 16'b0000000000011111;
        weights1[41924] <= 16'b0000000000001001;
        weights1[41925] <= 16'b0000000000011000;
        weights1[41926] <= 16'b0000000000100101;
        weights1[41927] <= 16'b0000000000010101;
        weights1[41928] <= 16'b0000000000000111;
        weights1[41929] <= 16'b0000000000010010;
        weights1[41930] <= 16'b1111111111110011;
        weights1[41931] <= 16'b0000000000011000;
        weights1[41932] <= 16'b0000000000001010;
        weights1[41933] <= 16'b0000000000010011;
        weights1[41934] <= 16'b0000000000001101;
        weights1[41935] <= 16'b1111111111111111;
        weights1[41936] <= 16'b0000000000101001;
        weights1[41937] <= 16'b1111111111111011;
        weights1[41938] <= 16'b0000000000000100;
        weights1[41939] <= 16'b0000000000000101;
        weights1[41940] <= 16'b1111111111111110;
        weights1[41941] <= 16'b0000000000000110;
        weights1[41942] <= 16'b0000000000000011;
        weights1[41943] <= 16'b0000000000010000;
        weights1[41944] <= 16'b0000000000001001;
        weights1[41945] <= 16'b0000000000011010;
        weights1[41946] <= 16'b0000000000110001;
        weights1[41947] <= 16'b0000000000011111;
        weights1[41948] <= 16'b0000000000011101;
        weights1[41949] <= 16'b0000000000101110;
        weights1[41950] <= 16'b0000000000101100;
        weights1[41951] <= 16'b0000000000111101;
        weights1[41952] <= 16'b0000000000100110;
        weights1[41953] <= 16'b0000000000110111;
        weights1[41954] <= 16'b0000000000000100;
        weights1[41955] <= 16'b0000000000001011;
        weights1[41956] <= 16'b0000000000000110;
        weights1[41957] <= 16'b0000000000010010;
        weights1[41958] <= 16'b0000000000010001;
        weights1[41959] <= 16'b0000000000001001;
        weights1[41960] <= 16'b0000000000001111;
        weights1[41961] <= 16'b0000000000001100;
        weights1[41962] <= 16'b0000000000001110;
        weights1[41963] <= 16'b0000000000011011;
        weights1[41964] <= 16'b0000000000010001;
        weights1[41965] <= 16'b0000000000001111;
        weights1[41966] <= 16'b0000000000011000;
        weights1[41967] <= 16'b0000000000100111;
        weights1[41968] <= 16'b0000000000001100;
        weights1[41969] <= 16'b0000000000011100;
        weights1[41970] <= 16'b0000000000010001;
        weights1[41971] <= 16'b0000000000000000;
        weights1[41972] <= 16'b0000000000001001;
        weights1[41973] <= 16'b0000000000001010;
        weights1[41974] <= 16'b0000000000011001;
        weights1[41975] <= 16'b0000000000011000;
        weights1[41976] <= 16'b0000000000101101;
        weights1[41977] <= 16'b0000000000110011;
        weights1[41978] <= 16'b0000000000011000;
        weights1[41979] <= 16'b0000000000110010;
        weights1[41980] <= 16'b0000000000101011;
        weights1[41981] <= 16'b0000000000011110;
        weights1[41982] <= 16'b0000000000010010;
        weights1[41983] <= 16'b0000000000010100;
        weights1[41984] <= 16'b0000000000001100;
        weights1[41985] <= 16'b0000000000000101;
        weights1[41986] <= 16'b0000000000011000;
        weights1[41987] <= 16'b0000000000100010;
        weights1[41988] <= 16'b0000000000011100;
        weights1[41989] <= 16'b0000000000100011;
        weights1[41990] <= 16'b0000000000011101;
        weights1[41991] <= 16'b0000000000010100;
        weights1[41992] <= 16'b0000000000101010;
        weights1[41993] <= 16'b0000000000101000;
        weights1[41994] <= 16'b0000000000010101;
        weights1[41995] <= 16'b0000000000011100;
        weights1[41996] <= 16'b0000000000001011;
        weights1[41997] <= 16'b1111111111111101;
        weights1[41998] <= 16'b0000000000001001;
        weights1[41999] <= 16'b0000000000001001;
        weights1[42000] <= 16'b1111111111111111;
        weights1[42001] <= 16'b0000000000000011;
        weights1[42002] <= 16'b0000000000000100;
        weights1[42003] <= 16'b0000000000000011;
        weights1[42004] <= 16'b0000000000010011;
        weights1[42005] <= 16'b0000000000011001;
        weights1[42006] <= 16'b0000000000010010;
        weights1[42007] <= 16'b0000000000010110;
        weights1[42008] <= 16'b0000000000100011;
        weights1[42009] <= 16'b0000000000001000;
        weights1[42010] <= 16'b0000000000010001;
        weights1[42011] <= 16'b0000000000001000;
        weights1[42012] <= 16'b0000000000011101;
        weights1[42013] <= 16'b0000000000010100;
        weights1[42014] <= 16'b0000000000001111;
        weights1[42015] <= 16'b0000000000011010;
        weights1[42016] <= 16'b0000000000011001;
        weights1[42017] <= 16'b0000000000100010;
        weights1[42018] <= 16'b0000000000001011;
        weights1[42019] <= 16'b0000000000001111;
        weights1[42020] <= 16'b0000000000010000;
        weights1[42021] <= 16'b0000000000011000;
        weights1[42022] <= 16'b1111111111111011;
        weights1[42023] <= 16'b0000000000001010;
        weights1[42024] <= 16'b0000000000001010;
        weights1[42025] <= 16'b0000000000000000;
        weights1[42026] <= 16'b1111111111111110;
        weights1[42027] <= 16'b0000000000000000;
        weights1[42028] <= 16'b1111111111101111;
        weights1[42029] <= 16'b1111111111101001;
        weights1[42030] <= 16'b1111111111100111;
        weights1[42031] <= 16'b1111111111101111;
        weights1[42032] <= 16'b1111111111110011;
        weights1[42033] <= 16'b1111111111110111;
        weights1[42034] <= 16'b1111111111110110;
        weights1[42035] <= 16'b1111111111110011;
        weights1[42036] <= 16'b1111111111110101;
        weights1[42037] <= 16'b1111111111100111;
        weights1[42038] <= 16'b1111111111110010;
        weights1[42039] <= 16'b0000000000011001;
        weights1[42040] <= 16'b1111111111111111;
        weights1[42041] <= 16'b0000000000001000;
        weights1[42042] <= 16'b0000000000000110;
        weights1[42043] <= 16'b0000000000001000;
        weights1[42044] <= 16'b0000000000000000;
        weights1[42045] <= 16'b0000000000000110;
        weights1[42046] <= 16'b0000000000001011;
        weights1[42047] <= 16'b1111111111110110;
        weights1[42048] <= 16'b0000000000000011;
        weights1[42049] <= 16'b0000000000000110;
        weights1[42050] <= 16'b1111111111101011;
        weights1[42051] <= 16'b1111111111111000;
        weights1[42052] <= 16'b1111111111101101;
        weights1[42053] <= 16'b1111111111111000;
        weights1[42054] <= 16'b1111111111111011;
        weights1[42055] <= 16'b1111111111111110;
        weights1[42056] <= 16'b1111111111100001;
        weights1[42057] <= 16'b1111111111010100;
        weights1[42058] <= 16'b1111111111001110;
        weights1[42059] <= 16'b1111111111000100;
        weights1[42060] <= 16'b1111111111011110;
        weights1[42061] <= 16'b1111111111010101;
        weights1[42062] <= 16'b1111111111010011;
        weights1[42063] <= 16'b1111111111001010;
        weights1[42064] <= 16'b1111111111000111;
        weights1[42065] <= 16'b1111111110111101;
        weights1[42066] <= 16'b1111111111010000;
        weights1[42067] <= 16'b1111111111011000;
        weights1[42068] <= 16'b1111111111011011;
        weights1[42069] <= 16'b1111111111100100;
        weights1[42070] <= 16'b1111111111101111;
        weights1[42071] <= 16'b1111111111111011;
        weights1[42072] <= 16'b1111111111110100;
        weights1[42073] <= 16'b1111111111110011;
        weights1[42074] <= 16'b1111111111110011;
        weights1[42075] <= 16'b1111111111100111;
        weights1[42076] <= 16'b1111111111110101;
        weights1[42077] <= 16'b1111111111101100;
        weights1[42078] <= 16'b1111111111001111;
        weights1[42079] <= 16'b1111111111011111;
        weights1[42080] <= 16'b1111111111011011;
        weights1[42081] <= 16'b1111111111101111;
        weights1[42082] <= 16'b1111111111110000;
        weights1[42083] <= 16'b1111111111111110;
        weights1[42084] <= 16'b1111111111011100;
        weights1[42085] <= 16'b1111111111010000;
        weights1[42086] <= 16'b1111111111000001;
        weights1[42087] <= 16'b1111111110101010;
        weights1[42088] <= 16'b1111111110110000;
        weights1[42089] <= 16'b1111111110001110;
        weights1[42090] <= 16'b1111111101110000;
        weights1[42091] <= 16'b1111111101111000;
        weights1[42092] <= 16'b1111111101111000;
        weights1[42093] <= 16'b1111111110101110;
        weights1[42094] <= 16'b1111111111000110;
        weights1[42095] <= 16'b1111111111001100;
        weights1[42096] <= 16'b1111111111001111;
        weights1[42097] <= 16'b1111111111100111;
        weights1[42098] <= 16'b1111111111111010;
        weights1[42099] <= 16'b1111111111100110;
        weights1[42100] <= 16'b1111111111101010;
        weights1[42101] <= 16'b1111111111111110;
        weights1[42102] <= 16'b1111111111100000;
        weights1[42103] <= 16'b1111111111110011;
        weights1[42104] <= 16'b1111111111100010;
        weights1[42105] <= 16'b1111111111011100;
        weights1[42106] <= 16'b1111111111010010;
        weights1[42107] <= 16'b1111111111010110;
        weights1[42108] <= 16'b1111111111011111;
        weights1[42109] <= 16'b1111111111111100;
        weights1[42110] <= 16'b1111111111110111;
        weights1[42111] <= 16'b1111111111111110;
        weights1[42112] <= 16'b1111111111011001;
        weights1[42113] <= 16'b1111111111010010;
        weights1[42114] <= 16'b1111111111000101;
        weights1[42115] <= 16'b1111111110110000;
        weights1[42116] <= 16'b1111111110011011;
        weights1[42117] <= 16'b1111111110010011;
        weights1[42118] <= 16'b1111111110010011;
        weights1[42119] <= 16'b1111111110100111;
        weights1[42120] <= 16'b1111111111010000;
        weights1[42121] <= 16'b1111111111111000;
        weights1[42122] <= 16'b1111111111111100;
        weights1[42123] <= 16'b0000000000000000;
        weights1[42124] <= 16'b0000000000000011;
        weights1[42125] <= 16'b0000000000000101;
        weights1[42126] <= 16'b0000000000001100;
        weights1[42127] <= 16'b0000000000010011;
        weights1[42128] <= 16'b1111111111100111;
        weights1[42129] <= 16'b1111111111111010;
        weights1[42130] <= 16'b0000000000000101;
        weights1[42131] <= 16'b1111111111011001;
        weights1[42132] <= 16'b1111111111010010;
        weights1[42133] <= 16'b1111111111100011;
        weights1[42134] <= 16'b1111111111101001;
        weights1[42135] <= 16'b1111111111100010;
        weights1[42136] <= 16'b0000000000000001;
        weights1[42137] <= 16'b1111111111111011;
        weights1[42138] <= 16'b1111111111110111;
        weights1[42139] <= 16'b1111111111111011;
        weights1[42140] <= 16'b1111111111100011;
        weights1[42141] <= 16'b1111111111011000;
        weights1[42142] <= 16'b1111111111001110;
        weights1[42143] <= 16'b1111111110110111;
        weights1[42144] <= 16'b1111111110101101;
        weights1[42145] <= 16'b1111111110101100;
        weights1[42146] <= 16'b1111111111000101;
        weights1[42147] <= 16'b0000000000000100;
        weights1[42148] <= 16'b0000000000010100;
        weights1[42149] <= 16'b0000000000100011;
        weights1[42150] <= 16'b0000000000011000;
        weights1[42151] <= 16'b0000000000001101;
        weights1[42152] <= 16'b0000000000001000;
        weights1[42153] <= 16'b1111111111101010;
        weights1[42154] <= 16'b1111111111101110;
        weights1[42155] <= 16'b1111111111110111;
        weights1[42156] <= 16'b1111111111011101;
        weights1[42157] <= 16'b1111111111100100;
        weights1[42158] <= 16'b1111111111110100;
        weights1[42159] <= 16'b1111111111011111;
        weights1[42160] <= 16'b1111111111101010;
        weights1[42161] <= 16'b1111111111111111;
        weights1[42162] <= 16'b1111111111100000;
        weights1[42163] <= 16'b1111111111011111;
        weights1[42164] <= 16'b1111111111111000;
        weights1[42165] <= 16'b1111111111111000;
        weights1[42166] <= 16'b1111111111110100;
        weights1[42167] <= 16'b1111111111111110;
        weights1[42168] <= 16'b1111111111100001;
        weights1[42169] <= 16'b1111111111010000;
        weights1[42170] <= 16'b1111111111001010;
        weights1[42171] <= 16'b1111111111000100;
        weights1[42172] <= 16'b1111111111001110;
        weights1[42173] <= 16'b1111111111101000;
        weights1[42174] <= 16'b0000000000000000;
        weights1[42175] <= 16'b0000000000100110;
        weights1[42176] <= 16'b0000000000110100;
        weights1[42177] <= 16'b0000000000000111;
        weights1[42178] <= 16'b0000000000011000;
        weights1[42179] <= 16'b1111111111111001;
        weights1[42180] <= 16'b1111111111110110;
        weights1[42181] <= 16'b1111111111110011;
        weights1[42182] <= 16'b1111111111111010;
        weights1[42183] <= 16'b1111111111110101;
        weights1[42184] <= 16'b1111111111111010;
        weights1[42185] <= 16'b1111111111111101;
        weights1[42186] <= 16'b1111111111110111;
        weights1[42187] <= 16'b1111111111101100;
        weights1[42188] <= 16'b1111111111110001;
        weights1[42189] <= 16'b1111111111111101;
        weights1[42190] <= 16'b1111111111101101;
        weights1[42191] <= 16'b1111111111100110;
        weights1[42192] <= 16'b1111111111111001;
        weights1[42193] <= 16'b1111111111101101;
        weights1[42194] <= 16'b0000000000000000;
        weights1[42195] <= 16'b0000000000000000;
        weights1[42196] <= 16'b1111111111011111;
        weights1[42197] <= 16'b1111111111011111;
        weights1[42198] <= 16'b1111111111010101;
        weights1[42199] <= 16'b1111111111001110;
        weights1[42200] <= 16'b1111111111011010;
        weights1[42201] <= 16'b1111111111111010;
        weights1[42202] <= 16'b0000000000100000;
        weights1[42203] <= 16'b0000000000011011;
        weights1[42204] <= 16'b0000000000000100;
        weights1[42205] <= 16'b1111111111110111;
        weights1[42206] <= 16'b1111111111110101;
        weights1[42207] <= 16'b0000000000000111;
        weights1[42208] <= 16'b1111111111111000;
        weights1[42209] <= 16'b0000000000001100;
        weights1[42210] <= 16'b1111111111111000;
        weights1[42211] <= 16'b1111111111011001;
        weights1[42212] <= 16'b1111111111101111;
        weights1[42213] <= 16'b0000000000010111;
        weights1[42214] <= 16'b1111111111111001;
        weights1[42215] <= 16'b1111111111100101;
        weights1[42216] <= 16'b1111111111011100;
        weights1[42217] <= 16'b1111111111101010;
        weights1[42218] <= 16'b1111111111011100;
        weights1[42219] <= 16'b1111111111011111;
        weights1[42220] <= 16'b1111111111110011;
        weights1[42221] <= 16'b1111111111111111;
        weights1[42222] <= 16'b0000000000000000;
        weights1[42223] <= 16'b1111111111111111;
        weights1[42224] <= 16'b1111111111101110;
        weights1[42225] <= 16'b1111111111101000;
        weights1[42226] <= 16'b1111111111100000;
        weights1[42227] <= 16'b1111111111110110;
        weights1[42228] <= 16'b1111111111111011;
        weights1[42229] <= 16'b0000000000010011;
        weights1[42230] <= 16'b0000000000100000;
        weights1[42231] <= 16'b0000000000100100;
        weights1[42232] <= 16'b0000000000001101;
        weights1[42233] <= 16'b0000000000001100;
        weights1[42234] <= 16'b1111111111110101;
        weights1[42235] <= 16'b1111111111110101;
        weights1[42236] <= 16'b1111111111110101;
        weights1[42237] <= 16'b0000000000000100;
        weights1[42238] <= 16'b1111111111111100;
        weights1[42239] <= 16'b1111111111010101;
        weights1[42240] <= 16'b1111111111111000;
        weights1[42241] <= 16'b1111111111110100;
        weights1[42242] <= 16'b1111111111111010;
        weights1[42243] <= 16'b1111111111010101;
        weights1[42244] <= 16'b1111111111111011;
        weights1[42245] <= 16'b1111111111110111;
        weights1[42246] <= 16'b1111111111110111;
        weights1[42247] <= 16'b1111111111111100;
        weights1[42248] <= 16'b1111111111110011;
        weights1[42249] <= 16'b1111111111110101;
        weights1[42250] <= 16'b1111111111111011;
        weights1[42251] <= 16'b1111111111111110;
        weights1[42252] <= 16'b1111111111111001;
        weights1[42253] <= 16'b1111111111110010;
        weights1[42254] <= 16'b1111111111110101;
        weights1[42255] <= 16'b1111111111111010;
        weights1[42256] <= 16'b0000000000011101;
        weights1[42257] <= 16'b0000000000010111;
        weights1[42258] <= 16'b0000000000010111;
        weights1[42259] <= 16'b0000000000000011;
        weights1[42260] <= 16'b0000000000001100;
        weights1[42261] <= 16'b1111111111110010;
        weights1[42262] <= 16'b1111111111110101;
        weights1[42263] <= 16'b1111111111110111;
        weights1[42264] <= 16'b1111111111011111;
        weights1[42265] <= 16'b0000000000001001;
        weights1[42266] <= 16'b1111111111111100;
        weights1[42267] <= 16'b0000000000000101;
        weights1[42268] <= 16'b0000000000011001;
        weights1[42269] <= 16'b0000000000000100;
        weights1[42270] <= 16'b0000000000000100;
        weights1[42271] <= 16'b1111111111110110;
        weights1[42272] <= 16'b1111111111101110;
        weights1[42273] <= 16'b1111111111111000;
        weights1[42274] <= 16'b0000000000000001;
        weights1[42275] <= 16'b0000000000000100;
        weights1[42276] <= 16'b1111111111111101;
        weights1[42277] <= 16'b1111111111111101;
        weights1[42278] <= 16'b1111111111111111;
        weights1[42279] <= 16'b1111111111111101;
        weights1[42280] <= 16'b1111111111111100;
        weights1[42281] <= 16'b1111111111111010;
        weights1[42282] <= 16'b1111111111111111;
        weights1[42283] <= 16'b0000000000000100;
        weights1[42284] <= 16'b0000000000011001;
        weights1[42285] <= 16'b0000000000010010;
        weights1[42286] <= 16'b0000000000010000;
        weights1[42287] <= 16'b1111111111110101;
        weights1[42288] <= 16'b1111111111101111;
        weights1[42289] <= 16'b1111111111111010;
        weights1[42290] <= 16'b1111111111101110;
        weights1[42291] <= 16'b1111111111110011;
        weights1[42292] <= 16'b0000000000000111;
        weights1[42293] <= 16'b0000000000000110;
        weights1[42294] <= 16'b1111111111111100;
        weights1[42295] <= 16'b1111111111101110;
        weights1[42296] <= 16'b0000000000000111;
        weights1[42297] <= 16'b1111111111111110;
        weights1[42298] <= 16'b1111111111110000;
        weights1[42299] <= 16'b1111111111110011;
        weights1[42300] <= 16'b1111111111101110;
        weights1[42301] <= 16'b1111111111110010;
        weights1[42302] <= 16'b1111111111110100;
        weights1[42303] <= 16'b1111111111111011;
        weights1[42304] <= 16'b1111111111111110;
        weights1[42305] <= 16'b0000000000000001;
        weights1[42306] <= 16'b0000000000000000;
        weights1[42307] <= 16'b0000000000000000;
        weights1[42308] <= 16'b1111111111111111;
        weights1[42309] <= 16'b1111111111111111;
        weights1[42310] <= 16'b0000000000000101;
        weights1[42311] <= 16'b0000000000001000;
        weights1[42312] <= 16'b0000000000010000;
        weights1[42313] <= 16'b0000000000000011;
        weights1[42314] <= 16'b1111111111110110;
        weights1[42315] <= 16'b1111111111110010;
        weights1[42316] <= 16'b1111111111101000;
        weights1[42317] <= 16'b1111111111101101;
        weights1[42318] <= 16'b1111111111111000;
        weights1[42319] <= 16'b1111111111110001;
        weights1[42320] <= 16'b1111111111100100;
        weights1[42321] <= 16'b1111111111101110;
        weights1[42322] <= 16'b1111111111110000;
        weights1[42323] <= 16'b1111111111101101;
        weights1[42324] <= 16'b1111111111111001;
        weights1[42325] <= 16'b1111111111111101;
        weights1[42326] <= 16'b1111111111110100;
        weights1[42327] <= 16'b1111111111110111;
        weights1[42328] <= 16'b1111111111111000;
        weights1[42329] <= 16'b1111111111110001;
        weights1[42330] <= 16'b1111111111111000;
        weights1[42331] <= 16'b1111111111110111;
        weights1[42332] <= 16'b1111111111111011;
        weights1[42333] <= 16'b1111111111111101;
        weights1[42334] <= 16'b1111111111111111;
        weights1[42335] <= 16'b0000000000000001;
        weights1[42336] <= 16'b0000000000000000;
        weights1[42337] <= 16'b0000000000000000;
        weights1[42338] <= 16'b0000000000000000;
        weights1[42339] <= 16'b0000000000000000;
        weights1[42340] <= 16'b0000000000000000;
        weights1[42341] <= 16'b0000000000000000;
        weights1[42342] <= 16'b0000000000000000;
        weights1[42343] <= 16'b0000000000000000;
        weights1[42344] <= 16'b0000000000000000;
        weights1[42345] <= 16'b0000000000000000;
        weights1[42346] <= 16'b0000000000000000;
        weights1[42347] <= 16'b0000000000000000;
        weights1[42348] <= 16'b0000000000000000;
        weights1[42349] <= 16'b0000000000000000;
        weights1[42350] <= 16'b0000000000000000;
        weights1[42351] <= 16'b0000000000000000;
        weights1[42352] <= 16'b0000000000000000;
        weights1[42353] <= 16'b0000000000000000;
        weights1[42354] <= 16'b0000000000000000;
        weights1[42355] <= 16'b0000000000000000;
        weights1[42356] <= 16'b0000000000000000;
        weights1[42357] <= 16'b0000000000000000;
        weights1[42358] <= 16'b0000000000000000;
        weights1[42359] <= 16'b0000000000000000;
        weights1[42360] <= 16'b0000000000000000;
        weights1[42361] <= 16'b0000000000000000;
        weights1[42362] <= 16'b0000000000000000;
        weights1[42363] <= 16'b0000000000000000;
        weights1[42364] <= 16'b0000000000000000;
        weights1[42365] <= 16'b0000000000000000;
        weights1[42366] <= 16'b0000000000000000;
        weights1[42367] <= 16'b0000000000000000;
        weights1[42368] <= 16'b0000000000000000;
        weights1[42369] <= 16'b0000000000000000;
        weights1[42370] <= 16'b0000000000000000;
        weights1[42371] <= 16'b0000000000000000;
        weights1[42372] <= 16'b0000000000000000;
        weights1[42373] <= 16'b0000000000000000;
        weights1[42374] <= 16'b0000000000000000;
        weights1[42375] <= 16'b0000000000000000;
        weights1[42376] <= 16'b0000000000000000;
        weights1[42377] <= 16'b0000000000000000;
        weights1[42378] <= 16'b0000000000000000;
        weights1[42379] <= 16'b0000000000000000;
        weights1[42380] <= 16'b0000000000000000;
        weights1[42381] <= 16'b0000000000000000;
        weights1[42382] <= 16'b0000000000000000;
        weights1[42383] <= 16'b0000000000000000;
        weights1[42384] <= 16'b0000000000000000;
        weights1[42385] <= 16'b0000000000000000;
        weights1[42386] <= 16'b0000000000000000;
        weights1[42387] <= 16'b0000000000000000;
        weights1[42388] <= 16'b0000000000000000;
        weights1[42389] <= 16'b0000000000000000;
        weights1[42390] <= 16'b0000000000000000;
        weights1[42391] <= 16'b0000000000000000;
        weights1[42392] <= 16'b0000000000000000;
        weights1[42393] <= 16'b0000000000000000;
        weights1[42394] <= 16'b0000000000000000;
        weights1[42395] <= 16'b0000000000000000;
        weights1[42396] <= 16'b0000000000000000;
        weights1[42397] <= 16'b0000000000000000;
        weights1[42398] <= 16'b0000000000000000;
        weights1[42399] <= 16'b0000000000000000;
        weights1[42400] <= 16'b0000000000000000;
        weights1[42401] <= 16'b0000000000000000;
        weights1[42402] <= 16'b0000000000000000;
        weights1[42403] <= 16'b0000000000000000;
        weights1[42404] <= 16'b0000000000000000;
        weights1[42405] <= 16'b0000000000000000;
        weights1[42406] <= 16'b0000000000000000;
        weights1[42407] <= 16'b0000000000000000;
        weights1[42408] <= 16'b0000000000000000;
        weights1[42409] <= 16'b0000000000000000;
        weights1[42410] <= 16'b0000000000000000;
        weights1[42411] <= 16'b0000000000000000;
        weights1[42412] <= 16'b0000000000000000;
        weights1[42413] <= 16'b0000000000000000;
        weights1[42414] <= 16'b0000000000000000;
        weights1[42415] <= 16'b0000000000000000;
        weights1[42416] <= 16'b0000000000000000;
        weights1[42417] <= 16'b0000000000000000;
        weights1[42418] <= 16'b0000000000000000;
        weights1[42419] <= 16'b0000000000000000;
        weights1[42420] <= 16'b0000000000000000;
        weights1[42421] <= 16'b0000000000000000;
        weights1[42422] <= 16'b0000000000000000;
        weights1[42423] <= 16'b0000000000000000;
        weights1[42424] <= 16'b0000000000000000;
        weights1[42425] <= 16'b0000000000000000;
        weights1[42426] <= 16'b0000000000000000;
        weights1[42427] <= 16'b0000000000000000;
        weights1[42428] <= 16'b0000000000000000;
        weights1[42429] <= 16'b0000000000000000;
        weights1[42430] <= 16'b0000000000000000;
        weights1[42431] <= 16'b0000000000000000;
        weights1[42432] <= 16'b0000000000000000;
        weights1[42433] <= 16'b0000000000000000;
        weights1[42434] <= 16'b0000000000000000;
        weights1[42435] <= 16'b0000000000000000;
        weights1[42436] <= 16'b0000000000000000;
        weights1[42437] <= 16'b0000000000000000;
        weights1[42438] <= 16'b0000000000000000;
        weights1[42439] <= 16'b0000000000000000;
        weights1[42440] <= 16'b0000000000000000;
        weights1[42441] <= 16'b0000000000000000;
        weights1[42442] <= 16'b0000000000000000;
        weights1[42443] <= 16'b0000000000000000;
        weights1[42444] <= 16'b0000000000000000;
        weights1[42445] <= 16'b0000000000000000;
        weights1[42446] <= 16'b0000000000000000;
        weights1[42447] <= 16'b0000000000000000;
        weights1[42448] <= 16'b0000000000000000;
        weights1[42449] <= 16'b0000000000000000;
        weights1[42450] <= 16'b0000000000000000;
        weights1[42451] <= 16'b0000000000000000;
        weights1[42452] <= 16'b0000000000000000;
        weights1[42453] <= 16'b0000000000000000;
        weights1[42454] <= 16'b0000000000000000;
        weights1[42455] <= 16'b0000000000000000;
        weights1[42456] <= 16'b0000000000000000;
        weights1[42457] <= 16'b0000000000000000;
        weights1[42458] <= 16'b0000000000000000;
        weights1[42459] <= 16'b0000000000000000;
        weights1[42460] <= 16'b0000000000000000;
        weights1[42461] <= 16'b0000000000000000;
        weights1[42462] <= 16'b0000000000000000;
        weights1[42463] <= 16'b0000000000000000;
        weights1[42464] <= 16'b0000000000000000;
        weights1[42465] <= 16'b0000000000000000;
        weights1[42466] <= 16'b0000000000000000;
        weights1[42467] <= 16'b0000000000000000;
        weights1[42468] <= 16'b0000000000000000;
        weights1[42469] <= 16'b0000000000000000;
        weights1[42470] <= 16'b0000000000000000;
        weights1[42471] <= 16'b0000000000000000;
        weights1[42472] <= 16'b0000000000000000;
        weights1[42473] <= 16'b0000000000000000;
        weights1[42474] <= 16'b0000000000000000;
        weights1[42475] <= 16'b0000000000000000;
        weights1[42476] <= 16'b0000000000000000;
        weights1[42477] <= 16'b0000000000000000;
        weights1[42478] <= 16'b0000000000000000;
        weights1[42479] <= 16'b0000000000000000;
        weights1[42480] <= 16'b0000000000000000;
        weights1[42481] <= 16'b0000000000000000;
        weights1[42482] <= 16'b0000000000000000;
        weights1[42483] <= 16'b0000000000000000;
        weights1[42484] <= 16'b0000000000000000;
        weights1[42485] <= 16'b0000000000000000;
        weights1[42486] <= 16'b0000000000000000;
        weights1[42487] <= 16'b0000000000000000;
        weights1[42488] <= 16'b0000000000000000;
        weights1[42489] <= 16'b0000000000000000;
        weights1[42490] <= 16'b0000000000000000;
        weights1[42491] <= 16'b0000000000000000;
        weights1[42492] <= 16'b0000000000000000;
        weights1[42493] <= 16'b0000000000000000;
        weights1[42494] <= 16'b0000000000000000;
        weights1[42495] <= 16'b0000000000000000;
        weights1[42496] <= 16'b0000000000000000;
        weights1[42497] <= 16'b0000000000000000;
        weights1[42498] <= 16'b0000000000000000;
        weights1[42499] <= 16'b0000000000000000;
        weights1[42500] <= 16'b0000000000000000;
        weights1[42501] <= 16'b0000000000000000;
        weights1[42502] <= 16'b0000000000000000;
        weights1[42503] <= 16'b0000000000000000;
        weights1[42504] <= 16'b0000000000000000;
        weights1[42505] <= 16'b0000000000000000;
        weights1[42506] <= 16'b0000000000000000;
        weights1[42507] <= 16'b0000000000000000;
        weights1[42508] <= 16'b0000000000000000;
        weights1[42509] <= 16'b0000000000000000;
        weights1[42510] <= 16'b0000000000000000;
        weights1[42511] <= 16'b0000000000000000;
        weights1[42512] <= 16'b0000000000000000;
        weights1[42513] <= 16'b0000000000000000;
        weights1[42514] <= 16'b0000000000000000;
        weights1[42515] <= 16'b0000000000000000;
        weights1[42516] <= 16'b0000000000000000;
        weights1[42517] <= 16'b0000000000000000;
        weights1[42518] <= 16'b0000000000000000;
        weights1[42519] <= 16'b0000000000000000;
        weights1[42520] <= 16'b0000000000000000;
        weights1[42521] <= 16'b0000000000000000;
        weights1[42522] <= 16'b0000000000000000;
        weights1[42523] <= 16'b0000000000000000;
        weights1[42524] <= 16'b0000000000000000;
        weights1[42525] <= 16'b0000000000000000;
        weights1[42526] <= 16'b0000000000000000;
        weights1[42527] <= 16'b0000000000000000;
        weights1[42528] <= 16'b0000000000000000;
        weights1[42529] <= 16'b0000000000000000;
        weights1[42530] <= 16'b0000000000000000;
        weights1[42531] <= 16'b0000000000000000;
        weights1[42532] <= 16'b0000000000000000;
        weights1[42533] <= 16'b0000000000000000;
        weights1[42534] <= 16'b0000000000000000;
        weights1[42535] <= 16'b0000000000000000;
        weights1[42536] <= 16'b0000000000000000;
        weights1[42537] <= 16'b0000000000000000;
        weights1[42538] <= 16'b0000000000000000;
        weights1[42539] <= 16'b0000000000000000;
        weights1[42540] <= 16'b0000000000000000;
        weights1[42541] <= 16'b0000000000000000;
        weights1[42542] <= 16'b0000000000000000;
        weights1[42543] <= 16'b0000000000000000;
        weights1[42544] <= 16'b0000000000000000;
        weights1[42545] <= 16'b0000000000000000;
        weights1[42546] <= 16'b0000000000000000;
        weights1[42547] <= 16'b0000000000000000;
        weights1[42548] <= 16'b0000000000000000;
        weights1[42549] <= 16'b0000000000000000;
        weights1[42550] <= 16'b0000000000000000;
        weights1[42551] <= 16'b0000000000000000;
        weights1[42552] <= 16'b0000000000000000;
        weights1[42553] <= 16'b0000000000000000;
        weights1[42554] <= 16'b0000000000000000;
        weights1[42555] <= 16'b0000000000000000;
        weights1[42556] <= 16'b0000000000000000;
        weights1[42557] <= 16'b0000000000000000;
        weights1[42558] <= 16'b0000000000000000;
        weights1[42559] <= 16'b0000000000000000;
        weights1[42560] <= 16'b0000000000000000;
        weights1[42561] <= 16'b0000000000000000;
        weights1[42562] <= 16'b0000000000000000;
        weights1[42563] <= 16'b0000000000000000;
        weights1[42564] <= 16'b0000000000000000;
        weights1[42565] <= 16'b0000000000000000;
        weights1[42566] <= 16'b0000000000000000;
        weights1[42567] <= 16'b0000000000000000;
        weights1[42568] <= 16'b0000000000000000;
        weights1[42569] <= 16'b0000000000000000;
        weights1[42570] <= 16'b0000000000000000;
        weights1[42571] <= 16'b0000000000000000;
        weights1[42572] <= 16'b0000000000000000;
        weights1[42573] <= 16'b0000000000000000;
        weights1[42574] <= 16'b0000000000000000;
        weights1[42575] <= 16'b0000000000000000;
        weights1[42576] <= 16'b0000000000000000;
        weights1[42577] <= 16'b0000000000000000;
        weights1[42578] <= 16'b0000000000000000;
        weights1[42579] <= 16'b0000000000000000;
        weights1[42580] <= 16'b0000000000000000;
        weights1[42581] <= 16'b0000000000000000;
        weights1[42582] <= 16'b0000000000000000;
        weights1[42583] <= 16'b0000000000000000;
        weights1[42584] <= 16'b0000000000000000;
        weights1[42585] <= 16'b0000000000000000;
        weights1[42586] <= 16'b0000000000000000;
        weights1[42587] <= 16'b0000000000000000;
        weights1[42588] <= 16'b0000000000000000;
        weights1[42589] <= 16'b0000000000000000;
        weights1[42590] <= 16'b0000000000000000;
        weights1[42591] <= 16'b0000000000000000;
        weights1[42592] <= 16'b0000000000000000;
        weights1[42593] <= 16'b0000000000000000;
        weights1[42594] <= 16'b0000000000000000;
        weights1[42595] <= 16'b0000000000000000;
        weights1[42596] <= 16'b0000000000000000;
        weights1[42597] <= 16'b0000000000000000;
        weights1[42598] <= 16'b0000000000000000;
        weights1[42599] <= 16'b0000000000000000;
        weights1[42600] <= 16'b0000000000000000;
        weights1[42601] <= 16'b0000000000000000;
        weights1[42602] <= 16'b0000000000000000;
        weights1[42603] <= 16'b0000000000000000;
        weights1[42604] <= 16'b0000000000000000;
        weights1[42605] <= 16'b0000000000000000;
        weights1[42606] <= 16'b0000000000000000;
        weights1[42607] <= 16'b0000000000000000;
        weights1[42608] <= 16'b0000000000000000;
        weights1[42609] <= 16'b0000000000000000;
        weights1[42610] <= 16'b0000000000000000;
        weights1[42611] <= 16'b0000000000000000;
        weights1[42612] <= 16'b0000000000000000;
        weights1[42613] <= 16'b0000000000000000;
        weights1[42614] <= 16'b0000000000000000;
        weights1[42615] <= 16'b0000000000000000;
        weights1[42616] <= 16'b0000000000000000;
        weights1[42617] <= 16'b0000000000000000;
        weights1[42618] <= 16'b0000000000000000;
        weights1[42619] <= 16'b0000000000000000;
        weights1[42620] <= 16'b0000000000000000;
        weights1[42621] <= 16'b0000000000000000;
        weights1[42622] <= 16'b0000000000000000;
        weights1[42623] <= 16'b0000000000000000;
        weights1[42624] <= 16'b0000000000000000;
        weights1[42625] <= 16'b0000000000000000;
        weights1[42626] <= 16'b0000000000000000;
        weights1[42627] <= 16'b0000000000000000;
        weights1[42628] <= 16'b0000000000000000;
        weights1[42629] <= 16'b0000000000000000;
        weights1[42630] <= 16'b0000000000000000;
        weights1[42631] <= 16'b0000000000000000;
        weights1[42632] <= 16'b0000000000000000;
        weights1[42633] <= 16'b0000000000000000;
        weights1[42634] <= 16'b0000000000000000;
        weights1[42635] <= 16'b0000000000000000;
        weights1[42636] <= 16'b0000000000000000;
        weights1[42637] <= 16'b0000000000000000;
        weights1[42638] <= 16'b0000000000000000;
        weights1[42639] <= 16'b0000000000000000;
        weights1[42640] <= 16'b0000000000000000;
        weights1[42641] <= 16'b0000000000000000;
        weights1[42642] <= 16'b0000000000000000;
        weights1[42643] <= 16'b0000000000000000;
        weights1[42644] <= 16'b0000000000000000;
        weights1[42645] <= 16'b0000000000000000;
        weights1[42646] <= 16'b0000000000000000;
        weights1[42647] <= 16'b0000000000000000;
        weights1[42648] <= 16'b0000000000000000;
        weights1[42649] <= 16'b0000000000000000;
        weights1[42650] <= 16'b0000000000000000;
        weights1[42651] <= 16'b0000000000000000;
        weights1[42652] <= 16'b0000000000000000;
        weights1[42653] <= 16'b0000000000000000;
        weights1[42654] <= 16'b0000000000000000;
        weights1[42655] <= 16'b0000000000000000;
        weights1[42656] <= 16'b0000000000000000;
        weights1[42657] <= 16'b0000000000000000;
        weights1[42658] <= 16'b0000000000000000;
        weights1[42659] <= 16'b0000000000000000;
        weights1[42660] <= 16'b0000000000000000;
        weights1[42661] <= 16'b0000000000000000;
        weights1[42662] <= 16'b0000000000000000;
        weights1[42663] <= 16'b0000000000000000;
        weights1[42664] <= 16'b0000000000000000;
        weights1[42665] <= 16'b0000000000000000;
        weights1[42666] <= 16'b0000000000000000;
        weights1[42667] <= 16'b0000000000000000;
        weights1[42668] <= 16'b0000000000000000;
        weights1[42669] <= 16'b0000000000000000;
        weights1[42670] <= 16'b0000000000000000;
        weights1[42671] <= 16'b0000000000000000;
        weights1[42672] <= 16'b0000000000000000;
        weights1[42673] <= 16'b0000000000000000;
        weights1[42674] <= 16'b0000000000000000;
        weights1[42675] <= 16'b0000000000000000;
        weights1[42676] <= 16'b0000000000000000;
        weights1[42677] <= 16'b0000000000000000;
        weights1[42678] <= 16'b0000000000000000;
        weights1[42679] <= 16'b0000000000000000;
        weights1[42680] <= 16'b0000000000000000;
        weights1[42681] <= 16'b0000000000000000;
        weights1[42682] <= 16'b0000000000000000;
        weights1[42683] <= 16'b0000000000000000;
        weights1[42684] <= 16'b0000000000000000;
        weights1[42685] <= 16'b0000000000000000;
        weights1[42686] <= 16'b0000000000000000;
        weights1[42687] <= 16'b0000000000000000;
        weights1[42688] <= 16'b0000000000000000;
        weights1[42689] <= 16'b0000000000000000;
        weights1[42690] <= 16'b0000000000000000;
        weights1[42691] <= 16'b0000000000000000;
        weights1[42692] <= 16'b0000000000000000;
        weights1[42693] <= 16'b0000000000000000;
        weights1[42694] <= 16'b0000000000000000;
        weights1[42695] <= 16'b0000000000000000;
        weights1[42696] <= 16'b0000000000000000;
        weights1[42697] <= 16'b0000000000000000;
        weights1[42698] <= 16'b0000000000000000;
        weights1[42699] <= 16'b0000000000000000;
        weights1[42700] <= 16'b0000000000000000;
        weights1[42701] <= 16'b0000000000000000;
        weights1[42702] <= 16'b0000000000000000;
        weights1[42703] <= 16'b0000000000000000;
        weights1[42704] <= 16'b0000000000000000;
        weights1[42705] <= 16'b0000000000000000;
        weights1[42706] <= 16'b0000000000000000;
        weights1[42707] <= 16'b0000000000000000;
        weights1[42708] <= 16'b0000000000000000;
        weights1[42709] <= 16'b0000000000000000;
        weights1[42710] <= 16'b0000000000000000;
        weights1[42711] <= 16'b0000000000000000;
        weights1[42712] <= 16'b0000000000000000;
        weights1[42713] <= 16'b0000000000000000;
        weights1[42714] <= 16'b0000000000000000;
        weights1[42715] <= 16'b0000000000000000;
        weights1[42716] <= 16'b0000000000000000;
        weights1[42717] <= 16'b0000000000000000;
        weights1[42718] <= 16'b0000000000000000;
        weights1[42719] <= 16'b0000000000000000;
        weights1[42720] <= 16'b0000000000000000;
        weights1[42721] <= 16'b0000000000000000;
        weights1[42722] <= 16'b0000000000000000;
        weights1[42723] <= 16'b0000000000000000;
        weights1[42724] <= 16'b0000000000000000;
        weights1[42725] <= 16'b0000000000000000;
        weights1[42726] <= 16'b0000000000000000;
        weights1[42727] <= 16'b0000000000000000;
        weights1[42728] <= 16'b0000000000000000;
        weights1[42729] <= 16'b0000000000000000;
        weights1[42730] <= 16'b0000000000000000;
        weights1[42731] <= 16'b0000000000000000;
        weights1[42732] <= 16'b0000000000000000;
        weights1[42733] <= 16'b0000000000000000;
        weights1[42734] <= 16'b0000000000000000;
        weights1[42735] <= 16'b0000000000000000;
        weights1[42736] <= 16'b0000000000000000;
        weights1[42737] <= 16'b0000000000000000;
        weights1[42738] <= 16'b0000000000000000;
        weights1[42739] <= 16'b0000000000000000;
        weights1[42740] <= 16'b0000000000000000;
        weights1[42741] <= 16'b0000000000000000;
        weights1[42742] <= 16'b0000000000000000;
        weights1[42743] <= 16'b0000000000000000;
        weights1[42744] <= 16'b0000000000000000;
        weights1[42745] <= 16'b0000000000000000;
        weights1[42746] <= 16'b0000000000000000;
        weights1[42747] <= 16'b0000000000000000;
        weights1[42748] <= 16'b0000000000000000;
        weights1[42749] <= 16'b0000000000000000;
        weights1[42750] <= 16'b0000000000000000;
        weights1[42751] <= 16'b0000000000000000;
        weights1[42752] <= 16'b0000000000000000;
        weights1[42753] <= 16'b0000000000000000;
        weights1[42754] <= 16'b0000000000000000;
        weights1[42755] <= 16'b0000000000000000;
        weights1[42756] <= 16'b0000000000000000;
        weights1[42757] <= 16'b0000000000000000;
        weights1[42758] <= 16'b0000000000000000;
        weights1[42759] <= 16'b0000000000000000;
        weights1[42760] <= 16'b0000000000000000;
        weights1[42761] <= 16'b0000000000000000;
        weights1[42762] <= 16'b0000000000000000;
        weights1[42763] <= 16'b0000000000000000;
        weights1[42764] <= 16'b0000000000000000;
        weights1[42765] <= 16'b0000000000000000;
        weights1[42766] <= 16'b0000000000000000;
        weights1[42767] <= 16'b0000000000000000;
        weights1[42768] <= 16'b0000000000000000;
        weights1[42769] <= 16'b0000000000000000;
        weights1[42770] <= 16'b0000000000000000;
        weights1[42771] <= 16'b0000000000000000;
        weights1[42772] <= 16'b0000000000000000;
        weights1[42773] <= 16'b0000000000000000;
        weights1[42774] <= 16'b0000000000000000;
        weights1[42775] <= 16'b0000000000000000;
        weights1[42776] <= 16'b0000000000000000;
        weights1[42777] <= 16'b0000000000000000;
        weights1[42778] <= 16'b0000000000000000;
        weights1[42779] <= 16'b0000000000000000;
        weights1[42780] <= 16'b0000000000000000;
        weights1[42781] <= 16'b0000000000000000;
        weights1[42782] <= 16'b0000000000000000;
        weights1[42783] <= 16'b0000000000000000;
        weights1[42784] <= 16'b0000000000000000;
        weights1[42785] <= 16'b0000000000000000;
        weights1[42786] <= 16'b0000000000000000;
        weights1[42787] <= 16'b0000000000000000;
        weights1[42788] <= 16'b0000000000000000;
        weights1[42789] <= 16'b0000000000000000;
        weights1[42790] <= 16'b0000000000000000;
        weights1[42791] <= 16'b0000000000000000;
        weights1[42792] <= 16'b0000000000000000;
        weights1[42793] <= 16'b0000000000000000;
        weights1[42794] <= 16'b0000000000000000;
        weights1[42795] <= 16'b0000000000000000;
        weights1[42796] <= 16'b0000000000000000;
        weights1[42797] <= 16'b0000000000000000;
        weights1[42798] <= 16'b0000000000000000;
        weights1[42799] <= 16'b0000000000000000;
        weights1[42800] <= 16'b0000000000000000;
        weights1[42801] <= 16'b0000000000000000;
        weights1[42802] <= 16'b0000000000000000;
        weights1[42803] <= 16'b0000000000000000;
        weights1[42804] <= 16'b0000000000000000;
        weights1[42805] <= 16'b0000000000000000;
        weights1[42806] <= 16'b0000000000000000;
        weights1[42807] <= 16'b0000000000000000;
        weights1[42808] <= 16'b0000000000000000;
        weights1[42809] <= 16'b0000000000000000;
        weights1[42810] <= 16'b0000000000000000;
        weights1[42811] <= 16'b0000000000000000;
        weights1[42812] <= 16'b0000000000000000;
        weights1[42813] <= 16'b0000000000000000;
        weights1[42814] <= 16'b0000000000000000;
        weights1[42815] <= 16'b0000000000000000;
        weights1[42816] <= 16'b0000000000000000;
        weights1[42817] <= 16'b0000000000000000;
        weights1[42818] <= 16'b0000000000000000;
        weights1[42819] <= 16'b0000000000000000;
        weights1[42820] <= 16'b0000000000000000;
        weights1[42821] <= 16'b0000000000000000;
        weights1[42822] <= 16'b0000000000000000;
        weights1[42823] <= 16'b0000000000000000;
        weights1[42824] <= 16'b0000000000000000;
        weights1[42825] <= 16'b0000000000000000;
        weights1[42826] <= 16'b0000000000000000;
        weights1[42827] <= 16'b0000000000000000;
        weights1[42828] <= 16'b0000000000000000;
        weights1[42829] <= 16'b0000000000000000;
        weights1[42830] <= 16'b0000000000000000;
        weights1[42831] <= 16'b0000000000000000;
        weights1[42832] <= 16'b0000000000000000;
        weights1[42833] <= 16'b0000000000000000;
        weights1[42834] <= 16'b0000000000000000;
        weights1[42835] <= 16'b0000000000000000;
        weights1[42836] <= 16'b0000000000000000;
        weights1[42837] <= 16'b0000000000000000;
        weights1[42838] <= 16'b0000000000000000;
        weights1[42839] <= 16'b0000000000000000;
        weights1[42840] <= 16'b0000000000000000;
        weights1[42841] <= 16'b0000000000000000;
        weights1[42842] <= 16'b0000000000000000;
        weights1[42843] <= 16'b0000000000000000;
        weights1[42844] <= 16'b0000000000000000;
        weights1[42845] <= 16'b0000000000000000;
        weights1[42846] <= 16'b0000000000000000;
        weights1[42847] <= 16'b0000000000000000;
        weights1[42848] <= 16'b0000000000000000;
        weights1[42849] <= 16'b0000000000000000;
        weights1[42850] <= 16'b0000000000000000;
        weights1[42851] <= 16'b0000000000000000;
        weights1[42852] <= 16'b0000000000000000;
        weights1[42853] <= 16'b0000000000000000;
        weights1[42854] <= 16'b0000000000000000;
        weights1[42855] <= 16'b0000000000000000;
        weights1[42856] <= 16'b0000000000000000;
        weights1[42857] <= 16'b0000000000000000;
        weights1[42858] <= 16'b0000000000000000;
        weights1[42859] <= 16'b0000000000000000;
        weights1[42860] <= 16'b0000000000000000;
        weights1[42861] <= 16'b0000000000000000;
        weights1[42862] <= 16'b0000000000000000;
        weights1[42863] <= 16'b0000000000000000;
        weights1[42864] <= 16'b0000000000000000;
        weights1[42865] <= 16'b0000000000000000;
        weights1[42866] <= 16'b0000000000000000;
        weights1[42867] <= 16'b0000000000000000;
        weights1[42868] <= 16'b0000000000000000;
        weights1[42869] <= 16'b0000000000000000;
        weights1[42870] <= 16'b0000000000000000;
        weights1[42871] <= 16'b0000000000000000;
        weights1[42872] <= 16'b0000000000000000;
        weights1[42873] <= 16'b0000000000000000;
        weights1[42874] <= 16'b0000000000000000;
        weights1[42875] <= 16'b0000000000000000;
        weights1[42876] <= 16'b0000000000000000;
        weights1[42877] <= 16'b0000000000000000;
        weights1[42878] <= 16'b0000000000000000;
        weights1[42879] <= 16'b0000000000000000;
        weights1[42880] <= 16'b0000000000000000;
        weights1[42881] <= 16'b0000000000000000;
        weights1[42882] <= 16'b0000000000000000;
        weights1[42883] <= 16'b0000000000000000;
        weights1[42884] <= 16'b0000000000000000;
        weights1[42885] <= 16'b0000000000000000;
        weights1[42886] <= 16'b0000000000000000;
        weights1[42887] <= 16'b0000000000000000;
        weights1[42888] <= 16'b0000000000000000;
        weights1[42889] <= 16'b0000000000000000;
        weights1[42890] <= 16'b0000000000000000;
        weights1[42891] <= 16'b0000000000000000;
        weights1[42892] <= 16'b0000000000000000;
        weights1[42893] <= 16'b0000000000000000;
        weights1[42894] <= 16'b0000000000000000;
        weights1[42895] <= 16'b0000000000000000;
        weights1[42896] <= 16'b0000000000000000;
        weights1[42897] <= 16'b0000000000000000;
        weights1[42898] <= 16'b0000000000000000;
        weights1[42899] <= 16'b0000000000000000;
        weights1[42900] <= 16'b0000000000000000;
        weights1[42901] <= 16'b0000000000000000;
        weights1[42902] <= 16'b0000000000000000;
        weights1[42903] <= 16'b0000000000000000;
        weights1[42904] <= 16'b0000000000000000;
        weights1[42905] <= 16'b0000000000000000;
        weights1[42906] <= 16'b0000000000000000;
        weights1[42907] <= 16'b0000000000000000;
        weights1[42908] <= 16'b0000000000000000;
        weights1[42909] <= 16'b0000000000000000;
        weights1[42910] <= 16'b0000000000000000;
        weights1[42911] <= 16'b0000000000000000;
        weights1[42912] <= 16'b0000000000000000;
        weights1[42913] <= 16'b0000000000000000;
        weights1[42914] <= 16'b0000000000000000;
        weights1[42915] <= 16'b0000000000000000;
        weights1[42916] <= 16'b0000000000000000;
        weights1[42917] <= 16'b0000000000000000;
        weights1[42918] <= 16'b0000000000000000;
        weights1[42919] <= 16'b0000000000000000;
        weights1[42920] <= 16'b0000000000000000;
        weights1[42921] <= 16'b0000000000000000;
        weights1[42922] <= 16'b0000000000000000;
        weights1[42923] <= 16'b0000000000000000;
        weights1[42924] <= 16'b0000000000000000;
        weights1[42925] <= 16'b0000000000000000;
        weights1[42926] <= 16'b0000000000000000;
        weights1[42927] <= 16'b0000000000000000;
        weights1[42928] <= 16'b0000000000000000;
        weights1[42929] <= 16'b0000000000000000;
        weights1[42930] <= 16'b0000000000000000;
        weights1[42931] <= 16'b0000000000000000;
        weights1[42932] <= 16'b0000000000000000;
        weights1[42933] <= 16'b0000000000000000;
        weights1[42934] <= 16'b0000000000000000;
        weights1[42935] <= 16'b0000000000000000;
        weights1[42936] <= 16'b0000000000000000;
        weights1[42937] <= 16'b0000000000000000;
        weights1[42938] <= 16'b0000000000000000;
        weights1[42939] <= 16'b0000000000000000;
        weights1[42940] <= 16'b0000000000000000;
        weights1[42941] <= 16'b0000000000000000;
        weights1[42942] <= 16'b0000000000000000;
        weights1[42943] <= 16'b0000000000000000;
        weights1[42944] <= 16'b0000000000000000;
        weights1[42945] <= 16'b0000000000000000;
        weights1[42946] <= 16'b0000000000000000;
        weights1[42947] <= 16'b0000000000000000;
        weights1[42948] <= 16'b0000000000000000;
        weights1[42949] <= 16'b0000000000000000;
        weights1[42950] <= 16'b0000000000000000;
        weights1[42951] <= 16'b0000000000000000;
        weights1[42952] <= 16'b0000000000000000;
        weights1[42953] <= 16'b0000000000000000;
        weights1[42954] <= 16'b0000000000000000;
        weights1[42955] <= 16'b0000000000000000;
        weights1[42956] <= 16'b0000000000000000;
        weights1[42957] <= 16'b0000000000000000;
        weights1[42958] <= 16'b0000000000000000;
        weights1[42959] <= 16'b0000000000000000;
        weights1[42960] <= 16'b0000000000000000;
        weights1[42961] <= 16'b0000000000000000;
        weights1[42962] <= 16'b0000000000000000;
        weights1[42963] <= 16'b0000000000000000;
        weights1[42964] <= 16'b0000000000000000;
        weights1[42965] <= 16'b0000000000000000;
        weights1[42966] <= 16'b0000000000000000;
        weights1[42967] <= 16'b0000000000000000;
        weights1[42968] <= 16'b0000000000000000;
        weights1[42969] <= 16'b0000000000000000;
        weights1[42970] <= 16'b0000000000000000;
        weights1[42971] <= 16'b0000000000000000;
        weights1[42972] <= 16'b0000000000000000;
        weights1[42973] <= 16'b0000000000000000;
        weights1[42974] <= 16'b0000000000000000;
        weights1[42975] <= 16'b0000000000000000;
        weights1[42976] <= 16'b0000000000000000;
        weights1[42977] <= 16'b0000000000000000;
        weights1[42978] <= 16'b0000000000000000;
        weights1[42979] <= 16'b0000000000000000;
        weights1[42980] <= 16'b0000000000000000;
        weights1[42981] <= 16'b0000000000000000;
        weights1[42982] <= 16'b0000000000000000;
        weights1[42983] <= 16'b0000000000000000;
        weights1[42984] <= 16'b0000000000000000;
        weights1[42985] <= 16'b0000000000000000;
        weights1[42986] <= 16'b0000000000000000;
        weights1[42987] <= 16'b0000000000000000;
        weights1[42988] <= 16'b0000000000000000;
        weights1[42989] <= 16'b0000000000000000;
        weights1[42990] <= 16'b0000000000000000;
        weights1[42991] <= 16'b0000000000000000;
        weights1[42992] <= 16'b0000000000000000;
        weights1[42993] <= 16'b0000000000000000;
        weights1[42994] <= 16'b0000000000000000;
        weights1[42995] <= 16'b0000000000000000;
        weights1[42996] <= 16'b0000000000000000;
        weights1[42997] <= 16'b0000000000000000;
        weights1[42998] <= 16'b0000000000000000;
        weights1[42999] <= 16'b0000000000000000;
        weights1[43000] <= 16'b0000000000000000;
        weights1[43001] <= 16'b0000000000000000;
        weights1[43002] <= 16'b0000000000000000;
        weights1[43003] <= 16'b0000000000000000;
        weights1[43004] <= 16'b0000000000000000;
        weights1[43005] <= 16'b0000000000000000;
        weights1[43006] <= 16'b0000000000000000;
        weights1[43007] <= 16'b0000000000000000;
        weights1[43008] <= 16'b0000000000000000;
        weights1[43009] <= 16'b0000000000000000;
        weights1[43010] <= 16'b0000000000000000;
        weights1[43011] <= 16'b0000000000000000;
        weights1[43012] <= 16'b0000000000000000;
        weights1[43013] <= 16'b0000000000000000;
        weights1[43014] <= 16'b0000000000000000;
        weights1[43015] <= 16'b0000000000000000;
        weights1[43016] <= 16'b0000000000000000;
        weights1[43017] <= 16'b0000000000000000;
        weights1[43018] <= 16'b0000000000000000;
        weights1[43019] <= 16'b0000000000000000;
        weights1[43020] <= 16'b0000000000000000;
        weights1[43021] <= 16'b0000000000000000;
        weights1[43022] <= 16'b0000000000000000;
        weights1[43023] <= 16'b0000000000000000;
        weights1[43024] <= 16'b0000000000000000;
        weights1[43025] <= 16'b0000000000000000;
        weights1[43026] <= 16'b0000000000000000;
        weights1[43027] <= 16'b0000000000000000;
        weights1[43028] <= 16'b0000000000000000;
        weights1[43029] <= 16'b0000000000000000;
        weights1[43030] <= 16'b0000000000000000;
        weights1[43031] <= 16'b0000000000000000;
        weights1[43032] <= 16'b0000000000000000;
        weights1[43033] <= 16'b0000000000000000;
        weights1[43034] <= 16'b0000000000000000;
        weights1[43035] <= 16'b0000000000000000;
        weights1[43036] <= 16'b0000000000000000;
        weights1[43037] <= 16'b0000000000000000;
        weights1[43038] <= 16'b0000000000000000;
        weights1[43039] <= 16'b0000000000000000;
        weights1[43040] <= 16'b0000000000000000;
        weights1[43041] <= 16'b0000000000000000;
        weights1[43042] <= 16'b0000000000000000;
        weights1[43043] <= 16'b0000000000000000;
        weights1[43044] <= 16'b0000000000000000;
        weights1[43045] <= 16'b0000000000000000;
        weights1[43046] <= 16'b0000000000000000;
        weights1[43047] <= 16'b0000000000000000;
        weights1[43048] <= 16'b0000000000000000;
        weights1[43049] <= 16'b0000000000000000;
        weights1[43050] <= 16'b0000000000000000;
        weights1[43051] <= 16'b0000000000000000;
        weights1[43052] <= 16'b0000000000000000;
        weights1[43053] <= 16'b0000000000000000;
        weights1[43054] <= 16'b0000000000000000;
        weights1[43055] <= 16'b0000000000000000;
        weights1[43056] <= 16'b0000000000000000;
        weights1[43057] <= 16'b0000000000000000;
        weights1[43058] <= 16'b0000000000000000;
        weights1[43059] <= 16'b0000000000000000;
        weights1[43060] <= 16'b0000000000000000;
        weights1[43061] <= 16'b0000000000000000;
        weights1[43062] <= 16'b0000000000000000;
        weights1[43063] <= 16'b0000000000000000;
        weights1[43064] <= 16'b0000000000000000;
        weights1[43065] <= 16'b0000000000000000;
        weights1[43066] <= 16'b0000000000000000;
        weights1[43067] <= 16'b0000000000000000;
        weights1[43068] <= 16'b0000000000000000;
        weights1[43069] <= 16'b0000000000000000;
        weights1[43070] <= 16'b0000000000000000;
        weights1[43071] <= 16'b0000000000000000;
        weights1[43072] <= 16'b0000000000000000;
        weights1[43073] <= 16'b0000000000000000;
        weights1[43074] <= 16'b0000000000000000;
        weights1[43075] <= 16'b0000000000000000;
        weights1[43076] <= 16'b0000000000000000;
        weights1[43077] <= 16'b0000000000000000;
        weights1[43078] <= 16'b0000000000000000;
        weights1[43079] <= 16'b0000000000000000;
        weights1[43080] <= 16'b0000000000000000;
        weights1[43081] <= 16'b0000000000000000;
        weights1[43082] <= 16'b0000000000000000;
        weights1[43083] <= 16'b0000000000000000;
        weights1[43084] <= 16'b0000000000000000;
        weights1[43085] <= 16'b0000000000000000;
        weights1[43086] <= 16'b0000000000000000;
        weights1[43087] <= 16'b0000000000000000;
        weights1[43088] <= 16'b0000000000000000;
        weights1[43089] <= 16'b0000000000000000;
        weights1[43090] <= 16'b0000000000000000;
        weights1[43091] <= 16'b0000000000000000;
        weights1[43092] <= 16'b0000000000000000;
        weights1[43093] <= 16'b0000000000000000;
        weights1[43094] <= 16'b0000000000000000;
        weights1[43095] <= 16'b0000000000000000;
        weights1[43096] <= 16'b0000000000000000;
        weights1[43097] <= 16'b0000000000000000;
        weights1[43098] <= 16'b0000000000000000;
        weights1[43099] <= 16'b0000000000000000;
        weights1[43100] <= 16'b0000000000000000;
        weights1[43101] <= 16'b0000000000000000;
        weights1[43102] <= 16'b0000000000000000;
        weights1[43103] <= 16'b0000000000000000;
        weights1[43104] <= 16'b0000000000000000;
        weights1[43105] <= 16'b0000000000000000;
        weights1[43106] <= 16'b0000000000000000;
        weights1[43107] <= 16'b0000000000000000;
        weights1[43108] <= 16'b0000000000000000;
        weights1[43109] <= 16'b0000000000000000;
        weights1[43110] <= 16'b0000000000000000;
        weights1[43111] <= 16'b0000000000000000;
        weights1[43112] <= 16'b0000000000000000;
        weights1[43113] <= 16'b0000000000000000;
        weights1[43114] <= 16'b0000000000000000;
        weights1[43115] <= 16'b0000000000000000;
        weights1[43116] <= 16'b0000000000000000;
        weights1[43117] <= 16'b0000000000000000;
        weights1[43118] <= 16'b0000000000000000;
        weights1[43119] <= 16'b0000000000000000;
        weights1[43120] <= 16'b0000000000000000;
        weights1[43121] <= 16'b1111111111111111;
        weights1[43122] <= 16'b1111111111111111;
        weights1[43123] <= 16'b0000000000000000;
        weights1[43124] <= 16'b0000000000000000;
        weights1[43125] <= 16'b0000000000000000;
        weights1[43126] <= 16'b0000000000000000;
        weights1[43127] <= 16'b1111111111111111;
        weights1[43128] <= 16'b1111111111111111;
        weights1[43129] <= 16'b1111111111111110;
        weights1[43130] <= 16'b0000000000000001;
        weights1[43131] <= 16'b1111111111111010;
        weights1[43132] <= 16'b1111111111111010;
        weights1[43133] <= 16'b1111111111111101;
        weights1[43134] <= 16'b1111111111111110;
        weights1[43135] <= 16'b1111111111111100;
        weights1[43136] <= 16'b1111111111110110;
        weights1[43137] <= 16'b1111111111110100;
        weights1[43138] <= 16'b1111111111110110;
        weights1[43139] <= 16'b1111111111110110;
        weights1[43140] <= 16'b1111111111110101;
        weights1[43141] <= 16'b1111111111111000;
        weights1[43142] <= 16'b1111111111111010;
        weights1[43143] <= 16'b1111111111111100;
        weights1[43144] <= 16'b1111111111111101;
        weights1[43145] <= 16'b1111111111111111;
        weights1[43146] <= 16'b0000000000000000;
        weights1[43147] <= 16'b0000000000000000;
        weights1[43148] <= 16'b0000000000000000;
        weights1[43149] <= 16'b1111111111111110;
        weights1[43150] <= 16'b1111111111111110;
        weights1[43151] <= 16'b1111111111111111;
        weights1[43152] <= 16'b0000000000000000;
        weights1[43153] <= 16'b0000000000000100;
        weights1[43154] <= 16'b0000000000000101;
        weights1[43155] <= 16'b0000000000000010;
        weights1[43156] <= 16'b1111111111111100;
        weights1[43157] <= 16'b1111111111110111;
        weights1[43158] <= 16'b1111111111111011;
        weights1[43159] <= 16'b1111111111111011;
        weights1[43160] <= 16'b1111111111111010;
        weights1[43161] <= 16'b1111111111101111;
        weights1[43162] <= 16'b1111111111101110;
        weights1[43163] <= 16'b1111111111101100;
        weights1[43164] <= 16'b1111111111101111;
        weights1[43165] <= 16'b1111111111100111;
        weights1[43166] <= 16'b1111111111101001;
        weights1[43167] <= 16'b1111111111101110;
        weights1[43168] <= 16'b1111111111110001;
        weights1[43169] <= 16'b1111111111110101;
        weights1[43170] <= 16'b1111111111111000;
        weights1[43171] <= 16'b1111111111111001;
        weights1[43172] <= 16'b1111111111111100;
        weights1[43173] <= 16'b1111111111111111;
        weights1[43174] <= 16'b0000000000000001;
        weights1[43175] <= 16'b0000000000000000;
        weights1[43176] <= 16'b1111111111111111;
        weights1[43177] <= 16'b1111111111111111;
        weights1[43178] <= 16'b0000000000000001;
        weights1[43179] <= 16'b0000000000000000;
        weights1[43180] <= 16'b0000000000000010;
        weights1[43181] <= 16'b0000000000000100;
        weights1[43182] <= 16'b0000000000001011;
        weights1[43183] <= 16'b1111111111111110;
        weights1[43184] <= 16'b1111111111111001;
        weights1[43185] <= 16'b1111111111111000;
        weights1[43186] <= 16'b1111111111111010;
        weights1[43187] <= 16'b1111111111111000;
        weights1[43188] <= 16'b1111111111110001;
        weights1[43189] <= 16'b1111111111101011;
        weights1[43190] <= 16'b1111111111101100;
        weights1[43191] <= 16'b1111111111100100;
        weights1[43192] <= 16'b1111111111101010;
        weights1[43193] <= 16'b1111111111100110;
        weights1[43194] <= 16'b1111111111101100;
        weights1[43195] <= 16'b1111111111100101;
        weights1[43196] <= 16'b1111111111101001;
        weights1[43197] <= 16'b1111111111101001;
        weights1[43198] <= 16'b1111111111110001;
        weights1[43199] <= 16'b1111111111110111;
        weights1[43200] <= 16'b1111111111111111;
        weights1[43201] <= 16'b1111111111111111;
        weights1[43202] <= 16'b1111111111111110;
        weights1[43203] <= 16'b1111111111111110;
        weights1[43204] <= 16'b1111111111111111;
        weights1[43205] <= 16'b1111111111111110;
        weights1[43206] <= 16'b1111111111111111;
        weights1[43207] <= 16'b1111111111111110;
        weights1[43208] <= 16'b0000000000000000;
        weights1[43209] <= 16'b0000000000000010;
        weights1[43210] <= 16'b1111111111111111;
        weights1[43211] <= 16'b1111111111111110;
        weights1[43212] <= 16'b1111111111110100;
        weights1[43213] <= 16'b1111111111111110;
        weights1[43214] <= 16'b1111111111110101;
        weights1[43215] <= 16'b0000000000000010;
        weights1[43216] <= 16'b1111111111111100;
        weights1[43217] <= 16'b0000000000000110;
        weights1[43218] <= 16'b1111111111111101;
        weights1[43219] <= 16'b1111111111110001;
        weights1[43220] <= 16'b1111111111100011;
        weights1[43221] <= 16'b1111111111100011;
        weights1[43222] <= 16'b1111111111011100;
        weights1[43223] <= 16'b1111111111010111;
        weights1[43224] <= 16'b1111111111011110;
        weights1[43225] <= 16'b1111111111100011;
        weights1[43226] <= 16'b1111111111100101;
        weights1[43227] <= 16'b1111111111110110;
        weights1[43228] <= 16'b1111111111111000;
        weights1[43229] <= 16'b1111111111111011;
        weights1[43230] <= 16'b1111111111111000;
        weights1[43231] <= 16'b1111111111111010;
        weights1[43232] <= 16'b1111111111111111;
        weights1[43233] <= 16'b1111111111111110;
        weights1[43234] <= 16'b1111111111111110;
        weights1[43235] <= 16'b0000000000000001;
        weights1[43236] <= 16'b1111111111111100;
        weights1[43237] <= 16'b1111111111111100;
        weights1[43238] <= 16'b1111111111110111;
        weights1[43239] <= 16'b1111111111111000;
        weights1[43240] <= 16'b1111111111111000;
        weights1[43241] <= 16'b1111111111100011;
        weights1[43242] <= 16'b1111111111101000;
        weights1[43243] <= 16'b1111111111100100;
        weights1[43244] <= 16'b1111111111100010;
        weights1[43245] <= 16'b0000000000000001;
        weights1[43246] <= 16'b0000000000010001;
        weights1[43247] <= 16'b1111111111101010;
        weights1[43248] <= 16'b1111111111100000;
        weights1[43249] <= 16'b1111111111110011;
        weights1[43250] <= 16'b1111111111110100;
        weights1[43251] <= 16'b1111111111110000;
        weights1[43252] <= 16'b1111111111110010;
        weights1[43253] <= 16'b1111111111011110;
        weights1[43254] <= 16'b1111111111100101;
        weights1[43255] <= 16'b1111111111101001;
        weights1[43256] <= 16'b1111111111101101;
        weights1[43257] <= 16'b1111111111110010;
        weights1[43258] <= 16'b1111111111110100;
        weights1[43259] <= 16'b1111111111111100;
        weights1[43260] <= 16'b1111111111111111;
        weights1[43261] <= 16'b0000000000000001;
        weights1[43262] <= 16'b1111111111111010;
        weights1[43263] <= 16'b1111111111111010;
        weights1[43264] <= 16'b1111111111111100;
        weights1[43265] <= 16'b1111111111100101;
        weights1[43266] <= 16'b1111111111111000;
        weights1[43267] <= 16'b1111111111101110;
        weights1[43268] <= 16'b1111111111100000;
        weights1[43269] <= 16'b1111111111101010;
        weights1[43270] <= 16'b0000000000000010;
        weights1[43271] <= 16'b0000000000001101;
        weights1[43272] <= 16'b0000000000000100;
        weights1[43273] <= 16'b0000000000010000;
        weights1[43274] <= 16'b1111111111101000;
        weights1[43275] <= 16'b1111111111011011;
        weights1[43276] <= 16'b1111111111101010;
        weights1[43277] <= 16'b0000000000000000;
        weights1[43278] <= 16'b0000000000010011;
        weights1[43279] <= 16'b1111111111100100;
        weights1[43280] <= 16'b1111111111101100;
        weights1[43281] <= 16'b1111111111110111;
        weights1[43282] <= 16'b1111111111011111;
        weights1[43283] <= 16'b1111111111101010;
        weights1[43284] <= 16'b1111111111101011;
        weights1[43285] <= 16'b1111111111110011;
        weights1[43286] <= 16'b1111111111110100;
        weights1[43287] <= 16'b0000000000000000;
        weights1[43288] <= 16'b1111111111111111;
        weights1[43289] <= 16'b1111111111111111;
        weights1[43290] <= 16'b1111111111101010;
        weights1[43291] <= 16'b1111111111101111;
        weights1[43292] <= 16'b1111111111110100;
        weights1[43293] <= 16'b1111111111101010;
        weights1[43294] <= 16'b0000000000001111;
        weights1[43295] <= 16'b1111111111111111;
        weights1[43296] <= 16'b1111111111101101;
        weights1[43297] <= 16'b0000000000000001;
        weights1[43298] <= 16'b0000000000010111;
        weights1[43299] <= 16'b1111111111111011;
        weights1[43300] <= 16'b1111111111110011;
        weights1[43301] <= 16'b1111111111111100;
        weights1[43302] <= 16'b1111111111111111;
        weights1[43303] <= 16'b1111111111100000;
        weights1[43304] <= 16'b1111111111101111;
        weights1[43305] <= 16'b1111111111111100;
        weights1[43306] <= 16'b1111111111011011;
        weights1[43307] <= 16'b0000000000000101;
        weights1[43308] <= 16'b1111111111101110;
        weights1[43309] <= 16'b1111111111101101;
        weights1[43310] <= 16'b1111111111011000;
        weights1[43311] <= 16'b1111111111011011;
        weights1[43312] <= 16'b1111111111110000;
        weights1[43313] <= 16'b1111111111100100;
        weights1[43314] <= 16'b1111111111110011;
        weights1[43315] <= 16'b1111111111111100;
        weights1[43316] <= 16'b0000000000000000;
        weights1[43317] <= 16'b1111111111111110;
        weights1[43318] <= 16'b1111111111110001;
        weights1[43319] <= 16'b1111111111110011;
        weights1[43320] <= 16'b1111111111101000;
        weights1[43321] <= 16'b1111111111111000;
        weights1[43322] <= 16'b0000000000001101;
        weights1[43323] <= 16'b1111111111100100;
        weights1[43324] <= 16'b0000000000011000;
        weights1[43325] <= 16'b1111111111110101;
        weights1[43326] <= 16'b0000000000001000;
        weights1[43327] <= 16'b0000000000000010;
        weights1[43328] <= 16'b0000000000001001;
        weights1[43329] <= 16'b0000000000010010;
        weights1[43330] <= 16'b0000000000000100;
        weights1[43331] <= 16'b1111111111111011;
        weights1[43332] <= 16'b0000000000011001;
        weights1[43333] <= 16'b1111111111101101;
        weights1[43334] <= 16'b1111111111110010;
        weights1[43335] <= 16'b1111111111110010;
        weights1[43336] <= 16'b0000000000000010;
        weights1[43337] <= 16'b0000000000000011;
        weights1[43338] <= 16'b1111111111110001;
        weights1[43339] <= 16'b1111111111101101;
        weights1[43340] <= 16'b1111111111110000;
        weights1[43341] <= 16'b1111111111100011;
        weights1[43342] <= 16'b1111111111110001;
        weights1[43343] <= 16'b1111111111110100;
        weights1[43344] <= 16'b0000000000000001;
        weights1[43345] <= 16'b1111111111111100;
        weights1[43346] <= 16'b0000000000000000;
        weights1[43347] <= 16'b1111111111101010;
        weights1[43348] <= 16'b1111111111110110;
        weights1[43349] <= 16'b1111111111110010;
        weights1[43350] <= 16'b1111111111111011;
        weights1[43351] <= 16'b1111111111111001;
        weights1[43352] <= 16'b1111111111111111;
        weights1[43353] <= 16'b1111111111110011;
        weights1[43354] <= 16'b1111111111110011;
        weights1[43355] <= 16'b0000000000000110;
        weights1[43356] <= 16'b0000000000000010;
        weights1[43357] <= 16'b0000000000001100;
        weights1[43358] <= 16'b1111111111111001;
        weights1[43359] <= 16'b0000000000010000;
        weights1[43360] <= 16'b0000000000001101;
        weights1[43361] <= 16'b0000000000001100;
        weights1[43362] <= 16'b1111111111100100;
        weights1[43363] <= 16'b0000000000010011;
        weights1[43364] <= 16'b1111111111101100;
        weights1[43365] <= 16'b1111111111110000;
        weights1[43366] <= 16'b0000000000000010;
        weights1[43367] <= 16'b0000000000001001;
        weights1[43368] <= 16'b1111111111101100;
        weights1[43369] <= 16'b1111111111110110;
        weights1[43370] <= 16'b1111111111101100;
        weights1[43371] <= 16'b1111111111110110;
        weights1[43372] <= 16'b0000000000000000;
        weights1[43373] <= 16'b1111111111111101;
        weights1[43374] <= 16'b1111111111111110;
        weights1[43375] <= 16'b1111111111110011;
        weights1[43376] <= 16'b1111111111110111;
        weights1[43377] <= 16'b0000000000000110;
        weights1[43378] <= 16'b1111111111011000;
        weights1[43379] <= 16'b1111111111110001;
        weights1[43380] <= 16'b0000000000000000;
        weights1[43381] <= 16'b1111111111111000;
        weights1[43382] <= 16'b1111111111111011;
        weights1[43383] <= 16'b1111111111111110;
        weights1[43384] <= 16'b1111111111100101;
        weights1[43385] <= 16'b1111111111110001;
        weights1[43386] <= 16'b0000000000001011;
        weights1[43387] <= 16'b0000000000000000;
        weights1[43388] <= 16'b1111111111111111;
        weights1[43389] <= 16'b1111111111110001;
        weights1[43390] <= 16'b1111111111111010;
        weights1[43391] <= 16'b1111111111111011;
        weights1[43392] <= 16'b1111111111110111;
        weights1[43393] <= 16'b0000000000001101;
        weights1[43394] <= 16'b0000000000010001;
        weights1[43395] <= 16'b1111111111111011;
        weights1[43396] <= 16'b1111111111011110;
        weights1[43397] <= 16'b1111111111101010;
        weights1[43398] <= 16'b1111111111110010;
        weights1[43399] <= 16'b0000000000000001;
        weights1[43400] <= 16'b1111111111111111;
        weights1[43401] <= 16'b1111111111111101;
        weights1[43402] <= 16'b1111111111110010;
        weights1[43403] <= 16'b1111111111101111;
        weights1[43404] <= 16'b1111111111111001;
        weights1[43405] <= 16'b0000000000000111;
        weights1[43406] <= 16'b1111111111110111;
        weights1[43407] <= 16'b1111111111111010;
        weights1[43408] <= 16'b1111111111111110;
        weights1[43409] <= 16'b1111111111110111;
        weights1[43410] <= 16'b1111111111101100;
        weights1[43411] <= 16'b0000000000000001;
        weights1[43412] <= 16'b1111111111111010;
        weights1[43413] <= 16'b1111111111100110;
        weights1[43414] <= 16'b1111111111101001;
        weights1[43415] <= 16'b0000000000000100;
        weights1[43416] <= 16'b1111111111101110;
        weights1[43417] <= 16'b0000000000010110;
        weights1[43418] <= 16'b1111111111110001;
        weights1[43419] <= 16'b1111111111110100;
        weights1[43420] <= 16'b1111111111101111;
        weights1[43421] <= 16'b1111111111100110;
        weights1[43422] <= 16'b0000000000001101;
        weights1[43423] <= 16'b1111111111110001;
        weights1[43424] <= 16'b1111111111111010;
        weights1[43425] <= 16'b1111111111111100;
        weights1[43426] <= 16'b1111111111111010;
        weights1[43427] <= 16'b1111111111111111;
        weights1[43428] <= 16'b1111111111111001;
        weights1[43429] <= 16'b1111111111111110;
        weights1[43430] <= 16'b1111111111110010;
        weights1[43431] <= 16'b1111111111110000;
        weights1[43432] <= 16'b0000000000010011;
        weights1[43433] <= 16'b1111111111100110;
        weights1[43434] <= 16'b1111111111101101;
        weights1[43435] <= 16'b1111111111110110;
        weights1[43436] <= 16'b1111111111110001;
        weights1[43437] <= 16'b1111111111110111;
        weights1[43438] <= 16'b1111111111100110;
        weights1[43439] <= 16'b1111111111100111;
        weights1[43440] <= 16'b1111111111100110;
        weights1[43441] <= 16'b1111111111111111;
        weights1[43442] <= 16'b1111111111100011;
        weights1[43443] <= 16'b1111111111101111;
        weights1[43444] <= 16'b1111111111110100;
        weights1[43445] <= 16'b1111111111111000;
        weights1[43446] <= 16'b0000000000001110;
        weights1[43447] <= 16'b1111111111110001;
        weights1[43448] <= 16'b0000000000001000;
        weights1[43449] <= 16'b0000000000001101;
        weights1[43450] <= 16'b0000000000001001;
        weights1[43451] <= 16'b1111111111110010;
        weights1[43452] <= 16'b1111111111101100;
        weights1[43453] <= 16'b0000000000000001;
        weights1[43454] <= 16'b0000000000000010;
        weights1[43455] <= 16'b0000000000000011;
        weights1[43456] <= 16'b1111111111111100;
        weights1[43457] <= 16'b0000000000000011;
        weights1[43458] <= 16'b1111111111111010;
        weights1[43459] <= 16'b0000000000000000;
        weights1[43460] <= 16'b0000000000000000;
        weights1[43461] <= 16'b1111111111100010;
        weights1[43462] <= 16'b1111111111101110;
        weights1[43463] <= 16'b1111111111111001;
        weights1[43464] <= 16'b1111111111100101;
        weights1[43465] <= 16'b1111111111110011;
        weights1[43466] <= 16'b1111111111110011;
        weights1[43467] <= 16'b1111111111110110;
        weights1[43468] <= 16'b1111111111101111;
        weights1[43469] <= 16'b1111111111101001;
        weights1[43470] <= 16'b1111111111100000;
        weights1[43471] <= 16'b1111111111101100;
        weights1[43472] <= 16'b1111111111111001;
        weights1[43473] <= 16'b1111111111101000;
        weights1[43474] <= 16'b1111111111101101;
        weights1[43475] <= 16'b0000000000000100;
        weights1[43476] <= 16'b1111111111110000;
        weights1[43477] <= 16'b1111111111110010;
        weights1[43478] <= 16'b0000000000001011;
        weights1[43479] <= 16'b0000000000001100;
        weights1[43480] <= 16'b0000000000000000;
        weights1[43481] <= 16'b1111111111110110;
        weights1[43482] <= 16'b1111111111101000;
        weights1[43483] <= 16'b1111111111101111;
        weights1[43484] <= 16'b1111111111111011;
        weights1[43485] <= 16'b1111111111111000;
        weights1[43486] <= 16'b1111111111101101;
        weights1[43487] <= 16'b1111111111110010;
        weights1[43488] <= 16'b1111111111111111;
        weights1[43489] <= 16'b1111111111100101;
        weights1[43490] <= 16'b1111111111101000;
        weights1[43491] <= 16'b1111111111110101;
        weights1[43492] <= 16'b1111111111101110;
        weights1[43493] <= 16'b1111111111101000;
        weights1[43494] <= 16'b1111111111100100;
        weights1[43495] <= 16'b1111111111001111;
        weights1[43496] <= 16'b1111111111010000;
        weights1[43497] <= 16'b1111111111001101;
        weights1[43498] <= 16'b1111111111100101;
        weights1[43499] <= 16'b1111111111011000;
        weights1[43500] <= 16'b1111111111001000;
        weights1[43501] <= 16'b1111111111110100;
        weights1[43502] <= 16'b1111111111101101;
        weights1[43503] <= 16'b1111111111110111;
        weights1[43504] <= 16'b1111111111110001;
        weights1[43505] <= 16'b1111111111111001;
        weights1[43506] <= 16'b1111111111111010;
        weights1[43507] <= 16'b1111111111110101;
        weights1[43508] <= 16'b1111111111101101;
        weights1[43509] <= 16'b1111111111111000;
        weights1[43510] <= 16'b0000000000000011;
        weights1[43511] <= 16'b1111111111110110;
        weights1[43512] <= 16'b0000000000000110;
        weights1[43513] <= 16'b1111111111110110;
        weights1[43514] <= 16'b1111111111110000;
        weights1[43515] <= 16'b1111111111101000;
        weights1[43516] <= 16'b1111111111110000;
        weights1[43517] <= 16'b1111111111110010;
        weights1[43518] <= 16'b1111111111110000;
        weights1[43519] <= 16'b1111111111100111;
        weights1[43520] <= 16'b1111111111111111;
        weights1[43521] <= 16'b1111111111000100;
        weights1[43522] <= 16'b1111111111011010;
        weights1[43523] <= 16'b1111111111100011;
        weights1[43524] <= 16'b1111111111011101;
        weights1[43525] <= 16'b1111111111100100;
        weights1[43526] <= 16'b1111111111001001;
        weights1[43527] <= 16'b1111111111000110;
        weights1[43528] <= 16'b1111111111011011;
        weights1[43529] <= 16'b1111111111010111;
        weights1[43530] <= 16'b1111111111001101;
        weights1[43531] <= 16'b1111111110110111;
        weights1[43532] <= 16'b1111111111000101;
        weights1[43533] <= 16'b1111111111011101;
        weights1[43534] <= 16'b1111111111011111;
        weights1[43535] <= 16'b1111111111101100;
        weights1[43536] <= 16'b1111111111011110;
        weights1[43537] <= 16'b1111111111110001;
        weights1[43538] <= 16'b1111111111110100;
        weights1[43539] <= 16'b1111111111110101;
        weights1[43540] <= 16'b0000000000000001;
        weights1[43541] <= 16'b1111111111111000;
        weights1[43542] <= 16'b1111111111111000;
        weights1[43543] <= 16'b1111111111110010;
        weights1[43544] <= 16'b1111111111011110;
        weights1[43545] <= 16'b1111111111101100;
        weights1[43546] <= 16'b1111111111110011;
        weights1[43547] <= 16'b1111111111100111;
        weights1[43548] <= 16'b1111111111001010;
        weights1[43549] <= 16'b1111111110111111;
        weights1[43550] <= 16'b1111111110111111;
        weights1[43551] <= 16'b1111111111001000;
        weights1[43552] <= 16'b1111111110111101;
        weights1[43553] <= 16'b1111111111000111;
        weights1[43554] <= 16'b1111111111010100;
        weights1[43555] <= 16'b1111111110101111;
        weights1[43556] <= 16'b1111111111010000;
        weights1[43557] <= 16'b1111111110110001;
        weights1[43558] <= 16'b1111111110111000;
        weights1[43559] <= 16'b1111111110111100;
        weights1[43560] <= 16'b1111111111000011;
        weights1[43561] <= 16'b1111111111001001;
        weights1[43562] <= 16'b1111111111011110;
        weights1[43563] <= 16'b1111111111001111;
        weights1[43564] <= 16'b1111111111110000;
        weights1[43565] <= 16'b1111111111101010;
        weights1[43566] <= 16'b1111111111101111;
        weights1[43567] <= 16'b1111111111110111;
        weights1[43568] <= 16'b0000000000001001;
        weights1[43569] <= 16'b0000000000000011;
        weights1[43570] <= 16'b0000000000000110;
        weights1[43571] <= 16'b0000000000000000;
        weights1[43572] <= 16'b0000000000000000;
        weights1[43573] <= 16'b1111111111111011;
        weights1[43574] <= 16'b1111111111100101;
        weights1[43575] <= 16'b1111111110111110;
        weights1[43576] <= 16'b1111111111001001;
        weights1[43577] <= 16'b1111111110101011;
        weights1[43578] <= 16'b1111111110110111;
        weights1[43579] <= 16'b1111111110111101;
        weights1[43580] <= 16'b1111111111011100;
        weights1[43581] <= 16'b1111111111001111;
        weights1[43582] <= 16'b1111111111001101;
        weights1[43583] <= 16'b1111111110111110;
        weights1[43584] <= 16'b1111111111100101;
        weights1[43585] <= 16'b1111111110111000;
        weights1[43586] <= 16'b1111111111010010;
        weights1[43587] <= 16'b1111111111000110;
        weights1[43588] <= 16'b1111111111000110;
        weights1[43589] <= 16'b1111111111000011;
        weights1[43590] <= 16'b1111111111001001;
        weights1[43591] <= 16'b1111111111001110;
        weights1[43592] <= 16'b1111111111100101;
        weights1[43593] <= 16'b1111111111101100;
        weights1[43594] <= 16'b1111111111111001;
        weights1[43595] <= 16'b1111111111111111;
        weights1[43596] <= 16'b0000000000000101;
        weights1[43597] <= 16'b0000000000010110;
        weights1[43598] <= 16'b0000000000011100;
        weights1[43599] <= 16'b0000000000010011;
        weights1[43600] <= 16'b0000000000011111;
        weights1[43601] <= 16'b0000000000011110;
        weights1[43602] <= 16'b0000000000010001;
        weights1[43603] <= 16'b0000000000100100;
        weights1[43604] <= 16'b1111111111101110;
        weights1[43605] <= 16'b1111111111101111;
        weights1[43606] <= 16'b1111111111011010;
        weights1[43607] <= 16'b1111111111010001;
        weights1[43608] <= 16'b1111111111101011;
        weights1[43609] <= 16'b1111111111011010;
        weights1[43610] <= 16'b1111111110111000;
        weights1[43611] <= 16'b1111111111010001;
        weights1[43612] <= 16'b1111111110110101;
        weights1[43613] <= 16'b1111111111000011;
        weights1[43614] <= 16'b1111111111001001;
        weights1[43615] <= 16'b1111111111001110;
        weights1[43616] <= 16'b1111111110111001;
        weights1[43617] <= 16'b1111111110111011;
        weights1[43618] <= 16'b1111111111011011;
        weights1[43619] <= 16'b1111111111101001;
        weights1[43620] <= 16'b1111111111100011;
        weights1[43621] <= 16'b1111111111110100;
        weights1[43622] <= 16'b0000000000010010;
        weights1[43623] <= 16'b0000000000010110;
        weights1[43624] <= 16'b0000000000010000;
        weights1[43625] <= 16'b0000000000100011;
        weights1[43626] <= 16'b0000000000101101;
        weights1[43627] <= 16'b0000000000011110;
        weights1[43628] <= 16'b0000000000101001;
        weights1[43629] <= 16'b0000000000110100;
        weights1[43630] <= 16'b0000000000010000;
        weights1[43631] <= 16'b0000000000100101;
        weights1[43632] <= 16'b0000000000100110;
        weights1[43633] <= 16'b0000000000011001;
        weights1[43634] <= 16'b0000000000000010;
        weights1[43635] <= 16'b1111111111110101;
        weights1[43636] <= 16'b1111111111111001;
        weights1[43637] <= 16'b1111111111110011;
        weights1[43638] <= 16'b1111111110111100;
        weights1[43639] <= 16'b1111111111010001;
        weights1[43640] <= 16'b1111111111100101;
        weights1[43641] <= 16'b1111111111001101;
        weights1[43642] <= 16'b1111111111011100;
        weights1[43643] <= 16'b1111111111010111;
        weights1[43644] <= 16'b1111111111100000;
        weights1[43645] <= 16'b1111111111011011;
        weights1[43646] <= 16'b1111111111111010;
        weights1[43647] <= 16'b1111111111110000;
        weights1[43648] <= 16'b1111111111100111;
        weights1[43649] <= 16'b0000000000000101;
        weights1[43650] <= 16'b0000000000011011;
        weights1[43651] <= 16'b0000000000100010;
        weights1[43652] <= 16'b0000000000011011;
        weights1[43653] <= 16'b0000000000101000;
        weights1[43654] <= 16'b0000000000101101;
        weights1[43655] <= 16'b0000000000100111;
        weights1[43656] <= 16'b0000000000101000;
        weights1[43657] <= 16'b0000000000010001;
        weights1[43658] <= 16'b0000000000011111;
        weights1[43659] <= 16'b0000000000101111;
        weights1[43660] <= 16'b0000000000100000;
        weights1[43661] <= 16'b0000000000001000;
        weights1[43662] <= 16'b0000000000001111;
        weights1[43663] <= 16'b0000000000001100;
        weights1[43664] <= 16'b0000000000000101;
        weights1[43665] <= 16'b1111111111111111;
        weights1[43666] <= 16'b1111111111110110;
        weights1[43667] <= 16'b1111111111110001;
        weights1[43668] <= 16'b1111111111100110;
        weights1[43669] <= 16'b1111111111101000;
        weights1[43670] <= 16'b1111111111110011;
        weights1[43671] <= 16'b1111111111111011;
        weights1[43672] <= 16'b0000000000000111;
        weights1[43673] <= 16'b1111111111110101;
        weights1[43674] <= 16'b1111111111110100;
        weights1[43675] <= 16'b1111111111111100;
        weights1[43676] <= 16'b0000000000001111;
        weights1[43677] <= 16'b0000000000100001;
        weights1[43678] <= 16'b0000000000011110;
        weights1[43679] <= 16'b0000000000100011;
        weights1[43680] <= 16'b0000000000011100;
        weights1[43681] <= 16'b0000000000101000;
        weights1[43682] <= 16'b0000000000011011;
        weights1[43683] <= 16'b0000000000110010;
        weights1[43684] <= 16'b0000000000100010;
        weights1[43685] <= 16'b0000000000101111;
        weights1[43686] <= 16'b0000000000101100;
        weights1[43687] <= 16'b0000000000100100;
        weights1[43688] <= 16'b0000000000011010;
        weights1[43689] <= 16'b0000000000111001;
        weights1[43690] <= 16'b0000000001001001;
        weights1[43691] <= 16'b0000000000010110;
        weights1[43692] <= 16'b0000000000111100;
        weights1[43693] <= 16'b0000000000111001;
        weights1[43694] <= 16'b0000000000111101;
        weights1[43695] <= 16'b0000000000011001;
        weights1[43696] <= 16'b0000000000101010;
        weights1[43697] <= 16'b1111111111111111;
        weights1[43698] <= 16'b0000000000101010;
        weights1[43699] <= 16'b0000000000100000;
        weights1[43700] <= 16'b0000000000001001;
        weights1[43701] <= 16'b0000000000010010;
        weights1[43702] <= 16'b0000000000110000;
        weights1[43703] <= 16'b0000000000101010;
        weights1[43704] <= 16'b0000000000101100;
        weights1[43705] <= 16'b0000000000110000;
        weights1[43706] <= 16'b0000000000100100;
        weights1[43707] <= 16'b0000000000100000;
        weights1[43708] <= 16'b0000000000011111;
        weights1[43709] <= 16'b0000000000101001;
        weights1[43710] <= 16'b0000000000101000;
        weights1[43711] <= 16'b0000000000101000;
        weights1[43712] <= 16'b0000000000011100;
        weights1[43713] <= 16'b0000000000100111;
        weights1[43714] <= 16'b0000000001000001;
        weights1[43715] <= 16'b0000000000101000;
        weights1[43716] <= 16'b0000000000100110;
        weights1[43717] <= 16'b0000000000110000;
        weights1[43718] <= 16'b0000000000111010;
        weights1[43719] <= 16'b0000000001010011;
        weights1[43720] <= 16'b0000000000111101;
        weights1[43721] <= 16'b0000000000111110;
        weights1[43722] <= 16'b0000000001011011;
        weights1[43723] <= 16'b0000000001011001;
        weights1[43724] <= 16'b0000000001001001;
        weights1[43725] <= 16'b0000000001001110;
        weights1[43726] <= 16'b0000000001001010;
        weights1[43727] <= 16'b0000000001000101;
        weights1[43728] <= 16'b0000000000111111;
        weights1[43729] <= 16'b0000000000101110;
        weights1[43730] <= 16'b0000000000111000;
        weights1[43731] <= 16'b0000000000111001;
        weights1[43732] <= 16'b0000000000110010;
        weights1[43733] <= 16'b0000000000111001;
        weights1[43734] <= 16'b0000000000101100;
        weights1[43735] <= 16'b0000000000100101;
        weights1[43736] <= 16'b0000000000011011;
        weights1[43737] <= 16'b0000000000100011;
        weights1[43738] <= 16'b0000000000100011;
        weights1[43739] <= 16'b0000000000100011;
        weights1[43740] <= 16'b0000000000100000;
        weights1[43741] <= 16'b0000000000110000;
        weights1[43742] <= 16'b0000000000111101;
        weights1[43743] <= 16'b0000000000100111;
        weights1[43744] <= 16'b0000000000111111;
        weights1[43745] <= 16'b0000000001000101;
        weights1[43746] <= 16'b0000000000011110;
        weights1[43747] <= 16'b0000000001000000;
        weights1[43748] <= 16'b0000000000101111;
        weights1[43749] <= 16'b0000000000110110;
        weights1[43750] <= 16'b0000000000110100;
        weights1[43751] <= 16'b0000000001000010;
        weights1[43752] <= 16'b0000000000110011;
        weights1[43753] <= 16'b0000000001000011;
        weights1[43754] <= 16'b0000000000011001;
        weights1[43755] <= 16'b0000000000011010;
        weights1[43756] <= 16'b0000000001001100;
        weights1[43757] <= 16'b0000000000101110;
        weights1[43758] <= 16'b0000000000111010;
        weights1[43759] <= 16'b0000000000101101;
        weights1[43760] <= 16'b0000000000111001;
        weights1[43761] <= 16'b0000000000111100;
        weights1[43762] <= 16'b0000000000101101;
        weights1[43763] <= 16'b0000000000011100;
        weights1[43764] <= 16'b0000000000011010;
        weights1[43765] <= 16'b0000000000011101;
        weights1[43766] <= 16'b0000000000101110;
        weights1[43767] <= 16'b0000000000001101;
        weights1[43768] <= 16'b0000000000101000;
        weights1[43769] <= 16'b0000000000100111;
        weights1[43770] <= 16'b0000000000010111;
        weights1[43771] <= 16'b0000000000101001;
        weights1[43772] <= 16'b0000000000100110;
        weights1[43773] <= 16'b0000000000110101;
        weights1[43774] <= 16'b0000000000100000;
        weights1[43775] <= 16'b0000000000110101;
        weights1[43776] <= 16'b0000000000111100;
        weights1[43777] <= 16'b0000000000101110;
        weights1[43778] <= 16'b0000000000100000;
        weights1[43779] <= 16'b0000000001001101;
        weights1[43780] <= 16'b0000000001000011;
        weights1[43781] <= 16'b0000000000111001;
        weights1[43782] <= 16'b0000000000101000;
        weights1[43783] <= 16'b0000000001001011;
        weights1[43784] <= 16'b0000000000111100;
        weights1[43785] <= 16'b0000000000101110;
        weights1[43786] <= 16'b0000000000101111;
        weights1[43787] <= 16'b0000000000101111;
        weights1[43788] <= 16'b0000000000110010;
        weights1[43789] <= 16'b0000000000111010;
        weights1[43790] <= 16'b0000000000101001;
        weights1[43791] <= 16'b0000000000011001;
        weights1[43792] <= 16'b0000000000010001;
        weights1[43793] <= 16'b0000000000001110;
        weights1[43794] <= 16'b0000000000011000;
        weights1[43795] <= 16'b0000000000010011;
        weights1[43796] <= 16'b0000000000010100;
        weights1[43797] <= 16'b0000000000001010;
        weights1[43798] <= 16'b0000000000100100;
        weights1[43799] <= 16'b0000000000110000;
        weights1[43800] <= 16'b0000000000010001;
        weights1[43801] <= 16'b0000000000001110;
        weights1[43802] <= 16'b0000000000001010;
        weights1[43803] <= 16'b0000000000100110;
        weights1[43804] <= 16'b0000000000100001;
        weights1[43805] <= 16'b0000000000111110;
        weights1[43806] <= 16'b0000000001000010;
        weights1[43807] <= 16'b0000000000101001;
        weights1[43808] <= 16'b0000000000101011;
        weights1[43809] <= 16'b0000000001000101;
        weights1[43810] <= 16'b0000000001000000;
        weights1[43811] <= 16'b0000000000110100;
        weights1[43812] <= 16'b0000000000110100;
        weights1[43813] <= 16'b0000000001000011;
        weights1[43814] <= 16'b0000000000110011;
        weights1[43815] <= 16'b0000000000101110;
        weights1[43816] <= 16'b0000000000101111;
        weights1[43817] <= 16'b0000000000100010;
        weights1[43818] <= 16'b0000000000100000;
        weights1[43819] <= 16'b0000000000010010;
        weights1[43820] <= 16'b0000000000000100;
        weights1[43821] <= 16'b0000000000001011;
        weights1[43822] <= 16'b0000000000001111;
        weights1[43823] <= 16'b0000000000001100;
        weights1[43824] <= 16'b0000000000011001;
        weights1[43825] <= 16'b0000000000000011;
        weights1[43826] <= 16'b0000000000010011;
        weights1[43827] <= 16'b1111111111110110;
        weights1[43828] <= 16'b0000000000100010;
        weights1[43829] <= 16'b0000000000010001;
        weights1[43830] <= 16'b0000000000011101;
        weights1[43831] <= 16'b0000000000100100;
        weights1[43832] <= 16'b0000000000010100;
        weights1[43833] <= 16'b0000000000011011;
        weights1[43834] <= 16'b0000000000001101;
        weights1[43835] <= 16'b0000000000100000;
        weights1[43836] <= 16'b0000000000101001;
        weights1[43837] <= 16'b0000000000111010;
        weights1[43838] <= 16'b0000000000110011;
        weights1[43839] <= 16'b0000000001001011;
        weights1[43840] <= 16'b0000000000101011;
        weights1[43841] <= 16'b0000000000011000;
        weights1[43842] <= 16'b0000000000101010;
        weights1[43843] <= 16'b0000000000110010;
        weights1[43844] <= 16'b0000000000100011;
        weights1[43845] <= 16'b0000000000100001;
        weights1[43846] <= 16'b0000000000010110;
        weights1[43847] <= 16'b0000000000000110;
        weights1[43848] <= 16'b0000000000000011;
        weights1[43849] <= 16'b0000000000000111;
        weights1[43850] <= 16'b1111111111111111;
        weights1[43851] <= 16'b0000000000000010;
        weights1[43852] <= 16'b0000000000010110;
        weights1[43853] <= 16'b0000000000000111;
        weights1[43854] <= 16'b0000000000000110;
        weights1[43855] <= 16'b0000000000000100;
        weights1[43856] <= 16'b0000000000010011;
        weights1[43857] <= 16'b0000000000001001;
        weights1[43858] <= 16'b0000000000010101;
        weights1[43859] <= 16'b0000000000011011;
        weights1[43860] <= 16'b0000000000001100;
        weights1[43861] <= 16'b1111111111111011;
        weights1[43862] <= 16'b0000000000001110;
        weights1[43863] <= 16'b0000000000001101;
        weights1[43864] <= 16'b0000000000000011;
        weights1[43865] <= 16'b1111111111110110;
        weights1[43866] <= 16'b1111111111111110;
        weights1[43867] <= 16'b0000000000001111;
        weights1[43868] <= 16'b0000000000001010;
        weights1[43869] <= 16'b0000000000100001;
        weights1[43870] <= 16'b0000000000100000;
        weights1[43871] <= 16'b0000000000011001;
        weights1[43872] <= 16'b0000000000001111;
        weights1[43873] <= 16'b0000000000000001;
        weights1[43874] <= 16'b0000000000000111;
        weights1[43875] <= 16'b0000000000000001;
        weights1[43876] <= 16'b1111111111111101;
        weights1[43877] <= 16'b1111111111111010;
        weights1[43878] <= 16'b0000000000000010;
        weights1[43879] <= 16'b0000000000000111;
        weights1[43880] <= 16'b0000000000001001;
        weights1[43881] <= 16'b1111111111111101;
        weights1[43882] <= 16'b0000000000010000;
        weights1[43883] <= 16'b0000000000001000;
        weights1[43884] <= 16'b1111111111111110;
        weights1[43885] <= 16'b1111111111101011;
        weights1[43886] <= 16'b1111111111110101;
        weights1[43887] <= 16'b1111111111110101;
        weights1[43888] <= 16'b1111111111110001;
        weights1[43889] <= 16'b1111111111100110;
        weights1[43890] <= 16'b1111111111101101;
        weights1[43891] <= 16'b1111111111110110;
        weights1[43892] <= 16'b1111111111111111;
        weights1[43893] <= 16'b0000000000000100;
        weights1[43894] <= 16'b0000000000001110;
        weights1[43895] <= 16'b0000000000000110;
        weights1[43896] <= 16'b1111111111101101;
        weights1[43897] <= 16'b0000000000001010;
        weights1[43898] <= 16'b0000000000011011;
        weights1[43899] <= 16'b0000000000001000;
        weights1[43900] <= 16'b0000000000000110;
        weights1[43901] <= 16'b0000000000000010;
        weights1[43902] <= 16'b0000000000000001;
        weights1[43903] <= 16'b0000000000000000;
        weights1[43904] <= 16'b0000000000000000;
        weights1[43905] <= 16'b1111111111111111;
        weights1[43906] <= 16'b1111111111111011;
        weights1[43907] <= 16'b1111111111110101;
        weights1[43908] <= 16'b1111111111110010;
        weights1[43909] <= 16'b1111111111110001;
        weights1[43910] <= 16'b1111111111101110;
        weights1[43911] <= 16'b1111111111100111;
        weights1[43912] <= 16'b1111111111100100;
        weights1[43913] <= 16'b1111111111100101;
        weights1[43914] <= 16'b1111111111101000;
        weights1[43915] <= 16'b1111111111101100;
        weights1[43916] <= 16'b1111111111101111;
        weights1[43917] <= 16'b1111111111110111;
        weights1[43918] <= 16'b1111111111111010;
        weights1[43919] <= 16'b1111111111110100;
        weights1[43920] <= 16'b1111111111110010;
        weights1[43921] <= 16'b1111111111101010;
        weights1[43922] <= 16'b1111111111110001;
        weights1[43923] <= 16'b1111111111101011;
        weights1[43924] <= 16'b1111111111110011;
        weights1[43925] <= 16'b1111111111111000;
        weights1[43926] <= 16'b0000000000000011;
        weights1[43927] <= 16'b1111111111111010;
        weights1[43928] <= 16'b0000000000000101;
        weights1[43929] <= 16'b1111111111111110;
        weights1[43930] <= 16'b0000000000000001;
        weights1[43931] <= 16'b1111111111111100;
        weights1[43932] <= 16'b0000000000000000;
        weights1[43933] <= 16'b1111111111111101;
        weights1[43934] <= 16'b1111111111110101;
        weights1[43935] <= 16'b1111111111101110;
        weights1[43936] <= 16'b1111111111101100;
        weights1[43937] <= 16'b1111111111101010;
        weights1[43938] <= 16'b1111111111100010;
        weights1[43939] <= 16'b1111111111011100;
        weights1[43940] <= 16'b1111111111100001;
        weights1[43941] <= 16'b1111111111011000;
        weights1[43942] <= 16'b1111111111011000;
        weights1[43943] <= 16'b1111111111011000;
        weights1[43944] <= 16'b1111111111100010;
        weights1[43945] <= 16'b1111111111100011;
        weights1[43946] <= 16'b1111111111101000;
        weights1[43947] <= 16'b1111111111011100;
        weights1[43948] <= 16'b1111111111010011;
        weights1[43949] <= 16'b1111111111011110;
        weights1[43950] <= 16'b1111111111100100;
        weights1[43951] <= 16'b1111111111100110;
        weights1[43952] <= 16'b1111111111101010;
        weights1[43953] <= 16'b1111111111110010;
        weights1[43954] <= 16'b1111111111101011;
        weights1[43955] <= 16'b1111111111110010;
        weights1[43956] <= 16'b1111111111111101;
        weights1[43957] <= 16'b0000000000000011;
        weights1[43958] <= 16'b1111111111111001;
        weights1[43959] <= 16'b1111111111110110;
        weights1[43960] <= 16'b1111111111111101;
        weights1[43961] <= 16'b1111111111111001;
        weights1[43962] <= 16'b1111111111110010;
        weights1[43963] <= 16'b1111111111101001;
        weights1[43964] <= 16'b1111111111100100;
        weights1[43965] <= 16'b1111111111011111;
        weights1[43966] <= 16'b1111111111011001;
        weights1[43967] <= 16'b1111111111010000;
        weights1[43968] <= 16'b1111111111001100;
        weights1[43969] <= 16'b1111111111000100;
        weights1[43970] <= 16'b1111111111001000;
        weights1[43971] <= 16'b1111111111001000;
        weights1[43972] <= 16'b1111111111001011;
        weights1[43973] <= 16'b1111111111000010;
        weights1[43974] <= 16'b1111111110110110;
        weights1[43975] <= 16'b1111111110111110;
        weights1[43976] <= 16'b1111111111000100;
        weights1[43977] <= 16'b1111111111001111;
        weights1[43978] <= 16'b1111111111001011;
        weights1[43979] <= 16'b1111111111001001;
        weights1[43980] <= 16'b1111111111011001;
        weights1[43981] <= 16'b1111111111011100;
        weights1[43982] <= 16'b1111111111100000;
        weights1[43983] <= 16'b1111111111110011;
        weights1[43984] <= 16'b1111111111101001;
        weights1[43985] <= 16'b1111111111101001;
        weights1[43986] <= 16'b1111111111110010;
        weights1[43987] <= 16'b1111111111110000;
        weights1[43988] <= 16'b1111111111111101;
        weights1[43989] <= 16'b1111111111110010;
        weights1[43990] <= 16'b1111111111101100;
        weights1[43991] <= 16'b1111111111100010;
        weights1[43992] <= 16'b1111111111011110;
        weights1[43993] <= 16'b1111111111010111;
        weights1[43994] <= 16'b1111111111001100;
        weights1[43995] <= 16'b1111111111000011;
        weights1[43996] <= 16'b1111111111000010;
        weights1[43997] <= 16'b1111111110111100;
        weights1[43998] <= 16'b1111111110110001;
        weights1[43999] <= 16'b1111111110101101;
        weights1[44000] <= 16'b1111111110101100;
        weights1[44001] <= 16'b1111111110111001;
        weights1[44002] <= 16'b1111111111001110;
        weights1[44003] <= 16'b1111111110111010;
        weights1[44004] <= 16'b1111111111001110;
        weights1[44005] <= 16'b1111111111010100;
        weights1[44006] <= 16'b1111111111100000;
        weights1[44007] <= 16'b1111111111001101;
        weights1[44008] <= 16'b1111111111001110;
        weights1[44009] <= 16'b1111111111010101;
        weights1[44010] <= 16'b1111111111010000;
        weights1[44011] <= 16'b1111111111100011;
        weights1[44012] <= 16'b1111111111101110;
        weights1[44013] <= 16'b1111111111101110;
        weights1[44014] <= 16'b1111111111111010;
        weights1[44015] <= 16'b0000000000000011;
        weights1[44016] <= 16'b1111111111111001;
        weights1[44017] <= 16'b1111111111110000;
        weights1[44018] <= 16'b1111111111101010;
        weights1[44019] <= 16'b1111111111100110;
        weights1[44020] <= 16'b1111111111100011;
        weights1[44021] <= 16'b1111111111010000;
        weights1[44022] <= 16'b1111111111000010;
        weights1[44023] <= 16'b1111111110110010;
        weights1[44024] <= 16'b1111111111000000;
        weights1[44025] <= 16'b1111111111000010;
        weights1[44026] <= 16'b1111111111000110;
        weights1[44027] <= 16'b1111111111001010;
        weights1[44028] <= 16'b1111111111011000;
        weights1[44029] <= 16'b1111111111001010;
        weights1[44030] <= 16'b1111111111110101;
        weights1[44031] <= 16'b1111111111101011;
        weights1[44032] <= 16'b1111111111111001;
        weights1[44033] <= 16'b1111111111011000;
        weights1[44034] <= 16'b1111111111100100;
        weights1[44035] <= 16'b1111111111101001;
        weights1[44036] <= 16'b1111111111001110;
        weights1[44037] <= 16'b1111111111010111;
        weights1[44038] <= 16'b1111111111010001;
        weights1[44039] <= 16'b0000000000001010;
        weights1[44040] <= 16'b1111111111111000;
        weights1[44041] <= 16'b1111111111110101;
        weights1[44042] <= 16'b0000000000000110;
        weights1[44043] <= 16'b0000000000001001;
        weights1[44044] <= 16'b1111111111111100;
        weights1[44045] <= 16'b1111111111110010;
        weights1[44046] <= 16'b1111111111100110;
        weights1[44047] <= 16'b1111111111101001;
        weights1[44048] <= 16'b1111111111100111;
        weights1[44049] <= 16'b1111111111110010;
        weights1[44050] <= 16'b1111111111011011;
        weights1[44051] <= 16'b1111111111110110;
        weights1[44052] <= 16'b1111111111111001;
        weights1[44053] <= 16'b0000000000000001;
        weights1[44054] <= 16'b0000000000001100;
        weights1[44055] <= 16'b0000000000010101;
        weights1[44056] <= 16'b1111111111111110;
        weights1[44057] <= 16'b1111111111110011;
        weights1[44058] <= 16'b1111111111110000;
        weights1[44059] <= 16'b1111111111111101;
        weights1[44060] <= 16'b1111111111110100;
        weights1[44061] <= 16'b0000000000000111;
        weights1[44062] <= 16'b1111111111111000;
        weights1[44063] <= 16'b1111111111111101;
        weights1[44064] <= 16'b1111111111111111;
        weights1[44065] <= 16'b1111111111100110;
        weights1[44066] <= 16'b1111111111110011;
        weights1[44067] <= 16'b1111111111110001;
        weights1[44068] <= 16'b1111111111100000;
        weights1[44069] <= 16'b1111111111110011;
        weights1[44070] <= 16'b0000000000001101;
        weights1[44071] <= 16'b0000000000010101;
        weights1[44072] <= 16'b1111111111111100;
        weights1[44073] <= 16'b1111111111111000;
        weights1[44074] <= 16'b1111111111111001;
        weights1[44075] <= 16'b1111111111111000;
        weights1[44076] <= 16'b0000000000000100;
        weights1[44077] <= 16'b1111111111100100;
        weights1[44078] <= 16'b1111111111111110;
        weights1[44079] <= 16'b0000000000001111;
        weights1[44080] <= 16'b0000000000011110;
        weights1[44081] <= 16'b0000000000000100;
        weights1[44082] <= 16'b1111111111110011;
        weights1[44083] <= 16'b1111111111110111;
        weights1[44084] <= 16'b0000000000001111;
        weights1[44085] <= 16'b0000000000001001;
        weights1[44086] <= 16'b0000000000010000;
        weights1[44087] <= 16'b1111111111111111;
        weights1[44088] <= 16'b1111111111110001;
        weights1[44089] <= 16'b0000000000000001;
        weights1[44090] <= 16'b1111111111111011;
        weights1[44091] <= 16'b1111111111110110;
        weights1[44092] <= 16'b0000000000000110;
        weights1[44093] <= 16'b0000000000011001;
        weights1[44094] <= 16'b1111111111111101;
        weights1[44095] <= 16'b1111111111111001;
        weights1[44096] <= 16'b1111111111101101;
        weights1[44097] <= 16'b0000000000000111;
        weights1[44098] <= 16'b0000000000000011;
        weights1[44099] <= 16'b0000000000001000;
        weights1[44100] <= 16'b1111111111111110;
        weights1[44101] <= 16'b0000000000000000;
        weights1[44102] <= 16'b1111111111111101;
        weights1[44103] <= 16'b0000000000000100;
        weights1[44104] <= 16'b0000000000000100;
        weights1[44105] <= 16'b0000000000000101;
        weights1[44106] <= 16'b0000000000000010;
        weights1[44107] <= 16'b1111111111110001;
        weights1[44108] <= 16'b1111111111111101;
        weights1[44109] <= 16'b1111111111101011;
        weights1[44110] <= 16'b0000000000010001;
        weights1[44111] <= 16'b1111111111110111;
        weights1[44112] <= 16'b0000000000001011;
        weights1[44113] <= 16'b0000000000001110;
        weights1[44114] <= 16'b0000000000000101;
        weights1[44115] <= 16'b0000000000001100;
        weights1[44116] <= 16'b0000000000000111;
        weights1[44117] <= 16'b0000000000001001;
        weights1[44118] <= 16'b0000000000001101;
        weights1[44119] <= 16'b0000000000000001;
        weights1[44120] <= 16'b1111111111111110;
        weights1[44121] <= 16'b1111111111101110;
        weights1[44122] <= 16'b1111111111111010;
        weights1[44123] <= 16'b1111111111111011;
        weights1[44124] <= 16'b0000000000000001;
        weights1[44125] <= 16'b1111111111110101;
        weights1[44126] <= 16'b0000000000000011;
        weights1[44127] <= 16'b0000000000000101;
        weights1[44128] <= 16'b1111111111111100;
        weights1[44129] <= 16'b0000000000000110;
        weights1[44130] <= 16'b0000000000000000;
        weights1[44131] <= 16'b0000000000001000;
        weights1[44132] <= 16'b0000000000000010;
        weights1[44133] <= 16'b0000000000001110;
        weights1[44134] <= 16'b0000000000010101;
        weights1[44135] <= 16'b0000000000000010;
        weights1[44136] <= 16'b1111111111110011;
        weights1[44137] <= 16'b0000000000001111;
        weights1[44138] <= 16'b1111111111110010;
        weights1[44139] <= 16'b0000000000000001;
        weights1[44140] <= 16'b1111111111101110;
        weights1[44141] <= 16'b0000000000000001;
        weights1[44142] <= 16'b1111111111111110;
        weights1[44143] <= 16'b1111111111110100;
        weights1[44144] <= 16'b1111111111111111;
        weights1[44145] <= 16'b1111111111110111;
        weights1[44146] <= 16'b0000000000000011;
        weights1[44147] <= 16'b1111111111111110;
        weights1[44148] <= 16'b1111111111111000;
        weights1[44149] <= 16'b1111111111110010;
        weights1[44150] <= 16'b1111111111111100;
        weights1[44151] <= 16'b0000000000001000;
        weights1[44152] <= 16'b1111111111110100;
        weights1[44153] <= 16'b0000000000001010;
        weights1[44154] <= 16'b1111111111111110;
        weights1[44155] <= 16'b0000000000001010;
        weights1[44156] <= 16'b0000000000000111;
        weights1[44157] <= 16'b0000000000001110;
        weights1[44158] <= 16'b0000000000000101;
        weights1[44159] <= 16'b1111111111111111;
        weights1[44160] <= 16'b0000000000000111;
        weights1[44161] <= 16'b1111111111110010;
        weights1[44162] <= 16'b0000000000010010;
        weights1[44163] <= 16'b0000000000000001;
        weights1[44164] <= 16'b1111111111110101;
        weights1[44165] <= 16'b0000000000000101;
        weights1[44166] <= 16'b0000000000000010;
        weights1[44167] <= 16'b0000000000001011;
        weights1[44168] <= 16'b0000000000010001;
        weights1[44169] <= 16'b1111111111111011;
        weights1[44170] <= 16'b0000000000000010;
        weights1[44171] <= 16'b0000000000000101;
        weights1[44172] <= 16'b0000000000000000;
        weights1[44173] <= 16'b0000000000001011;
        weights1[44174] <= 16'b1111111111111001;
        weights1[44175] <= 16'b1111111111111100;
        weights1[44176] <= 16'b0000000000010010;
        weights1[44177] <= 16'b1111111111111110;
        weights1[44178] <= 16'b1111111111111110;
        weights1[44179] <= 16'b1111111111101101;
        weights1[44180] <= 16'b0000000000000011;
        weights1[44181] <= 16'b0000000000000101;
        weights1[44182] <= 16'b1111111111111010;
        weights1[44183] <= 16'b0000000000001001;
        weights1[44184] <= 16'b0000000000010110;
        weights1[44185] <= 16'b0000000000010011;
        weights1[44186] <= 16'b1111111111111110;
        weights1[44187] <= 16'b0000000000010100;
        weights1[44188] <= 16'b0000000000000110;
        weights1[44189] <= 16'b1111111111110001;
        weights1[44190] <= 16'b0000000000001001;
        weights1[44191] <= 16'b1111111111111001;
        weights1[44192] <= 16'b1111111111111001;
        weights1[44193] <= 16'b0000000000001111;
        weights1[44194] <= 16'b0000000000001000;
        weights1[44195] <= 16'b0000000000010001;
        weights1[44196] <= 16'b1111111111111011;
        weights1[44197] <= 16'b0000000000000011;
        weights1[44198] <= 16'b1111111111110111;
        weights1[44199] <= 16'b1111111111110111;
        weights1[44200] <= 16'b1111111111110101;
        weights1[44201] <= 16'b1111111111111111;
        weights1[44202] <= 16'b0000000000000010;
        weights1[44203] <= 16'b1111111111111011;
        weights1[44204] <= 16'b1111111111110011;
        weights1[44205] <= 16'b0000000000000001;
        weights1[44206] <= 16'b1111111111111100;
        weights1[44207] <= 16'b1111111111111111;
        weights1[44208] <= 16'b1111111111101000;
        weights1[44209] <= 16'b1111111111111101;
        weights1[44210] <= 16'b1111111111111001;
        weights1[44211] <= 16'b0000000000000000;
        weights1[44212] <= 16'b0000000000001000;
        weights1[44213] <= 16'b0000000000010010;
        weights1[44214] <= 16'b0000000000000001;
        weights1[44215] <= 16'b1111111111111101;
        weights1[44216] <= 16'b1111111111101100;
        weights1[44217] <= 16'b1111111111111110;
        weights1[44218] <= 16'b1111111111111000;
        weights1[44219] <= 16'b1111111111111011;
        weights1[44220] <= 16'b0000000000010001;
        weights1[44221] <= 16'b0000000000010010;
        weights1[44222] <= 16'b0000000000001000;
        weights1[44223] <= 16'b0000000000001110;
        weights1[44224] <= 16'b0000000000000000;
        weights1[44225] <= 16'b1111111111111010;
        weights1[44226] <= 16'b0000000000000111;
        weights1[44227] <= 16'b1111111111110000;
        weights1[44228] <= 16'b0000000000000110;
        weights1[44229] <= 16'b1111111111111101;
        weights1[44230] <= 16'b0000000000010010;
        weights1[44231] <= 16'b0000000000000101;
        weights1[44232] <= 16'b0000000000000100;
        weights1[44233] <= 16'b1111111111111011;
        weights1[44234] <= 16'b1111111111110101;
        weights1[44235] <= 16'b1111111111111111;
        weights1[44236] <= 16'b0000000000000010;
        weights1[44237] <= 16'b1111111111111001;
        weights1[44238] <= 16'b1111111111111001;
        weights1[44239] <= 16'b0000000000001110;
        weights1[44240] <= 16'b0000000000000000;
        weights1[44241] <= 16'b0000000000000100;
        weights1[44242] <= 16'b0000000000000100;
        weights1[44243] <= 16'b1111111111110010;
        weights1[44244] <= 16'b1111111111111110;
        weights1[44245] <= 16'b1111111111111100;
        weights1[44246] <= 16'b1111111111111011;
        weights1[44247] <= 16'b0000000000000001;
        weights1[44248] <= 16'b1111111111110000;
        weights1[44249] <= 16'b1111111111100001;
        weights1[44250] <= 16'b1111111111101100;
        weights1[44251] <= 16'b1111111111101101;
        weights1[44252] <= 16'b0000000000000101;
        weights1[44253] <= 16'b1111111111110101;
        weights1[44254] <= 16'b1111111111111000;
        weights1[44255] <= 16'b1111111111110111;
        weights1[44256] <= 16'b0000000000000000;
        weights1[44257] <= 16'b1111111111110010;
        weights1[44258] <= 16'b1111111111110011;
        weights1[44259] <= 16'b0000000000000001;
        weights1[44260] <= 16'b1111111111111110;
        weights1[44261] <= 16'b1111111111111011;
        weights1[44262] <= 16'b1111111111111010;
        weights1[44263] <= 16'b0000000000011000;
        weights1[44264] <= 16'b0000000000001100;
        weights1[44265] <= 16'b1111111111111111;
        weights1[44266] <= 16'b0000000000001110;
        weights1[44267] <= 16'b0000000000000011;
        weights1[44268] <= 16'b0000000000000011;
        weights1[44269] <= 16'b0000000000001000;
        weights1[44270] <= 16'b1111111111100100;
        weights1[44271] <= 16'b1111111111101111;
        weights1[44272] <= 16'b0000000000000100;
        weights1[44273] <= 16'b1111111111110111;
        weights1[44274] <= 16'b0000000000000100;
        weights1[44275] <= 16'b0000000000001110;
        weights1[44276] <= 16'b1111111111111100;
        weights1[44277] <= 16'b1111111111111111;
        weights1[44278] <= 16'b0000000000001110;
        weights1[44279] <= 16'b1111111111111001;
        weights1[44280] <= 16'b1111111111110010;
        weights1[44281] <= 16'b0000000000001001;
        weights1[44282] <= 16'b0000000000000100;
        weights1[44283] <= 16'b0000000000000000;
        weights1[44284] <= 16'b1111111111111000;
        weights1[44285] <= 16'b0000000000000101;
        weights1[44286] <= 16'b0000000000000110;
        weights1[44287] <= 16'b0000000000000000;
        weights1[44288] <= 16'b0000000000000001;
        weights1[44289] <= 16'b0000000000000011;
        weights1[44290] <= 16'b1111111111111111;
        weights1[44291] <= 16'b1111111111111100;
        weights1[44292] <= 16'b1111111111111110;
        weights1[44293] <= 16'b0000000000000001;
        weights1[44294] <= 16'b0000000000001011;
        weights1[44295] <= 16'b0000000000001011;
        weights1[44296] <= 16'b1111111111111110;
        weights1[44297] <= 16'b1111111111111011;
        weights1[44298] <= 16'b1111111111110010;
        weights1[44299] <= 16'b1111111111111011;
        weights1[44300] <= 16'b0000000000010101;
        weights1[44301] <= 16'b1111111111110001;
        weights1[44302] <= 16'b1111111111101111;
        weights1[44303] <= 16'b0000000000000000;
        weights1[44304] <= 16'b0000000000000001;
        weights1[44305] <= 16'b0000000000001101;
        weights1[44306] <= 16'b0000000000001100;
        weights1[44307] <= 16'b1111111111111001;
        weights1[44308] <= 16'b1111111111110111;
        weights1[44309] <= 16'b0000000000001101;
        weights1[44310] <= 16'b0000000000010100;
        weights1[44311] <= 16'b0000000000001111;
        weights1[44312] <= 16'b0000000000000111;
        weights1[44313] <= 16'b0000000000001011;
        weights1[44314] <= 16'b1111111111101110;
        weights1[44315] <= 16'b0000000000000101;
        weights1[44316] <= 16'b0000000000000001;
        weights1[44317] <= 16'b0000000000000010;
        weights1[44318] <= 16'b0000000000000100;
        weights1[44319] <= 16'b1111111111110100;
        weights1[44320] <= 16'b0000000000000111;
        weights1[44321] <= 16'b0000000000000100;
        weights1[44322] <= 16'b1111111111111101;
        weights1[44323] <= 16'b0000000000001111;
        weights1[44324] <= 16'b1111111111110001;
        weights1[44325] <= 16'b1111111111101111;
        weights1[44326] <= 16'b1111111111101010;
        weights1[44327] <= 16'b1111111111111101;
        weights1[44328] <= 16'b0000000000000010;
        weights1[44329] <= 16'b0000000000011011;
        weights1[44330] <= 16'b0000000000010101;
        weights1[44331] <= 16'b0000000000000010;
        weights1[44332] <= 16'b0000000000001111;
        weights1[44333] <= 16'b0000000000001100;
        weights1[44334] <= 16'b0000000000010011;
        weights1[44335] <= 16'b0000000000010010;
        weights1[44336] <= 16'b0000000000011101;
        weights1[44337] <= 16'b0000000000001100;
        weights1[44338] <= 16'b0000000000000111;
        weights1[44339] <= 16'b1111111111111001;
        weights1[44340] <= 16'b0000000000010001;
        weights1[44341] <= 16'b0000000000000010;
        weights1[44342] <= 16'b1111111111110110;
        weights1[44343] <= 16'b1111111111111110;
        weights1[44344] <= 16'b1111111111111010;
        weights1[44345] <= 16'b1111111111111110;
        weights1[44346] <= 16'b1111111111101010;
        weights1[44347] <= 16'b1111111111111011;
        weights1[44348] <= 16'b1111111111110100;
        weights1[44349] <= 16'b0000000000000000;
        weights1[44350] <= 16'b1111111111111100;
        weights1[44351] <= 16'b1111111111111100;
        weights1[44352] <= 16'b1111111111101000;
        weights1[44353] <= 16'b1111111111100001;
        weights1[44354] <= 16'b1111111111100001;
        weights1[44355] <= 16'b1111111111010101;
        weights1[44356] <= 16'b0000000000000100;
        weights1[44357] <= 16'b0000000000100101;
        weights1[44358] <= 16'b0000000000100000;
        weights1[44359] <= 16'b0000000000100110;
        weights1[44360] <= 16'b0000000000101011;
        weights1[44361] <= 16'b0000000000011011;
        weights1[44362] <= 16'b0000000000100101;
        weights1[44363] <= 16'b0000000000010101;
        weights1[44364] <= 16'b0000000000010011;
        weights1[44365] <= 16'b0000000000001101;
        weights1[44366] <= 16'b0000000000000011;
        weights1[44367] <= 16'b0000000000001111;
        weights1[44368] <= 16'b0000000000000100;
        weights1[44369] <= 16'b0000000000001010;
        weights1[44370] <= 16'b0000000000001001;
        weights1[44371] <= 16'b0000000000000110;
        weights1[44372] <= 16'b1111111111110100;
        weights1[44373] <= 16'b0000000000000001;
        weights1[44374] <= 16'b0000000000000100;
        weights1[44375] <= 16'b0000000000000111;
        weights1[44376] <= 16'b1111111111111001;
        weights1[44377] <= 16'b1111111111111101;
        weights1[44378] <= 16'b1111111111111011;
        weights1[44379] <= 16'b0000000000000010;
        weights1[44380] <= 16'b1111111111100000;
        weights1[44381] <= 16'b1111111111010010;
        weights1[44382] <= 16'b1111111111000001;
        weights1[44383] <= 16'b1111111111000000;
        weights1[44384] <= 16'b1111111111000101;
        weights1[44385] <= 16'b1111111111111111;
        weights1[44386] <= 16'b0000000000010011;
        weights1[44387] <= 16'b0000000000010110;
        weights1[44388] <= 16'b0000000000010101;
        weights1[44389] <= 16'b0000000000011101;
        weights1[44390] <= 16'b0000000000101001;
        weights1[44391] <= 16'b0000000000010110;
        weights1[44392] <= 16'b0000000000001100;
        weights1[44393] <= 16'b0000000000001001;
        weights1[44394] <= 16'b1111111111111101;
        weights1[44395] <= 16'b0000000000011010;
        weights1[44396] <= 16'b0000000000001111;
        weights1[44397] <= 16'b0000000000000100;
        weights1[44398] <= 16'b0000000000001000;
        weights1[44399] <= 16'b0000000000010001;
        weights1[44400] <= 16'b0000000000001001;
        weights1[44401] <= 16'b0000000000001100;
        weights1[44402] <= 16'b0000000000001011;
        weights1[44403] <= 16'b0000000000010100;
        weights1[44404] <= 16'b0000000000000111;
        weights1[44405] <= 16'b1111111111111001;
        weights1[44406] <= 16'b1111111111111100;
        weights1[44407] <= 16'b1111111111111001;
        weights1[44408] <= 16'b1111111111011011;
        weights1[44409] <= 16'b1111111111000000;
        weights1[44410] <= 16'b1111111110110101;
        weights1[44411] <= 16'b1111111110010101;
        weights1[44412] <= 16'b1111111101110110;
        weights1[44413] <= 16'b1111111111001011;
        weights1[44414] <= 16'b1111111111011011;
        weights1[44415] <= 16'b1111111111100111;
        weights1[44416] <= 16'b0000000000010011;
        weights1[44417] <= 16'b0000000000011000;
        weights1[44418] <= 16'b0000000000011100;
        weights1[44419] <= 16'b0000000000100111;
        weights1[44420] <= 16'b0000000000010011;
        weights1[44421] <= 16'b0000000000011000;
        weights1[44422] <= 16'b0000000000000111;
        weights1[44423] <= 16'b1111111111111110;
        weights1[44424] <= 16'b0000000000001101;
        weights1[44425] <= 16'b0000000000000110;
        weights1[44426] <= 16'b1111111111111110;
        weights1[44427] <= 16'b0000000000000100;
        weights1[44428] <= 16'b0000000000011000;
        weights1[44429] <= 16'b0000000000001000;
        weights1[44430] <= 16'b1111111111111001;
        weights1[44431] <= 16'b0000000000000010;
        weights1[44432] <= 16'b1111111111110010;
        weights1[44433] <= 16'b0000000000011000;
        weights1[44434] <= 16'b0000000000000010;
        weights1[44435] <= 16'b1111111111111111;
        weights1[44436] <= 16'b1111111111011110;
        weights1[44437] <= 16'b1111111111001001;
        weights1[44438] <= 16'b1111111110101101;
        weights1[44439] <= 16'b1111111110000000;
        weights1[44440] <= 16'b1111111101100011;
        weights1[44441] <= 16'b1111111101101010;
        weights1[44442] <= 16'b1111111110000011;
        weights1[44443] <= 16'b1111111110100000;
        weights1[44444] <= 16'b1111111110100010;
        weights1[44445] <= 16'b1111111110111110;
        weights1[44446] <= 16'b1111111111011110;
        weights1[44447] <= 16'b1111111111100111;
        weights1[44448] <= 16'b1111111111101101;
        weights1[44449] <= 16'b1111111111101010;
        weights1[44450] <= 16'b1111111111110001;
        weights1[44451] <= 16'b1111111111110101;
        weights1[44452] <= 16'b1111111111110010;
        weights1[44453] <= 16'b1111111111110000;
        weights1[44454] <= 16'b0000000000000001;
        weights1[44455] <= 16'b1111111111111100;
        weights1[44456] <= 16'b1111111111110100;
        weights1[44457] <= 16'b0000000000000100;
        weights1[44458] <= 16'b1111111111111000;
        weights1[44459] <= 16'b1111111111111011;
        weights1[44460] <= 16'b1111111111110000;
        weights1[44461] <= 16'b0000000000000101;
        weights1[44462] <= 16'b0000000000000001;
        weights1[44463] <= 16'b0000000000000011;
        weights1[44464] <= 16'b1111111111011111;
        weights1[44465] <= 16'b1111111111011010;
        weights1[44466] <= 16'b1111111111010001;
        weights1[44467] <= 16'b1111111110011111;
        weights1[44468] <= 16'b1111111101111101;
        weights1[44469] <= 16'b1111111101000000;
        weights1[44470] <= 16'b1111111100100000;
        weights1[44471] <= 16'b1111111100001100;
        weights1[44472] <= 16'b1111111011101101;
        weights1[44473] <= 16'b1111111011111111;
        weights1[44474] <= 16'b1111111100010000;
        weights1[44475] <= 16'b1111111101101000;
        weights1[44476] <= 16'b1111111110010011;
        weights1[44477] <= 16'b1111111110110110;
        weights1[44478] <= 16'b1111111111010101;
        weights1[44479] <= 16'b1111111111010000;
        weights1[44480] <= 16'b1111111111101111;
        weights1[44481] <= 16'b1111111111111100;
        weights1[44482] <= 16'b1111111111111101;
        weights1[44483] <= 16'b0000000000000011;
        weights1[44484] <= 16'b0000000000000000;
        weights1[44485] <= 16'b0000000000010000;
        weights1[44486] <= 16'b0000000000000110;
        weights1[44487] <= 16'b0000000000000000;
        weights1[44488] <= 16'b1111111111111011;
        weights1[44489] <= 16'b0000000000010010;
        weights1[44490] <= 16'b1111111111110101;
        weights1[44491] <= 16'b1111111111101001;
        weights1[44492] <= 16'b1111111111110000;
        weights1[44493] <= 16'b1111111111110101;
        weights1[44494] <= 16'b1111111111101101;
        weights1[44495] <= 16'b1111111111011101;
        weights1[44496] <= 16'b1111111111000110;
        weights1[44497] <= 16'b1111111110101001;
        weights1[44498] <= 16'b1111111110101100;
        weights1[44499] <= 16'b1111111110000111;
        weights1[44500] <= 16'b1111111101110111;
        weights1[44501] <= 16'b1111111110000010;
        weights1[44502] <= 16'b1111111110011110;
        weights1[44503] <= 16'b1111111110101010;
        weights1[44504] <= 16'b1111111111000000;
        weights1[44505] <= 16'b1111111111011001;
        weights1[44506] <= 16'b1111111111110001;
        weights1[44507] <= 16'b1111111111111001;
        weights1[44508] <= 16'b1111111111110010;
        weights1[44509] <= 16'b1111111111110111;
        weights1[44510] <= 16'b0000000000001111;
        weights1[44511] <= 16'b1111111111111110;
        weights1[44512] <= 16'b0000000000010001;
        weights1[44513] <= 16'b0000000000000010;
        weights1[44514] <= 16'b0000000000001000;
        weights1[44515] <= 16'b0000000000001101;
        weights1[44516] <= 16'b1111111111111111;
        weights1[44517] <= 16'b0000000000000110;
        weights1[44518] <= 16'b1111111111111100;
        weights1[44519] <= 16'b1111111111100111;
        weights1[44520] <= 16'b1111111111101011;
        weights1[44521] <= 16'b1111111111110101;
        weights1[44522] <= 16'b0000000000001100;
        weights1[44523] <= 16'b0000000000010011;
        weights1[44524] <= 16'b0000000000001000;
        weights1[44525] <= 16'b0000000000000000;
        weights1[44526] <= 16'b0000000000001101;
        weights1[44527] <= 16'b0000000000001011;
        weights1[44528] <= 16'b0000000001000000;
        weights1[44529] <= 16'b0000000000100010;
        weights1[44530] <= 16'b0000000000111000;
        weights1[44531] <= 16'b0000000000101101;
        weights1[44532] <= 16'b0000000000011101;
        weights1[44533] <= 16'b0000000000010001;
        weights1[44534] <= 16'b0000000000000110;
        weights1[44535] <= 16'b0000000000000100;
        weights1[44536] <= 16'b0000000000000010;
        weights1[44537] <= 16'b0000000000000000;
        weights1[44538] <= 16'b1111111111101110;
        weights1[44539] <= 16'b1111111111101111;
        weights1[44540] <= 16'b0000000000001111;
        weights1[44541] <= 16'b1111111111111101;
        weights1[44542] <= 16'b0000000000000110;
        weights1[44543] <= 16'b0000000000000101;
        weights1[44544] <= 16'b0000000000000010;
        weights1[44545] <= 16'b0000000000000011;
        weights1[44546] <= 16'b1111111111110011;
        weights1[44547] <= 16'b1111111111101101;
        weights1[44548] <= 16'b1111111111110110;
        weights1[44549] <= 16'b1111111111110110;
        weights1[44550] <= 16'b0000000000001100;
        weights1[44551] <= 16'b0000000000011111;
        weights1[44552] <= 16'b0000000000101000;
        weights1[44553] <= 16'b0000000000110111;
        weights1[44554] <= 16'b0000000001000101;
        weights1[44555] <= 16'b0000000001001100;
        weights1[44556] <= 16'b0000000000111100;
        weights1[44557] <= 16'b0000000001010001;
        weights1[44558] <= 16'b0000000001000010;
        weights1[44559] <= 16'b0000000000101101;
        weights1[44560] <= 16'b0000000000011010;
        weights1[44561] <= 16'b0000000000010110;
        weights1[44562] <= 16'b0000000000000111;
        weights1[44563] <= 16'b0000000000000000;
        weights1[44564] <= 16'b1111111111110001;
        weights1[44565] <= 16'b0000000000000010;
        weights1[44566] <= 16'b1111111111110011;
        weights1[44567] <= 16'b0000000000000001;
        weights1[44568] <= 16'b1111111111111110;
        weights1[44569] <= 16'b1111111111111100;
        weights1[44570] <= 16'b0000000000000010;
        weights1[44571] <= 16'b0000000000000101;
        weights1[44572] <= 16'b1111111111111111;
        weights1[44573] <= 16'b0000000000000011;
        weights1[44574] <= 16'b1111111111111110;
        weights1[44575] <= 16'b1111111111101101;
        weights1[44576] <= 16'b1111111111111111;
        weights1[44577] <= 16'b0000000000000000;
        weights1[44578] <= 16'b1111111111111111;
        weights1[44579] <= 16'b0000000000010101;
        weights1[44580] <= 16'b0000000000100101;
        weights1[44581] <= 16'b0000000000101110;
        weights1[44582] <= 16'b0000000000110111;
        weights1[44583] <= 16'b0000000000101011;
        weights1[44584] <= 16'b0000000000100000;
        weights1[44585] <= 16'b0000000000100001;
        weights1[44586] <= 16'b0000000000011110;
        weights1[44587] <= 16'b0000000000000101;
        weights1[44588] <= 16'b0000000000010101;
        weights1[44589] <= 16'b0000000000000011;
        weights1[44590] <= 16'b0000000000010000;
        weights1[44591] <= 16'b1111111111111001;
        weights1[44592] <= 16'b1111111111111000;
        weights1[44593] <= 16'b0000000000000011;
        weights1[44594] <= 16'b1111111111111001;
        weights1[44595] <= 16'b1111111111101010;
        weights1[44596] <= 16'b1111111111111011;
        weights1[44597] <= 16'b0000000000001010;
        weights1[44598] <= 16'b0000000000001110;
        weights1[44599] <= 16'b0000000000010010;
        weights1[44600] <= 16'b0000000000000000;
        weights1[44601] <= 16'b1111111111100100;
        weights1[44602] <= 16'b1111111111111100;
        weights1[44603] <= 16'b1111111111110010;
        weights1[44604] <= 16'b0000000000000101;
        weights1[44605] <= 16'b0000000000000110;
        weights1[44606] <= 16'b0000000000010011;
        weights1[44607] <= 16'b0000000000100000;
        weights1[44608] <= 16'b0000000000011101;
        weights1[44609] <= 16'b0000000000111111;
        weights1[44610] <= 16'b0000000000011110;
        weights1[44611] <= 16'b0000000000001110;
        weights1[44612] <= 16'b0000000000001110;
        weights1[44613] <= 16'b0000000000011001;
        weights1[44614] <= 16'b0000000000000100;
        weights1[44615] <= 16'b0000000000010010;
        weights1[44616] <= 16'b0000000000000011;
        weights1[44617] <= 16'b1111111111111100;
        weights1[44618] <= 16'b0000000000000100;
        weights1[44619] <= 16'b0000000000000011;
        weights1[44620] <= 16'b0000000000000110;
        weights1[44621] <= 16'b0000000000000011;
        weights1[44622] <= 16'b1111111111111111;
        weights1[44623] <= 16'b1111111111111111;
        weights1[44624] <= 16'b0000000000000000;
        weights1[44625] <= 16'b1111111111110100;
        weights1[44626] <= 16'b1111111111111110;
        weights1[44627] <= 16'b0000000000001111;
        weights1[44628] <= 16'b0000000000001101;
        weights1[44629] <= 16'b0000000000000100;
        weights1[44630] <= 16'b1111111111111000;
        weights1[44631] <= 16'b1111111111111100;
        weights1[44632] <= 16'b0000000000000011;
        weights1[44633] <= 16'b0000000000001001;
        weights1[44634] <= 16'b0000000000001111;
        weights1[44635] <= 16'b0000000000011010;
        weights1[44636] <= 16'b0000000000001000;
        weights1[44637] <= 16'b0000000000011111;
        weights1[44638] <= 16'b0000000000010101;
        weights1[44639] <= 16'b0000000000000101;
        weights1[44640] <= 16'b0000000000011011;
        weights1[44641] <= 16'b0000000000001110;
        weights1[44642] <= 16'b0000000000000111;
        weights1[44643] <= 16'b0000000000000110;
        weights1[44644] <= 16'b0000000000001001;
        weights1[44645] <= 16'b0000000000010000;
        weights1[44646] <= 16'b0000000000000110;
        weights1[44647] <= 16'b1111111111111000;
        weights1[44648] <= 16'b0000000000000000;
        weights1[44649] <= 16'b1111111111101110;
        weights1[44650] <= 16'b0000000000000000;
        weights1[44651] <= 16'b1111111111111010;
        weights1[44652] <= 16'b1111111111111011;
        weights1[44653] <= 16'b0000000000000010;
        weights1[44654] <= 16'b1111111111111000;
        weights1[44655] <= 16'b1111111111110111;
        weights1[44656] <= 16'b1111111111111111;
        weights1[44657] <= 16'b0000000000000011;
        weights1[44658] <= 16'b1111111111111001;
        weights1[44659] <= 16'b0000000000000010;
        weights1[44660] <= 16'b0000000000001010;
        weights1[44661] <= 16'b0000000000010100;
        weights1[44662] <= 16'b0000000000010100;
        weights1[44663] <= 16'b0000000000001001;
        weights1[44664] <= 16'b0000000000011010;
        weights1[44665] <= 16'b0000000000011011;
        weights1[44666] <= 16'b0000000000010000;
        weights1[44667] <= 16'b0000000000000011;
        weights1[44668] <= 16'b0000000000001100;
        weights1[44669] <= 16'b0000000000000101;
        weights1[44670] <= 16'b0000000000000011;
        weights1[44671] <= 16'b0000000000000000;
        weights1[44672] <= 16'b1111111111111010;
        weights1[44673] <= 16'b1111111111110011;
        weights1[44674] <= 16'b1111111111110111;
        weights1[44675] <= 16'b1111111111110100;
        weights1[44676] <= 16'b0000000000000100;
        weights1[44677] <= 16'b1111111111111110;
        weights1[44678] <= 16'b1111111111111001;
        weights1[44679] <= 16'b1111111111110011;
        weights1[44680] <= 16'b1111111111110111;
        weights1[44681] <= 16'b1111111111110110;
        weights1[44682] <= 16'b0000000000000001;
        weights1[44683] <= 16'b1111111111111011;
        weights1[44684] <= 16'b1111111111110110;
        weights1[44685] <= 16'b0000000000000001;
        weights1[44686] <= 16'b1111111111111011;
        weights1[44687] <= 16'b0000000000000000;
        weights1[44688] <= 16'b1111111111111111;
        weights1[44689] <= 16'b0000000000000000;
        weights1[44690] <= 16'b0000000000000000;
        weights1[44691] <= 16'b0000000000000001;
        weights1[44692] <= 16'b0000000000000011;
        weights1[44693] <= 16'b0000000000001111;
        weights1[44694] <= 16'b0000000000011111;
        weights1[44695] <= 16'b0000000000101000;
        weights1[44696] <= 16'b0000000000100010;
        weights1[44697] <= 16'b0000000000011110;
        weights1[44698] <= 16'b0000000000001000;
        weights1[44699] <= 16'b1111111111001110;
        weights1[44700] <= 16'b1111111110100111;
        weights1[44701] <= 16'b1111111110011001;
        weights1[44702] <= 16'b1111111110011111;
        weights1[44703] <= 16'b1111111110111111;
        weights1[44704] <= 16'b1111111111010011;
        weights1[44705] <= 16'b1111111111110110;
        weights1[44706] <= 16'b0000000000000011;
        weights1[44707] <= 16'b0000000000001101;
        weights1[44708] <= 16'b0000000000001110;
        weights1[44709] <= 16'b0000000000010010;
        weights1[44710] <= 16'b0000000000000001;
        weights1[44711] <= 16'b1111111111111010;
        weights1[44712] <= 16'b1111111111110100;
        weights1[44713] <= 16'b1111111111111000;
        weights1[44714] <= 16'b1111111111111001;
        weights1[44715] <= 16'b0000000000000001;
        weights1[44716] <= 16'b1111111111111111;
        weights1[44717] <= 16'b0000000000000011;
        weights1[44718] <= 16'b0000000000000111;
        weights1[44719] <= 16'b0000000000000100;
        weights1[44720] <= 16'b0000000000001011;
        weights1[44721] <= 16'b0000000000001110;
        weights1[44722] <= 16'b0000000000100100;
        weights1[44723] <= 16'b0000000000101111;
        weights1[44724] <= 16'b0000000000011011;
        weights1[44725] <= 16'b0000000000010100;
        weights1[44726] <= 16'b1111111111110101;
        weights1[44727] <= 16'b1111111111001010;
        weights1[44728] <= 16'b1111111110001000;
        weights1[44729] <= 16'b1111111110000001;
        weights1[44730] <= 16'b1111111110101011;
        weights1[44731] <= 16'b1111111111100100;
        weights1[44732] <= 16'b1111111111101011;
        weights1[44733] <= 16'b1111111111111101;
        weights1[44734] <= 16'b0000000000001111;
        weights1[44735] <= 16'b0000000000010101;
        weights1[44736] <= 16'b0000000000010110;
        weights1[44737] <= 16'b0000000000010001;
        weights1[44738] <= 16'b0000000000000111;
        weights1[44739] <= 16'b1111111111111011;
        weights1[44740] <= 16'b1111111111101111;
        weights1[44741] <= 16'b1111111111100101;
        weights1[44742] <= 16'b1111111111110011;
        weights1[44743] <= 16'b1111111111111010;
        weights1[44744] <= 16'b1111111111111111;
        weights1[44745] <= 16'b0000000000000011;
        weights1[44746] <= 16'b0000000000000000;
        weights1[44747] <= 16'b1111111111111111;
        weights1[44748] <= 16'b0000000000000001;
        weights1[44749] <= 16'b0000000000010100;
        weights1[44750] <= 16'b0000000000100010;
        weights1[44751] <= 16'b0000000000110110;
        weights1[44752] <= 16'b0000000000011011;
        weights1[44753] <= 16'b0000000000001110;
        weights1[44754] <= 16'b1111111111100010;
        weights1[44755] <= 16'b1111111110011011;
        weights1[44756] <= 16'b1111111101101101;
        weights1[44757] <= 16'b1111111110001100;
        weights1[44758] <= 16'b1111111110111100;
        weights1[44759] <= 16'b1111111111110010;
        weights1[44760] <= 16'b0000000000011011;
        weights1[44761] <= 16'b0000000000001111;
        weights1[44762] <= 16'b0000000000011111;
        weights1[44763] <= 16'b0000000000010101;
        weights1[44764] <= 16'b0000000000010001;
        weights1[44765] <= 16'b1111111111111110;
        weights1[44766] <= 16'b1111111111111000;
        weights1[44767] <= 16'b1111111111011101;
        weights1[44768] <= 16'b1111111111010011;
        weights1[44769] <= 16'b1111111111100010;
        weights1[44770] <= 16'b1111111111100110;
        weights1[44771] <= 16'b1111111111101111;
        weights1[44772] <= 16'b0000000000000011;
        weights1[44773] <= 16'b0000000000000011;
        weights1[44774] <= 16'b1111111111111001;
        weights1[44775] <= 16'b0000000000000001;
        weights1[44776] <= 16'b0000000000000110;
        weights1[44777] <= 16'b0000000000011110;
        weights1[44778] <= 16'b0000000000011101;
        weights1[44779] <= 16'b0000000000101010;
        weights1[44780] <= 16'b0000000000010101;
        weights1[44781] <= 16'b0000000000010101;
        weights1[44782] <= 16'b1111111111110000;
        weights1[44783] <= 16'b1111111110000011;
        weights1[44784] <= 16'b1111111101010011;
        weights1[44785] <= 16'b1111111101100110;
        weights1[44786] <= 16'b1111111110110001;
        weights1[44787] <= 16'b1111111111110111;
        weights1[44788] <= 16'b1111111111101011;
        weights1[44789] <= 16'b0000000000000011;
        weights1[44790] <= 16'b0000000000110100;
        weights1[44791] <= 16'b0000000000101010;
        weights1[44792] <= 16'b0000000000011001;
        weights1[44793] <= 16'b0000000000001101;
        weights1[44794] <= 16'b1111111111101111;
        weights1[44795] <= 16'b1111111111000111;
        weights1[44796] <= 16'b1111111111000011;
        weights1[44797] <= 16'b1111111111011000;
        weights1[44798] <= 16'b1111111111100101;
        weights1[44799] <= 16'b1111111111110110;
        weights1[44800] <= 16'b0000000000000001;
        weights1[44801] <= 16'b1111111111111100;
        weights1[44802] <= 16'b1111111111111110;
        weights1[44803] <= 16'b0000000000000110;
        weights1[44804] <= 16'b0000000000001110;
        weights1[44805] <= 16'b0000000000101010;
        weights1[44806] <= 16'b0000000000010010;
        weights1[44807] <= 16'b0000000000100001;
        weights1[44808] <= 16'b0000000000100000;
        weights1[44809] <= 16'b0000000000100000;
        weights1[44810] <= 16'b1111111111100011;
        weights1[44811] <= 16'b1111111101100101;
        weights1[44812] <= 16'b1111111100111110;
        weights1[44813] <= 16'b1111111101001101;
        weights1[44814] <= 16'b1111111111001111;
        weights1[44815] <= 16'b0000000000001111;
        weights1[44816] <= 16'b0000000000001011;
        weights1[44817] <= 16'b0000000000011111;
        weights1[44818] <= 16'b0000000000010010;
        weights1[44819] <= 16'b0000000000001100;
        weights1[44820] <= 16'b0000000000001111;
        weights1[44821] <= 16'b1111111111011110;
        weights1[44822] <= 16'b1111111111001110;
        weights1[44823] <= 16'b1111111110111001;
        weights1[44824] <= 16'b1111111110111000;
        weights1[44825] <= 16'b1111111111011001;
        weights1[44826] <= 16'b1111111111101101;
        weights1[44827] <= 16'b1111111111111100;
        weights1[44828] <= 16'b1111111111111100;
        weights1[44829] <= 16'b1111111111111001;
        weights1[44830] <= 16'b1111111111110111;
        weights1[44831] <= 16'b1111111111110101;
        weights1[44832] <= 16'b0000000000000011;
        weights1[44833] <= 16'b0000000000011110;
        weights1[44834] <= 16'b0000000000100011;
        weights1[44835] <= 16'b0000000000111000;
        weights1[44836] <= 16'b0000000000100100;
        weights1[44837] <= 16'b0000000000011111;
        weights1[44838] <= 16'b1111111111010011;
        weights1[44839] <= 16'b1111111101001000;
        weights1[44840] <= 16'b1111111100101000;
        weights1[44841] <= 16'b1111111101110101;
        weights1[44842] <= 16'b0000000000111111;
        weights1[44843] <= 16'b0000000000111100;
        weights1[44844] <= 16'b0000000000011001;
        weights1[44845] <= 16'b0000000000110101;
        weights1[44846] <= 16'b0000000000101101;
        weights1[44847] <= 16'b0000000000011000;
        weights1[44848] <= 16'b1111111111110010;
        weights1[44849] <= 16'b1111111111001000;
        weights1[44850] <= 16'b1111111110110010;
        weights1[44851] <= 16'b1111111110101111;
        weights1[44852] <= 16'b1111111111000110;
        weights1[44853] <= 16'b1111111111011101;
        weights1[44854] <= 16'b1111111111101011;
        weights1[44855] <= 16'b1111111111110011;
        weights1[44856] <= 16'b1111111111110100;
        weights1[44857] <= 16'b1111111111110010;
        weights1[44858] <= 16'b1111111111101000;
        weights1[44859] <= 16'b1111111111110111;
        weights1[44860] <= 16'b1111111111111011;
        weights1[44861] <= 16'b0000000000000010;
        weights1[44862] <= 16'b0000000000011101;
        weights1[44863] <= 16'b0000000000100011;
        weights1[44864] <= 16'b0000000000101100;
        weights1[44865] <= 16'b0000000000111011;
        weights1[44866] <= 16'b1111111110110001;
        weights1[44867] <= 16'b1111111101001111;
        weights1[44868] <= 16'b1111111100111001;
        weights1[44869] <= 16'b1111111111000000;
        weights1[44870] <= 16'b0000000000100000;
        weights1[44871] <= 16'b0000000000111010;
        weights1[44872] <= 16'b0000000000011111;
        weights1[44873] <= 16'b0000000000010111;
        weights1[44874] <= 16'b0000000000001101;
        weights1[44875] <= 16'b0000000000010011;
        weights1[44876] <= 16'b1111111111001110;
        weights1[44877] <= 16'b1111111110101100;
        weights1[44878] <= 16'b1111111110010001;
        weights1[44879] <= 16'b1111111110010110;
        weights1[44880] <= 16'b1111111111001011;
        weights1[44881] <= 16'b1111111111100001;
        weights1[44882] <= 16'b1111111111111010;
        weights1[44883] <= 16'b0000000000000100;
        weights1[44884] <= 16'b1111111111110010;
        weights1[44885] <= 16'b1111111111011111;
        weights1[44886] <= 16'b1111111111011101;
        weights1[44887] <= 16'b1111111111110111;
        weights1[44888] <= 16'b1111111111100101;
        weights1[44889] <= 16'b1111111111111111;
        weights1[44890] <= 16'b0000000000010101;
        weights1[44891] <= 16'b0000000000011001;
        weights1[44892] <= 16'b0000000000101101;
        weights1[44893] <= 16'b0000000000111110;
        weights1[44894] <= 16'b1111111111000100;
        weights1[44895] <= 16'b1111111100100101;
        weights1[44896] <= 16'b1111111101100110;
        weights1[44897] <= 16'b1111111111110101;
        weights1[44898] <= 16'b0000000000100101;
        weights1[44899] <= 16'b0000000000101101;
        weights1[44900] <= 16'b0000000000011111;
        weights1[44901] <= 16'b0000000000101011;
        weights1[44902] <= 16'b0000000000001001;
        weights1[44903] <= 16'b1111111111111101;
        weights1[44904] <= 16'b1111111111011001;
        weights1[44905] <= 16'b1111111110010111;
        weights1[44906] <= 16'b1111111110011010;
        weights1[44907] <= 16'b1111111111000101;
        weights1[44908] <= 16'b1111111111111100;
        weights1[44909] <= 16'b1111111111111101;
        weights1[44910] <= 16'b0000000000010000;
        weights1[44911] <= 16'b0000000000001111;
        weights1[44912] <= 16'b1111111111110110;
        weights1[44913] <= 16'b1111111111101011;
        weights1[44914] <= 16'b1111111111101011;
        weights1[44915] <= 16'b1111111111111000;
        weights1[44916] <= 16'b0000000000001100;
        weights1[44917] <= 16'b0000000000001000;
        weights1[44918] <= 16'b0000000000010000;
        weights1[44919] <= 16'b0000000000011110;
        weights1[44920] <= 16'b0000000000111000;
        weights1[44921] <= 16'b0000000000101100;
        weights1[44922] <= 16'b1111111111000110;
        weights1[44923] <= 16'b1111111101001000;
        weights1[44924] <= 16'b1111111110111100;
        weights1[44925] <= 16'b1111111111110000;
        weights1[44926] <= 16'b0000000000001101;
        weights1[44927] <= 16'b0000000000111010;
        weights1[44928] <= 16'b0000000000011101;
        weights1[44929] <= 16'b0000000000010010;
        weights1[44930] <= 16'b0000000000000010;
        weights1[44931] <= 16'b1111111111011110;
        weights1[44932] <= 16'b1111111110111001;
        weights1[44933] <= 16'b1111111110010011;
        weights1[44934] <= 16'b1111111111001110;
        weights1[44935] <= 16'b0000000000001101;
        weights1[44936] <= 16'b0000000000010100;
        weights1[44937] <= 16'b0000000000010001;
        weights1[44938] <= 16'b0000000000100010;
        weights1[44939] <= 16'b0000000000011111;
        weights1[44940] <= 16'b1111111111110111;
        weights1[44941] <= 16'b1111111111101100;
        weights1[44942] <= 16'b1111111111110100;
        weights1[44943] <= 16'b1111111111101001;
        weights1[44944] <= 16'b0000000000000010;
        weights1[44945] <= 16'b0000000000000001;
        weights1[44946] <= 16'b0000000000000100;
        weights1[44947] <= 16'b0000000000010101;
        weights1[44948] <= 16'b0000000000001110;
        weights1[44949] <= 16'b0000000000110110;
        weights1[44950] <= 16'b1111111111001001;
        weights1[44951] <= 16'b1111111110100100;
        weights1[44952] <= 16'b1111111111000100;
        weights1[44953] <= 16'b1111111111111100;
        weights1[44954] <= 16'b0000000000011011;
        weights1[44955] <= 16'b0000000000011011;
        weights1[44956] <= 16'b0000000000010011;
        weights1[44957] <= 16'b0000000000011111;
        weights1[44958] <= 16'b1111111111101011;
        weights1[44959] <= 16'b1111111111011110;
        weights1[44960] <= 16'b1111111110101110;
        weights1[44961] <= 16'b1111111110110001;
        weights1[44962] <= 16'b0000000000001001;
        weights1[44963] <= 16'b0000000000100100;
        weights1[44964] <= 16'b0000000000011110;
        weights1[44965] <= 16'b0000000000010000;
        weights1[44966] <= 16'b0000000000011110;
        weights1[44967] <= 16'b0000000000001110;
        weights1[44968] <= 16'b1111111111110111;
        weights1[44969] <= 16'b1111111111110010;
        weights1[44970] <= 16'b1111111111111011;
        weights1[44971] <= 16'b0000000000001001;
        weights1[44972] <= 16'b0000000000001100;
        weights1[44973] <= 16'b1111111111111100;
        weights1[44974] <= 16'b1111111111111100;
        weights1[44975] <= 16'b0000000000010010;
        weights1[44976] <= 16'b0000000000010011;
        weights1[44977] <= 16'b0000000000100000;
        weights1[44978] <= 16'b1111111111011011;
        weights1[44979] <= 16'b1111111111000100;
        weights1[44980] <= 16'b1111111111100101;
        weights1[44981] <= 16'b0000000000000001;
        weights1[44982] <= 16'b0000000000000100;
        weights1[44983] <= 16'b0000000000100001;
        weights1[44984] <= 16'b0000000000001111;
        weights1[44985] <= 16'b0000000000000010;
        weights1[44986] <= 16'b1111111111101101;
        weights1[44987] <= 16'b1111111111010100;
        weights1[44988] <= 16'b1111111111001011;
        weights1[44989] <= 16'b1111111111101000;
        weights1[44990] <= 16'b0000000000100101;
        weights1[44991] <= 16'b0000000000010111;
        weights1[44992] <= 16'b0000000000011111;
        weights1[44993] <= 16'b0000000000101000;
        weights1[44994] <= 16'b0000000000001111;
        weights1[44995] <= 16'b0000000000001001;
        weights1[44996] <= 16'b1111111111110111;
        weights1[44997] <= 16'b1111111111110110;
        weights1[44998] <= 16'b1111111111101001;
        weights1[44999] <= 16'b1111111111111001;
        weights1[45000] <= 16'b1111111111110100;
        weights1[45001] <= 16'b1111111111110100;
        weights1[45002] <= 16'b0000000000010001;
        weights1[45003] <= 16'b1111111111110001;
        weights1[45004] <= 16'b0000000000001101;
        weights1[45005] <= 16'b0000000000010110;
        weights1[45006] <= 16'b1111111111101111;
        weights1[45007] <= 16'b1111111111100001;
        weights1[45008] <= 16'b1111111111100010;
        weights1[45009] <= 16'b0000000000001000;
        weights1[45010] <= 16'b0000000000001000;
        weights1[45011] <= 16'b1111111111111011;
        weights1[45012] <= 16'b1111111111111011;
        weights1[45013] <= 16'b1111111111111010;
        weights1[45014] <= 16'b1111111111111110;
        weights1[45015] <= 16'b1111111111000010;
        weights1[45016] <= 16'b1111111111101100;
        weights1[45017] <= 16'b1111111111111101;
        weights1[45018] <= 16'b0000000000010010;
        weights1[45019] <= 16'b0000000000010010;
        weights1[45020] <= 16'b0000000000000111;
        weights1[45021] <= 16'b0000000000001100;
        weights1[45022] <= 16'b1111111111111111;
        weights1[45023] <= 16'b0000000000001001;
        weights1[45024] <= 16'b1111111111110100;
        weights1[45025] <= 16'b1111111111110010;
        weights1[45026] <= 16'b0000000000000111;
        weights1[45027] <= 16'b0000000000000000;
        weights1[45028] <= 16'b1111111111111100;
        weights1[45029] <= 16'b0000000000000100;
        weights1[45030] <= 16'b0000000000001010;
        weights1[45031] <= 16'b0000000000000101;
        weights1[45032] <= 16'b0000000000010101;
        weights1[45033] <= 16'b0000000000001010;
        weights1[45034] <= 16'b1111111111111100;
        weights1[45035] <= 16'b1111111111100100;
        weights1[45036] <= 16'b1111111111110001;
        weights1[45037] <= 16'b0000000000001111;
        weights1[45038] <= 16'b0000000000000000;
        weights1[45039] <= 16'b0000000000000011;
        weights1[45040] <= 16'b0000000000010010;
        weights1[45041] <= 16'b1111111111110001;
        weights1[45042] <= 16'b1111111111101111;
        weights1[45043] <= 16'b1111111111010001;
        weights1[45044] <= 16'b1111111111110100;
        weights1[45045] <= 16'b0000000000010101;
        weights1[45046] <= 16'b0000000000010111;
        weights1[45047] <= 16'b0000000000000011;
        weights1[45048] <= 16'b0000000000001010;
        weights1[45049] <= 16'b0000000000001000;
        weights1[45050] <= 16'b0000000000000110;
        weights1[45051] <= 16'b0000000000001111;
        weights1[45052] <= 16'b1111111111110011;
        weights1[45053] <= 16'b1111111111111100;
        weights1[45054] <= 16'b1111111111111010;
        weights1[45055] <= 16'b1111111111110010;
        weights1[45056] <= 16'b0000000000000001;
        weights1[45057] <= 16'b0000000000001000;
        weights1[45058] <= 16'b0000000000000000;
        weights1[45059] <= 16'b0000000000000100;
        weights1[45060] <= 16'b0000000000000010;
        weights1[45061] <= 16'b0000000000010000;
        weights1[45062] <= 16'b0000000000001001;
        weights1[45063] <= 16'b0000000000000001;
        weights1[45064] <= 16'b0000000000000011;
        weights1[45065] <= 16'b1111111111111100;
        weights1[45066] <= 16'b1111111111110010;
        weights1[45067] <= 16'b0000000000000000;
        weights1[45068] <= 16'b1111111111110011;
        weights1[45069] <= 16'b1111111111100010;
        weights1[45070] <= 16'b0000000000000000;
        weights1[45071] <= 16'b1111111111101110;
        weights1[45072] <= 16'b0000000000000111;
        weights1[45073] <= 16'b0000000000001001;
        weights1[45074] <= 16'b0000000000010111;
        weights1[45075] <= 16'b0000000000001100;
        weights1[45076] <= 16'b1111111111110010;
        weights1[45077] <= 16'b0000000000000000;
        weights1[45078] <= 16'b0000000000001000;
        weights1[45079] <= 16'b0000000000010001;
        weights1[45080] <= 16'b1111111111111011;
        weights1[45081] <= 16'b1111111111110011;
        weights1[45082] <= 16'b1111111111101010;
        weights1[45083] <= 16'b1111111111111100;
        weights1[45084] <= 16'b1111111111101101;
        weights1[45085] <= 16'b0000000000001111;
        weights1[45086] <= 16'b1111111111111011;
        weights1[45087] <= 16'b0000000000001010;
        weights1[45088] <= 16'b0000000000001110;
        weights1[45089] <= 16'b0000000000000111;
        weights1[45090] <= 16'b0000000000000011;
        weights1[45091] <= 16'b0000000000001111;
        weights1[45092] <= 16'b1111111111111101;
        weights1[45093] <= 16'b0000000000000100;
        weights1[45094] <= 16'b0000000000000101;
        weights1[45095] <= 16'b1111111111110110;
        weights1[45096] <= 16'b1111111111111010;
        weights1[45097] <= 16'b0000000000010000;
        weights1[45098] <= 16'b0000000000000001;
        weights1[45099] <= 16'b0000000000001101;
        weights1[45100] <= 16'b0000000000001010;
        weights1[45101] <= 16'b0000000000000110;
        weights1[45102] <= 16'b0000000000000101;
        weights1[45103] <= 16'b1111111111111000;
        weights1[45104] <= 16'b0000000000001110;
        weights1[45105] <= 16'b0000000000000101;
        weights1[45106] <= 16'b0000000000000101;
        weights1[45107] <= 16'b1111111111111110;
        weights1[45108] <= 16'b1111111111110100;
        weights1[45109] <= 16'b1111111111110011;
        weights1[45110] <= 16'b1111111111111101;
        weights1[45111] <= 16'b1111111111110010;
        weights1[45112] <= 16'b1111111111111011;
        weights1[45113] <= 16'b0000000000001010;
        weights1[45114] <= 16'b0000000000000000;
        weights1[45115] <= 16'b0000000000010110;
        weights1[45116] <= 16'b0000000000010010;
        weights1[45117] <= 16'b0000000000010100;
        weights1[45118] <= 16'b1111111111111101;
        weights1[45119] <= 16'b0000000000010101;
        weights1[45120] <= 16'b1111111111110110;
        weights1[45121] <= 16'b1111111111110000;
        weights1[45122] <= 16'b0000000000000001;
        weights1[45123] <= 16'b1111111111111010;
        weights1[45124] <= 16'b1111111111100010;
        weights1[45125] <= 16'b0000000000001011;
        weights1[45126] <= 16'b1111111111111101;
        weights1[45127] <= 16'b0000000000001000;
        weights1[45128] <= 16'b0000000000010011;
        weights1[45129] <= 16'b0000000000010001;
        weights1[45130] <= 16'b0000000000000110;
        weights1[45131] <= 16'b0000000000001010;
        weights1[45132] <= 16'b0000000000000111;
        weights1[45133] <= 16'b1111111111111011;
        weights1[45134] <= 16'b0000000000000100;
        weights1[45135] <= 16'b1111111111111110;
        weights1[45136] <= 16'b1111111111111000;
        weights1[45137] <= 16'b1111111111111011;
        weights1[45138] <= 16'b0000000000000101;
        weights1[45139] <= 16'b1111111111111111;
        weights1[45140] <= 16'b0000000000000111;
        weights1[45141] <= 16'b0000000000001101;
        weights1[45142] <= 16'b0000000000001110;
        weights1[45143] <= 16'b0000000000000010;
        weights1[45144] <= 16'b1111111111111010;
        weights1[45145] <= 16'b0000000000001001;
        weights1[45146] <= 16'b0000000000001000;
        weights1[45147] <= 16'b1111111111110101;
        weights1[45148] <= 16'b0000000000010110;
        weights1[45149] <= 16'b0000000000001001;
        weights1[45150] <= 16'b0000000000000000;
        weights1[45151] <= 16'b1111111111110011;
        weights1[45152] <= 16'b0000000000000001;
        weights1[45153] <= 16'b0000000000000110;
        weights1[45154] <= 16'b1111111111111001;
        weights1[45155] <= 16'b0000000000001000;
        weights1[45156] <= 16'b0000000000001000;
        weights1[45157] <= 16'b0000000000001100;
        weights1[45158] <= 16'b0000000000000000;
        weights1[45159] <= 16'b0000000000000101;
        weights1[45160] <= 16'b1111111111111111;
        weights1[45161] <= 16'b0000000000001001;
        weights1[45162] <= 16'b0000000000010100;
        weights1[45163] <= 16'b1111111111111011;
        weights1[45164] <= 16'b1111111111111101;
        weights1[45165] <= 16'b0000000000001111;
        weights1[45166] <= 16'b0000000000011010;
        weights1[45167] <= 16'b0000000000010011;
        weights1[45168] <= 16'b0000000000011011;
        weights1[45169] <= 16'b0000000000001000;
        weights1[45170] <= 16'b0000000000000101;
        weights1[45171] <= 16'b0000000000000100;
        weights1[45172] <= 16'b0000000000001011;
        weights1[45173] <= 16'b1111111111111110;
        weights1[45174] <= 16'b1111111111111001;
        weights1[45175] <= 16'b0000000000001000;
        weights1[45176] <= 16'b1111111111101101;
        weights1[45177] <= 16'b0000000000000000;
        weights1[45178] <= 16'b0000000000000000;
        weights1[45179] <= 16'b1111111111110000;
        weights1[45180] <= 16'b0000000000000000;
        weights1[45181] <= 16'b1111111111110010;
        weights1[45182] <= 16'b0000000000000011;
        weights1[45183] <= 16'b0000000000001000;
        weights1[45184] <= 16'b0000000000000111;
        weights1[45185] <= 16'b1111111111110101;
        weights1[45186] <= 16'b0000000000000011;
        weights1[45187] <= 16'b0000000000001000;
        weights1[45188] <= 16'b1111111111110101;
        weights1[45189] <= 16'b0000000000001000;
        weights1[45190] <= 16'b0000000000010011;
        weights1[45191] <= 16'b0000000000010110;
        weights1[45192] <= 16'b0000000000000110;
        weights1[45193] <= 16'b0000000000001110;
        weights1[45194] <= 16'b0000000000000101;
        weights1[45195] <= 16'b0000000000010100;
        weights1[45196] <= 16'b1111111111111111;
        weights1[45197] <= 16'b1111111111101100;
        weights1[45198] <= 16'b0000000000000101;
        weights1[45199] <= 16'b1111111111111101;
        weights1[45200] <= 16'b1111111111111000;
        weights1[45201] <= 16'b0000000000011000;
        weights1[45202] <= 16'b1111111111111111;
        weights1[45203] <= 16'b0000000000000001;
        weights1[45204] <= 16'b0000000000000011;
        weights1[45205] <= 16'b1111111111111101;
        weights1[45206] <= 16'b1111111111110110;
        weights1[45207] <= 16'b0000000000000100;
        weights1[45208] <= 16'b1111111111111111;
        weights1[45209] <= 16'b0000000000000000;
        weights1[45210] <= 16'b0000000000001001;
        weights1[45211] <= 16'b0000000000000000;
        weights1[45212] <= 16'b0000000000000011;
        weights1[45213] <= 16'b0000000000011000;
        weights1[45214] <= 16'b1111111111110101;
        weights1[45215] <= 16'b0000000000010010;
        weights1[45216] <= 16'b1111111111110010;
        weights1[45217] <= 16'b0000000000001001;
        weights1[45218] <= 16'b0000000000001110;
        weights1[45219] <= 16'b0000000000010100;
        weights1[45220] <= 16'b0000000000000100;
        weights1[45221] <= 16'b0000000000001011;
        weights1[45222] <= 16'b0000000000001001;
        weights1[45223] <= 16'b1111111111110001;
        weights1[45224] <= 16'b0000000000010000;
        weights1[45225] <= 16'b0000000000010101;
        weights1[45226] <= 16'b0000000000000100;
        weights1[45227] <= 16'b1111111111110100;
        weights1[45228] <= 16'b1111111111110000;
        weights1[45229] <= 16'b0000000000000110;
        weights1[45230] <= 16'b1111111111101011;
        weights1[45231] <= 16'b0000000000000010;
        weights1[45232] <= 16'b0000000000001001;
        weights1[45233] <= 16'b0000000000000010;
        weights1[45234] <= 16'b1111111111110010;
        weights1[45235] <= 16'b0000000000010111;
        weights1[45236] <= 16'b1111111111111101;
        weights1[45237] <= 16'b1111111111110100;
        weights1[45238] <= 16'b0000000000001110;
        weights1[45239] <= 16'b1111111111110110;
        weights1[45240] <= 16'b0000000000000111;
        weights1[45241] <= 16'b1111111111111001;
        weights1[45242] <= 16'b1111111111110001;
        weights1[45243] <= 16'b0000000000010110;
        weights1[45244] <= 16'b0000000000000000;
        weights1[45245] <= 16'b0000000000001011;
        weights1[45246] <= 16'b0000000000001010;
        weights1[45247] <= 16'b0000000000001101;
        weights1[45248] <= 16'b0000000000001010;
        weights1[45249] <= 16'b1111111111110001;
        weights1[45250] <= 16'b0000000000000111;
        weights1[45251] <= 16'b1111111111111100;
        weights1[45252] <= 16'b1111111111111111;
        weights1[45253] <= 16'b1111111111111010;
        weights1[45254] <= 16'b1111111111111100;
        weights1[45255] <= 16'b1111111111100111;
        weights1[45256] <= 16'b0000000000001110;
        weights1[45257] <= 16'b1111111111111000;
        weights1[45258] <= 16'b1111111111110001;
        weights1[45259] <= 16'b0000000000001110;
        weights1[45260] <= 16'b1111111111111010;
        weights1[45261] <= 16'b1111111111101001;
        weights1[45262] <= 16'b1111111111111111;
        weights1[45263] <= 16'b1111111111111110;
        weights1[45264] <= 16'b1111111111111111;
        weights1[45265] <= 16'b0000000000001101;
        weights1[45266] <= 16'b0000000000001101;
        weights1[45267] <= 16'b1111111111111010;
        weights1[45268] <= 16'b0000000000010100;
        weights1[45269] <= 16'b0000000000001111;
        weights1[45270] <= 16'b1111111111110100;
        weights1[45271] <= 16'b1111111111111111;
        weights1[45272] <= 16'b1111111111111111;
        weights1[45273] <= 16'b0000000000010100;
        weights1[45274] <= 16'b0000000000001001;
        weights1[45275] <= 16'b0000000000000101;
        weights1[45276] <= 16'b0000000000010011;
        weights1[45277] <= 16'b0000000000000100;
        weights1[45278] <= 16'b0000000000000101;
        weights1[45279] <= 16'b0000000000000000;
        weights1[45280] <= 16'b0000000000001110;
        weights1[45281] <= 16'b0000000000000010;
        weights1[45282] <= 16'b1111111111101100;
        weights1[45283] <= 16'b0000000000001001;
        weights1[45284] <= 16'b1111111111111000;
        weights1[45285] <= 16'b1111111111110111;
        weights1[45286] <= 16'b1111111111110011;
        weights1[45287] <= 16'b0000000000001110;
        weights1[45288] <= 16'b0000000000001010;
        weights1[45289] <= 16'b0000000000000100;
        weights1[45290] <= 16'b1111111111111110;
        weights1[45291] <= 16'b0000000000000101;
        weights1[45292] <= 16'b1111111111111111;
        weights1[45293] <= 16'b1111111111110111;
        weights1[45294] <= 16'b1111111111111110;
        weights1[45295] <= 16'b1111111111111101;
        weights1[45296] <= 16'b1111111111110110;
        weights1[45297] <= 16'b0000000000000010;
        weights1[45298] <= 16'b0000000000001101;
        weights1[45299] <= 16'b0000000000000100;
        weights1[45300] <= 16'b0000000000001111;
        weights1[45301] <= 16'b0000000000000100;
        weights1[45302] <= 16'b0000000000000000;
        weights1[45303] <= 16'b1111111111111011;
        weights1[45304] <= 16'b0000000000000111;
        weights1[45305] <= 16'b0000000000000100;
        weights1[45306] <= 16'b0000000000000101;
        weights1[45307] <= 16'b1111111111110011;
        weights1[45308] <= 16'b1111111111111110;
        weights1[45309] <= 16'b1111111111110110;
        weights1[45310] <= 16'b1111111111111010;
        weights1[45311] <= 16'b0000000000000111;
        weights1[45312] <= 16'b1111111111101010;
        weights1[45313] <= 16'b1111111111110010;
        weights1[45314] <= 16'b0000000000000100;
        weights1[45315] <= 16'b1111111111100101;
        weights1[45316] <= 16'b1111111111111010;
        weights1[45317] <= 16'b0000000000001100;
        weights1[45318] <= 16'b0000000000001001;
        weights1[45319] <= 16'b0000000000000101;
        weights1[45320] <= 16'b0000000000000000;
        weights1[45321] <= 16'b1111111111111110;
        weights1[45322] <= 16'b1111111111111011;
        weights1[45323] <= 16'b0000000000000011;
        weights1[45324] <= 16'b1111111111111100;
        weights1[45325] <= 16'b0000000000001110;
        weights1[45326] <= 16'b0000000000000000;
        weights1[45327] <= 16'b0000000000000011;
        weights1[45328] <= 16'b0000000000000111;
        weights1[45329] <= 16'b1111111111111011;
        weights1[45330] <= 16'b1111111111110101;
        weights1[45331] <= 16'b1111111111110110;
        weights1[45332] <= 16'b1111111111111010;
        weights1[45333] <= 16'b1111111111111011;
        weights1[45334] <= 16'b1111111111110011;
        weights1[45335] <= 16'b0000000000000010;
        weights1[45336] <= 16'b1111111111111010;
        weights1[45337] <= 16'b0000000000010001;
        weights1[45338] <= 16'b1111111111110101;
        weights1[45339] <= 16'b1111111111111101;
        weights1[45340] <= 16'b1111111111101100;
        weights1[45341] <= 16'b0000000000000001;
        weights1[45342] <= 16'b1111111111111001;
        weights1[45343] <= 16'b0000000000000010;
        weights1[45344] <= 16'b1111111111110011;
        weights1[45345] <= 16'b1111111111111001;
        weights1[45346] <= 16'b0000000000001111;
        weights1[45347] <= 16'b1111111111111100;
        weights1[45348] <= 16'b0000000000001001;
        weights1[45349] <= 16'b0000000000001001;
        weights1[45350] <= 16'b0000000000001101;
        weights1[45351] <= 16'b0000000000001100;
        weights1[45352] <= 16'b0000000000000011;
        weights1[45353] <= 16'b1111111111111001;
        weights1[45354] <= 16'b1111111111111110;
        weights1[45355] <= 16'b1111111111110110;
        weights1[45356] <= 16'b1111111111111011;
        weights1[45357] <= 16'b1111111111110101;
        weights1[45358] <= 16'b1111111111111010;
        weights1[45359] <= 16'b1111111111110000;
        weights1[45360] <= 16'b0000000000000000;
        weights1[45361] <= 16'b0000000000000011;
        weights1[45362] <= 16'b0000000000000101;
        weights1[45363] <= 16'b1111111111110101;
        weights1[45364] <= 16'b0000000000000100;
        weights1[45365] <= 16'b1111111111111011;
        weights1[45366] <= 16'b0000000000000001;
        weights1[45367] <= 16'b0000000000000100;
        weights1[45368] <= 16'b0000000000000011;
        weights1[45369] <= 16'b1111111111111010;
        weights1[45370] <= 16'b0000000000001101;
        weights1[45371] <= 16'b0000000000000010;
        weights1[45372] <= 16'b0000000000001000;
        weights1[45373] <= 16'b1111111111011110;
        weights1[45374] <= 16'b1111111111110000;
        weights1[45375] <= 16'b0000000000000110;
        weights1[45376] <= 16'b1111111111110000;
        weights1[45377] <= 16'b1111111111111111;
        weights1[45378] <= 16'b0000000000001000;
        weights1[45379] <= 16'b1111111111110010;
        weights1[45380] <= 16'b0000000000000000;
        weights1[45381] <= 16'b0000000000010101;
        weights1[45382] <= 16'b1111111111101111;
        weights1[45383] <= 16'b1111111111110011;
        weights1[45384] <= 16'b1111111111101011;
        weights1[45385] <= 16'b1111111111110001;
        weights1[45386] <= 16'b1111111111111000;
        weights1[45387] <= 16'b1111111111101011;
        weights1[45388] <= 16'b0000000000000000;
        weights1[45389] <= 16'b0000000000000000;
        weights1[45390] <= 16'b0000000000001000;
        weights1[45391] <= 16'b0000000000000010;
        weights1[45392] <= 16'b0000000000000000;
        weights1[45393] <= 16'b1111111111110000;
        weights1[45394] <= 16'b1111111111111111;
        weights1[45395] <= 16'b0000000000001101;
        weights1[45396] <= 16'b1111111111110010;
        weights1[45397] <= 16'b0000000000001010;
        weights1[45398] <= 16'b1111111111110000;
        weights1[45399] <= 16'b1111111111101111;
        weights1[45400] <= 16'b0000000000000110;
        weights1[45401] <= 16'b1111111111111011;
        weights1[45402] <= 16'b0000000000001010;
        weights1[45403] <= 16'b1111111111110100;
        weights1[45404] <= 16'b1111111111110100;
        weights1[45405] <= 16'b0000000000000001;
        weights1[45406] <= 16'b1111111111111100;
        weights1[45407] <= 16'b1111111111011010;
        weights1[45408] <= 16'b1111111111100110;
        weights1[45409] <= 16'b1111111111100010;
        weights1[45410] <= 16'b1111111111101001;
        weights1[45411] <= 16'b1111111111100100;
        weights1[45412] <= 16'b1111111111101100;
        weights1[45413] <= 16'b1111111111101100;
        weights1[45414] <= 16'b1111111111110111;
        weights1[45415] <= 16'b1111111111110101;
        weights1[45416] <= 16'b0000000000000010;
        weights1[45417] <= 16'b1111111111111010;
        weights1[45418] <= 16'b1111111111111101;
        weights1[45419] <= 16'b1111111111111110;
        weights1[45420] <= 16'b0000000000001100;
        weights1[45421] <= 16'b0000000000000000;
        weights1[45422] <= 16'b1111111111111100;
        weights1[45423] <= 16'b1111111111111111;
        weights1[45424] <= 16'b1111111111111010;
        weights1[45425] <= 16'b1111111111111001;
        weights1[45426] <= 16'b1111111111110110;
        weights1[45427] <= 16'b0000000000000100;
        weights1[45428] <= 16'b1111111111110100;
        weights1[45429] <= 16'b1111111111111011;
        weights1[45430] <= 16'b1111111111101101;
        weights1[45431] <= 16'b0000000000001000;
        weights1[45432] <= 16'b1111111111111001;
        weights1[45433] <= 16'b1111111111101010;
        weights1[45434] <= 16'b1111111111110100;
        weights1[45435] <= 16'b1111111111110001;
        weights1[45436] <= 16'b1111111111110010;
        weights1[45437] <= 16'b1111111111110000;
        weights1[45438] <= 16'b1111111111101011;
        weights1[45439] <= 16'b1111111111101110;
        weights1[45440] <= 16'b1111111111101001;
        weights1[45441] <= 16'b1111111111101000;
        weights1[45442] <= 16'b1111111111110010;
        weights1[45443] <= 16'b1111111111111001;
        weights1[45444] <= 16'b1111111111111110;
        weights1[45445] <= 16'b1111111111111110;
        weights1[45446] <= 16'b1111111111111001;
        weights1[45447] <= 16'b1111111111111110;
        weights1[45448] <= 16'b1111111111110100;
        weights1[45449] <= 16'b0000000000000011;
        weights1[45450] <= 16'b0000000000000000;
        weights1[45451] <= 16'b1111111111101010;
        weights1[45452] <= 16'b1111111111101111;
        weights1[45453] <= 16'b1111111111100000;
        weights1[45454] <= 16'b1111111111111011;
        weights1[45455] <= 16'b1111111111110100;
        weights1[45456] <= 16'b1111111111111001;
        weights1[45457] <= 16'b1111111111111011;
        weights1[45458] <= 16'b1111111111110001;
        weights1[45459] <= 16'b1111111111101001;
        weights1[45460] <= 16'b1111111111111010;
        weights1[45461] <= 16'b1111111111101101;
        weights1[45462] <= 16'b1111111111101101;
        weights1[45463] <= 16'b1111111111101101;
        weights1[45464] <= 16'b1111111111100011;
        weights1[45465] <= 16'b1111111111101010;
        weights1[45466] <= 16'b1111111111011101;
        weights1[45467] <= 16'b1111111111110000;
        weights1[45468] <= 16'b1111111111101101;
        weights1[45469] <= 16'b1111111111110010;
        weights1[45470] <= 16'b1111111111110111;
        weights1[45471] <= 16'b1111111111111110;
        weights1[45472] <= 16'b0000000000000000;
        weights1[45473] <= 16'b0000000000000000;
        weights1[45474] <= 16'b0000000000000011;
        weights1[45475] <= 16'b0000000000000011;
        weights1[45476] <= 16'b1111111111111101;
        weights1[45477] <= 16'b0000000000000000;
        weights1[45478] <= 16'b0000000000000000;
        weights1[45479] <= 16'b0000000000010100;
        weights1[45480] <= 16'b0000000000011111;
        weights1[45481] <= 16'b0000000000011100;
        weights1[45482] <= 16'b0000000000011111;
        weights1[45483] <= 16'b0000000000010110;
        weights1[45484] <= 16'b1111111111111101;
        weights1[45485] <= 16'b1111111111111001;
        weights1[45486] <= 16'b0000000000010110;
        weights1[45487] <= 16'b0000000000001111;
        weights1[45488] <= 16'b1111111111111111;
        weights1[45489] <= 16'b1111111111101001;
        weights1[45490] <= 16'b0000000000001010;
        weights1[45491] <= 16'b1111111111111110;
        weights1[45492] <= 16'b0000000000000101;
        weights1[45493] <= 16'b1111111111111110;
        weights1[45494] <= 16'b1111111111111001;
        weights1[45495] <= 16'b1111111111111100;
        weights1[45496] <= 16'b0000000000000001;
        weights1[45497] <= 16'b0000000000000010;
        weights1[45498] <= 16'b0000000000000000;
        weights1[45499] <= 16'b0000000000000000;
        weights1[45500] <= 16'b0000000000000001;
        weights1[45501] <= 16'b0000000000000001;
        weights1[45502] <= 16'b0000000000000000;
        weights1[45503] <= 16'b0000000000000101;
        weights1[45504] <= 16'b0000000000000011;
        weights1[45505] <= 16'b1111111111111010;
        weights1[45506] <= 16'b0000000000010000;
        weights1[45507] <= 16'b0000000000001110;
        weights1[45508] <= 16'b0000000000011110;
        weights1[45509] <= 16'b0000000000100000;
        weights1[45510] <= 16'b0000000000010111;
        weights1[45511] <= 16'b0000000000100111;
        weights1[45512] <= 16'b0000000000010001;
        weights1[45513] <= 16'b0000000000000100;
        weights1[45514] <= 16'b0000000000010000;
        weights1[45515] <= 16'b0000000000000011;
        weights1[45516] <= 16'b1111111111110100;
        weights1[45517] <= 16'b1111111111111111;
        weights1[45518] <= 16'b0000000000001011;
        weights1[45519] <= 16'b1111111111111110;
        weights1[45520] <= 16'b0000000000001011;
        weights1[45521] <= 16'b0000000000000010;
        weights1[45522] <= 16'b0000000000000011;
        weights1[45523] <= 16'b0000000000000100;
        weights1[45524] <= 16'b0000000000000110;
        weights1[45525] <= 16'b0000000000000010;
        weights1[45526] <= 16'b0000000000000010;
        weights1[45527] <= 16'b0000000000000001;
        weights1[45528] <= 16'b0000000000000011;
        weights1[45529] <= 16'b0000000000000011;
        weights1[45530] <= 16'b0000000000000101;
        weights1[45531] <= 16'b0000000000000011;
        weights1[45532] <= 16'b1111111111111111;
        weights1[45533] <= 16'b0000000000000100;
        weights1[45534] <= 16'b0000000000001110;
        weights1[45535] <= 16'b0000000000010111;
        weights1[45536] <= 16'b0000000000010000;
        weights1[45537] <= 16'b0000000000001110;
        weights1[45538] <= 16'b0000000000011010;
        weights1[45539] <= 16'b0000000000001011;
        weights1[45540] <= 16'b0000000000001001;
        weights1[45541] <= 16'b0000000000001010;
        weights1[45542] <= 16'b0000000000000000;
        weights1[45543] <= 16'b0000000000001111;
        weights1[45544] <= 16'b0000000000001100;
        weights1[45545] <= 16'b1111111111111100;
        weights1[45546] <= 16'b1111111111101111;
        weights1[45547] <= 16'b0000000000001101;
        weights1[45548] <= 16'b0000000000010000;
        weights1[45549] <= 16'b0000000000000001;
        weights1[45550] <= 16'b0000000000001100;
        weights1[45551] <= 16'b1111111111111111;
        weights1[45552] <= 16'b0000000000010001;
        weights1[45553] <= 16'b0000000000000010;
        weights1[45554] <= 16'b0000000000000011;
        weights1[45555] <= 16'b0000000000000010;
        weights1[45556] <= 16'b0000000000000111;
        weights1[45557] <= 16'b0000000000000010;
        weights1[45558] <= 16'b0000000000001000;
        weights1[45559] <= 16'b0000000000001000;
        weights1[45560] <= 16'b1111111111111100;
        weights1[45561] <= 16'b0000000000000100;
        weights1[45562] <= 16'b0000000000010100;
        weights1[45563] <= 16'b0000000000010110;
        weights1[45564] <= 16'b0000000000011001;
        weights1[45565] <= 16'b0000000000010111;
        weights1[45566] <= 16'b0000000000011000;
        weights1[45567] <= 16'b0000000000010101;
        weights1[45568] <= 16'b0000000000011000;
        weights1[45569] <= 16'b0000000000000100;
        weights1[45570] <= 16'b0000000000001100;
        weights1[45571] <= 16'b0000000000010111;
        weights1[45572] <= 16'b0000000000001000;
        weights1[45573] <= 16'b0000000000011011;
        weights1[45574] <= 16'b0000000000010011;
        weights1[45575] <= 16'b0000000000010000;
        weights1[45576] <= 16'b0000000000010111;
        weights1[45577] <= 16'b0000000000001111;
        weights1[45578] <= 16'b0000000000011110;
        weights1[45579] <= 16'b0000000000011111;
        weights1[45580] <= 16'b0000000000100000;
        weights1[45581] <= 16'b0000000000010010;
        weights1[45582] <= 16'b0000000000010000;
        weights1[45583] <= 16'b1111111111111110;
        weights1[45584] <= 16'b0000000000001001;
        weights1[45585] <= 16'b0000000000000111;
        weights1[45586] <= 16'b0000000000001001;
        weights1[45587] <= 16'b0000000000000000;
        weights1[45588] <= 16'b0000000000010001;
        weights1[45589] <= 16'b0000000000000001;
        weights1[45590] <= 16'b0000000000001111;
        weights1[45591] <= 16'b0000000000100011;
        weights1[45592] <= 16'b0000000000100001;
        weights1[45593] <= 16'b1111111111111100;
        weights1[45594] <= 16'b0000000000010100;
        weights1[45595] <= 16'b0000000000010010;
        weights1[45596] <= 16'b0000000000001000;
        weights1[45597] <= 16'b0000000000011001;
        weights1[45598] <= 16'b0000000000010010;
        weights1[45599] <= 16'b0000000000000001;
        weights1[45600] <= 16'b0000000000010100;
        weights1[45601] <= 16'b0000000000011010;
        weights1[45602] <= 16'b0000000000010011;
        weights1[45603] <= 16'b0000000000001011;
        weights1[45604] <= 16'b0000000000000010;
        weights1[45605] <= 16'b1111111111111001;
        weights1[45606] <= 16'b0000000000000100;
        weights1[45607] <= 16'b0000000000000110;
        weights1[45608] <= 16'b0000000000011000;
        weights1[45609] <= 16'b0000000000010100;
        weights1[45610] <= 16'b0000000000010000;
        weights1[45611] <= 16'b0000000000001010;
        weights1[45612] <= 16'b0000000000000110;
        weights1[45613] <= 16'b0000000000001101;
        weights1[45614] <= 16'b0000000000001011;
        weights1[45615] <= 16'b0000000000000100;
        weights1[45616] <= 16'b0000000000000000;
        weights1[45617] <= 16'b0000000000001110;
        weights1[45618] <= 16'b0000000000011010;
        weights1[45619] <= 16'b0000000000011100;
        weights1[45620] <= 16'b1111111111111011;
        weights1[45621] <= 16'b0000000000100110;
        weights1[45622] <= 16'b0000000000000100;
        weights1[45623] <= 16'b0000000000000001;
        weights1[45624] <= 16'b0000000000001001;
        weights1[45625] <= 16'b0000000000001110;
        weights1[45626] <= 16'b0000000000001111;
        weights1[45627] <= 16'b0000000000000011;
        weights1[45628] <= 16'b0000000000101010;
        weights1[45629] <= 16'b0000000000010101;
        weights1[45630] <= 16'b0000000000001101;
        weights1[45631] <= 16'b0000000000000100;
        weights1[45632] <= 16'b0000000000100100;
        weights1[45633] <= 16'b0000000000010000;
        weights1[45634] <= 16'b0000000000011010;
        weights1[45635] <= 16'b0000000000011100;
        weights1[45636] <= 16'b0000000000101011;
        weights1[45637] <= 16'b0000000000100100;
        weights1[45638] <= 16'b0000000000001010;
        weights1[45639] <= 16'b0000000000001101;
        weights1[45640] <= 16'b0000000000000101;
        weights1[45641] <= 16'b1111111111111111;
        weights1[45642] <= 16'b0000000000000000;
        weights1[45643] <= 16'b1111111111111010;
        weights1[45644] <= 16'b1111111111101101;
        weights1[45645] <= 16'b0000000000010011;
        weights1[45646] <= 16'b0000000000010011;
        weights1[45647] <= 16'b0000000000001100;
        weights1[45648] <= 16'b0000000000010011;
        weights1[45649] <= 16'b1111111111111001;
        weights1[45650] <= 16'b0000000000001001;
        weights1[45651] <= 16'b0000000000011100;
        weights1[45652] <= 16'b0000000000100001;
        weights1[45653] <= 16'b0000000000000011;
        weights1[45654] <= 16'b0000000000000111;
        weights1[45655] <= 16'b0000000000011110;
        weights1[45656] <= 16'b0000000000010100;
        weights1[45657] <= 16'b0000000000001011;
        weights1[45658] <= 16'b0000000000101000;
        weights1[45659] <= 16'b0000000000011111;
        weights1[45660] <= 16'b0000000000100111;
        weights1[45661] <= 16'b0000000000011111;
        weights1[45662] <= 16'b0000000000101110;
        weights1[45663] <= 16'b0000000000011101;
        weights1[45664] <= 16'b0000000000101100;
        weights1[45665] <= 16'b0000000000011111;
        weights1[45666] <= 16'b0000000000001010;
        weights1[45667] <= 16'b0000000000000100;
        weights1[45668] <= 16'b1111111111111111;
        weights1[45669] <= 16'b1111111111110111;
        weights1[45670] <= 16'b1111111111101011;
        weights1[45671] <= 16'b1111111111101110;
        weights1[45672] <= 16'b1111111111110101;
        weights1[45673] <= 16'b0000000000000011;
        weights1[45674] <= 16'b0000000000011110;
        weights1[45675] <= 16'b0000000000011111;
        weights1[45676] <= 16'b0000000000011000;
        weights1[45677] <= 16'b0000000000010000;
        weights1[45678] <= 16'b0000000000100111;
        weights1[45679] <= 16'b0000000000001111;
        weights1[45680] <= 16'b0000000000100010;
        weights1[45681] <= 16'b1111111111110101;
        weights1[45682] <= 16'b0000000000011010;
        weights1[45683] <= 16'b0000000000000000;
        weights1[45684] <= 16'b0000000000000100;
        weights1[45685] <= 16'b0000000000010101;
        weights1[45686] <= 16'b0000000000011010;
        weights1[45687] <= 16'b0000000000001101;
        weights1[45688] <= 16'b0000000000011011;
        weights1[45689] <= 16'b0000000000000110;
        weights1[45690] <= 16'b0000000000000101;
        weights1[45691] <= 16'b0000000001000011;
        weights1[45692] <= 16'b0000000000011001;
        weights1[45693] <= 16'b0000000000100000;
        weights1[45694] <= 16'b0000000000000110;
        weights1[45695] <= 16'b0000000000000111;
        weights1[45696] <= 16'b1111111111111000;
        weights1[45697] <= 16'b1111111111101101;
        weights1[45698] <= 16'b1111111111100101;
        weights1[45699] <= 16'b1111111111011101;
        weights1[45700] <= 16'b1111111111010110;
        weights1[45701] <= 16'b1111111111111110;
        weights1[45702] <= 16'b0000000000101101;
        weights1[45703] <= 16'b0000000000100010;
        weights1[45704] <= 16'b0000000000100110;
        weights1[45705] <= 16'b0000000000010001;
        weights1[45706] <= 16'b0000000000011001;
        weights1[45707] <= 16'b0000000000011110;
        weights1[45708] <= 16'b0000000000001101;
        weights1[45709] <= 16'b0000000000001011;
        weights1[45710] <= 16'b0000000000011001;
        weights1[45711] <= 16'b0000000000010110;
        weights1[45712] <= 16'b0000000000010000;
        weights1[45713] <= 16'b0000000000000111;
        weights1[45714] <= 16'b0000000000001111;
        weights1[45715] <= 16'b0000000000011111;
        weights1[45716] <= 16'b0000000000011111;
        weights1[45717] <= 16'b0000000000011111;
        weights1[45718] <= 16'b0000000000100011;
        weights1[45719] <= 16'b0000000000101000;
        weights1[45720] <= 16'b0000000000100011;
        weights1[45721] <= 16'b0000000000000001;
        weights1[45722] <= 16'b1111111111111000;
        weights1[45723] <= 16'b1111111111111111;
        weights1[45724] <= 16'b1111111111110010;
        weights1[45725] <= 16'b1111111111100010;
        weights1[45726] <= 16'b1111111111011110;
        weights1[45727] <= 16'b1111111111000110;
        weights1[45728] <= 16'b1111111111000100;
        weights1[45729] <= 16'b1111111111011001;
        weights1[45730] <= 16'b0000000000001101;
        weights1[45731] <= 16'b0000000000011001;
        weights1[45732] <= 16'b0000000000010001;
        weights1[45733] <= 16'b0000000000110011;
        weights1[45734] <= 16'b0000000000101100;
        weights1[45735] <= 16'b0000000000111011;
        weights1[45736] <= 16'b0000000000010010;
        weights1[45737] <= 16'b0000000000111000;
        weights1[45738] <= 16'b0000000000101100;
        weights1[45739] <= 16'b0000000000001100;
        weights1[45740] <= 16'b0000000000001101;
        weights1[45741] <= 16'b0000000000001111;
        weights1[45742] <= 16'b0000000000000101;
        weights1[45743] <= 16'b0000000000000110;
        weights1[45744] <= 16'b0000000000000101;
        weights1[45745] <= 16'b0000000000101011;
        weights1[45746] <= 16'b0000000000100001;
        weights1[45747] <= 16'b0000000000001001;
        weights1[45748] <= 16'b1111111111110011;
        weights1[45749] <= 16'b1111111111101100;
        weights1[45750] <= 16'b1111111111110001;
        weights1[45751] <= 16'b1111111111110011;
        weights1[45752] <= 16'b1111111111101010;
        weights1[45753] <= 16'b1111111111011101;
        weights1[45754] <= 16'b1111111111010100;
        weights1[45755] <= 16'b1111111111000010;
        weights1[45756] <= 16'b1111111110111010;
        weights1[45757] <= 16'b1111111110100010;
        weights1[45758] <= 16'b1111111111001111;
        weights1[45759] <= 16'b1111111111111111;
        weights1[45760] <= 16'b0000000000011000;
        weights1[45761] <= 16'b0000000000010100;
        weights1[45762] <= 16'b0000000000011011;
        weights1[45763] <= 16'b0000000000110001;
        weights1[45764] <= 16'b0000000000110000;
        weights1[45765] <= 16'b0000000000010010;
        weights1[45766] <= 16'b0000000000011100;
        weights1[45767] <= 16'b0000000000100010;
        weights1[45768] <= 16'b0000000000101001;
        weights1[45769] <= 16'b1111111111111101;
        weights1[45770] <= 16'b0000000000001110;
        weights1[45771] <= 16'b0000000000001001;
        weights1[45772] <= 16'b0000000000111011;
        weights1[45773] <= 16'b0000000001000000;
        weights1[45774] <= 16'b0000000000110010;
        weights1[45775] <= 16'b1111111111110010;
        weights1[45776] <= 16'b1111111111011000;
        weights1[45777] <= 16'b1111111111100110;
        weights1[45778] <= 16'b1111111111100000;
        weights1[45779] <= 16'b1111111111100101;
        weights1[45780] <= 16'b1111111111100111;
        weights1[45781] <= 16'b1111111111011100;
        weights1[45782] <= 16'b1111111111001111;
        weights1[45783] <= 16'b1111111111001110;
        weights1[45784] <= 16'b1111111110111001;
        weights1[45785] <= 16'b1111111110001010;
        weights1[45786] <= 16'b1111111110010001;
        weights1[45787] <= 16'b1111111111011000;
        weights1[45788] <= 16'b1111111111101010;
        weights1[45789] <= 16'b0000000000000110;
        weights1[45790] <= 16'b0000000000011111;
        weights1[45791] <= 16'b0000000000101110;
        weights1[45792] <= 16'b0000000000111101;
        weights1[45793] <= 16'b0000000000011100;
        weights1[45794] <= 16'b0000000000110000;
        weights1[45795] <= 16'b0000000000100101;
        weights1[45796] <= 16'b0000000000100101;
        weights1[45797] <= 16'b0000000000100001;
        weights1[45798] <= 16'b0000000000101000;
        weights1[45799] <= 16'b0000000000010000;
        weights1[45800] <= 16'b0000000000000010;
        weights1[45801] <= 16'b0000000000000001;
        weights1[45802] <= 16'b1111111111011100;
        weights1[45803] <= 16'b1111111111010000;
        weights1[45804] <= 16'b1111111111001000;
        weights1[45805] <= 16'b1111111111011110;
        weights1[45806] <= 16'b1111111111100111;
        weights1[45807] <= 16'b1111111111100011;
        weights1[45808] <= 16'b1111111111100111;
        weights1[45809] <= 16'b1111111111100100;
        weights1[45810] <= 16'b1111111111100001;
        weights1[45811] <= 16'b1111111111011010;
        weights1[45812] <= 16'b1111111111010100;
        weights1[45813] <= 16'b1111111110110011;
        weights1[45814] <= 16'b1111111110010100;
        weights1[45815] <= 16'b1111111110010110;
        weights1[45816] <= 16'b1111111110110001;
        weights1[45817] <= 16'b1111111111111100;
        weights1[45818] <= 16'b1111111111111111;
        weights1[45819] <= 16'b0000000000101010;
        weights1[45820] <= 16'b0000000000111000;
        weights1[45821] <= 16'b0000000000101111;
        weights1[45822] <= 16'b0000000000011111;
        weights1[45823] <= 16'b0000000000011001;
        weights1[45824] <= 16'b0000000000011001;
        weights1[45825] <= 16'b0000000000011010;
        weights1[45826] <= 16'b0000000000000111;
        weights1[45827] <= 16'b1111111111110010;
        weights1[45828] <= 16'b1111111111100000;
        weights1[45829] <= 16'b1111111111000010;
        weights1[45830] <= 16'b1111111110010111;
        weights1[45831] <= 16'b1111111110100011;
        weights1[45832] <= 16'b1111111110111001;
        weights1[45833] <= 16'b1111111111010110;
        weights1[45834] <= 16'b1111111111010111;
        weights1[45835] <= 16'b1111111111100000;
        weights1[45836] <= 16'b1111111111110011;
        weights1[45837] <= 16'b1111111111101111;
        weights1[45838] <= 16'b1111111111110110;
        weights1[45839] <= 16'b1111111111111001;
        weights1[45840] <= 16'b1111111111100001;
        weights1[45841] <= 16'b1111111111011110;
        weights1[45842] <= 16'b1111111110111110;
        weights1[45843] <= 16'b1111111110101110;
        weights1[45844] <= 16'b1111111110100001;
        weights1[45845] <= 16'b1111111110101111;
        weights1[45846] <= 16'b1111111111001010;
        weights1[45847] <= 16'b1111111111100100;
        weights1[45848] <= 16'b0000000000110001;
        weights1[45849] <= 16'b0000000000110101;
        weights1[45850] <= 16'b0000000000100111;
        weights1[45851] <= 16'b0000000000101010;
        weights1[45852] <= 16'b0000000000001000;
        weights1[45853] <= 16'b1111111111110110;
        weights1[45854] <= 16'b1111111111101110;
        weights1[45855] <= 16'b1111111111100100;
        weights1[45856] <= 16'b1111111110010110;
        weights1[45857] <= 16'b1111111101111011;
        weights1[45858] <= 16'b1111111110010101;
        weights1[45859] <= 16'b1111111110110100;
        weights1[45860] <= 16'b1111111111001100;
        weights1[45861] <= 16'b1111111111011100;
        weights1[45862] <= 16'b1111111111101000;
        weights1[45863] <= 16'b1111111111101100;
        weights1[45864] <= 16'b0000000000000011;
        weights1[45865] <= 16'b0000000000000000;
        weights1[45866] <= 16'b1111111111111110;
        weights1[45867] <= 16'b1111111111111000;
        weights1[45868] <= 16'b0000000000001001;
        weights1[45869] <= 16'b1111111111110001;
        weights1[45870] <= 16'b1111111111111001;
        weights1[45871] <= 16'b1111111111000010;
        weights1[45872] <= 16'b1111111110111110;
        weights1[45873] <= 16'b1111111110110101;
        weights1[45874] <= 16'b1111111111000001;
        weights1[45875] <= 16'b1111111110111111;
        weights1[45876] <= 16'b1111111111011100;
        weights1[45877] <= 16'b0000000000001011;
        weights1[45878] <= 16'b0000000000000000;
        weights1[45879] <= 16'b0000000000000000;
        weights1[45880] <= 16'b1111111111111101;
        weights1[45881] <= 16'b1111111111101110;
        weights1[45882] <= 16'b1111111111010011;
        weights1[45883] <= 16'b1111111111010011;
        weights1[45884] <= 16'b1111111110111010;
        weights1[45885] <= 16'b1111111110101001;
        weights1[45886] <= 16'b1111111111000001;
        weights1[45887] <= 16'b1111111110111101;
        weights1[45888] <= 16'b1111111111001100;
        weights1[45889] <= 16'b1111111111100111;
        weights1[45890] <= 16'b1111111111110010;
        weights1[45891] <= 16'b1111111111110001;
        weights1[45892] <= 16'b0000000000000000;
        weights1[45893] <= 16'b1111111111111000;
        weights1[45894] <= 16'b1111111111110011;
        weights1[45895] <= 16'b1111111111111010;
        weights1[45896] <= 16'b0000000000001110;
        weights1[45897] <= 16'b0000000000001110;
        weights1[45898] <= 16'b1111111111110101;
        weights1[45899] <= 16'b1111111111111110;
        weights1[45900] <= 16'b1111111111011111;
        weights1[45901] <= 16'b1111111111001010;
        weights1[45902] <= 16'b1111111110110110;
        weights1[45903] <= 16'b1111111110101110;
        weights1[45904] <= 16'b1111111111000111;
        weights1[45905] <= 16'b1111111111110101;
        weights1[45906] <= 16'b1111111111101001;
        weights1[45907] <= 16'b1111111111011111;
        weights1[45908] <= 16'b1111111111101000;
        weights1[45909] <= 16'b1111111111010100;
        weights1[45910] <= 16'b1111111111101100;
        weights1[45911] <= 16'b1111111111011110;
        weights1[45912] <= 16'b1111111111110101;
        weights1[45913] <= 16'b0000000000000010;
        weights1[45914] <= 16'b1111111111010010;
        weights1[45915] <= 16'b1111111111000111;
        weights1[45916] <= 16'b1111111111001110;
        weights1[45917] <= 16'b1111111111101100;
        weights1[45918] <= 16'b1111111111101111;
        weights1[45919] <= 16'b1111111111101111;
        weights1[45920] <= 16'b0000000000000101;
        weights1[45921] <= 16'b1111111111110101;
        weights1[45922] <= 16'b0000000000000010;
        weights1[45923] <= 16'b1111111111111001;
        weights1[45924] <= 16'b0000000000000100;
        weights1[45925] <= 16'b0000000000010011;
        weights1[45926] <= 16'b0000000000000111;
        weights1[45927] <= 16'b0000000000010001;
        weights1[45928] <= 16'b1111111111110110;
        weights1[45929] <= 16'b1111111111110010;
        weights1[45930] <= 16'b1111111111011110;
        weights1[45931] <= 16'b1111111111100011;
        weights1[45932] <= 16'b1111111110111100;
        weights1[45933] <= 16'b1111111110111101;
        weights1[45934] <= 16'b1111111111101000;
        weights1[45935] <= 16'b1111111111101110;
        weights1[45936] <= 16'b1111111111011100;
        weights1[45937] <= 16'b1111111111100110;
        weights1[45938] <= 16'b1111111111011100;
        weights1[45939] <= 16'b1111111111111100;
        weights1[45940] <= 16'b0000000000011000;
        weights1[45941] <= 16'b1111111111111000;
        weights1[45942] <= 16'b1111111110111101;
        weights1[45943] <= 16'b1111111110111010;
        weights1[45944] <= 16'b1111111111010100;
        weights1[45945] <= 16'b1111111111100111;
        weights1[45946] <= 16'b1111111111110010;
        weights1[45947] <= 16'b1111111111110110;
        weights1[45948] <= 16'b0000000000000000;
        weights1[45949] <= 16'b0000000000000011;
        weights1[45950] <= 16'b0000000000001101;
        weights1[45951] <= 16'b0000000000001100;
        weights1[45952] <= 16'b0000000000000000;
        weights1[45953] <= 16'b1111111111110111;
        weights1[45954] <= 16'b0000000000001101;
        weights1[45955] <= 16'b0000000000000010;
        weights1[45956] <= 16'b0000000000000011;
        weights1[45957] <= 16'b0000000000001010;
        weights1[45958] <= 16'b1111111111100101;
        weights1[45959] <= 16'b1111111111111001;
        weights1[45960] <= 16'b1111111111011101;
        weights1[45961] <= 16'b1111111111010000;
        weights1[45962] <= 16'b1111111111101100;
        weights1[45963] <= 16'b1111111111101000;
        weights1[45964] <= 16'b0000000000000110;
        weights1[45965] <= 16'b0000000000000101;
        weights1[45966] <= 16'b1111111111111100;
        weights1[45967] <= 16'b1111111111111010;
        weights1[45968] <= 16'b0000000000000001;
        weights1[45969] <= 16'b0000000000000111;
        weights1[45970] <= 16'b1111111111001110;
        weights1[45971] <= 16'b1111111111001001;
        weights1[45972] <= 16'b1111111111011011;
        weights1[45973] <= 16'b1111111111100010;
        weights1[45974] <= 16'b1111111111111000;
        weights1[45975] <= 16'b1111111111110101;
        weights1[45976] <= 16'b1111111111111110;
        weights1[45977] <= 16'b1111111111111011;
        weights1[45978] <= 16'b1111111111111101;
        weights1[45979] <= 16'b1111111111111010;
        weights1[45980] <= 16'b1111111111110111;
        weights1[45981] <= 16'b1111111111111000;
        weights1[45982] <= 16'b1111111111110111;
        weights1[45983] <= 16'b0000000000010000;
        weights1[45984] <= 16'b0000000000000101;
        weights1[45985] <= 16'b1111111111101101;
        weights1[45986] <= 16'b1111111111111101;
        weights1[45987] <= 16'b1111111111111011;
        weights1[45988] <= 16'b1111111111010001;
        weights1[45989] <= 16'b1111111111110000;
        weights1[45990] <= 16'b1111111111100111;
        weights1[45991] <= 16'b1111111111101011;
        weights1[45992] <= 16'b1111111111111001;
        weights1[45993] <= 16'b1111111111110111;
        weights1[45994] <= 16'b0000000000001000;
        weights1[45995] <= 16'b0000000000010111;
        weights1[45996] <= 16'b0000000000010110;
        weights1[45997] <= 16'b0000000000001111;
        weights1[45998] <= 16'b1111111111000110;
        weights1[45999] <= 16'b1111111111001111;
        weights1[46000] <= 16'b1111111111010100;
        weights1[46001] <= 16'b1111111111100010;
        weights1[46002] <= 16'b1111111111111001;
        weights1[46003] <= 16'b1111111111110111;
        weights1[46004] <= 16'b1111111111110111;
        weights1[46005] <= 16'b1111111111110001;
        weights1[46006] <= 16'b1111111111101101;
        weights1[46007] <= 16'b1111111111100101;
        weights1[46008] <= 16'b0000000000001101;
        weights1[46009] <= 16'b1111111111110110;
        weights1[46010] <= 16'b0000000000010101;
        weights1[46011] <= 16'b0000000000000011;
        weights1[46012] <= 16'b0000000000010001;
        weights1[46013] <= 16'b1111111111101100;
        weights1[46014] <= 16'b1111111111101000;
        weights1[46015] <= 16'b1111111111111000;
        weights1[46016] <= 16'b0000000000000011;
        weights1[46017] <= 16'b0000000000000100;
        weights1[46018] <= 16'b1111111111111111;
        weights1[46019] <= 16'b1111111111101000;
        weights1[46020] <= 16'b1111111111110100;
        weights1[46021] <= 16'b1111111111111011;
        weights1[46022] <= 16'b1111111111111001;
        weights1[46023] <= 16'b0000000000001010;
        weights1[46024] <= 16'b0000000000011100;
        weights1[46025] <= 16'b1111111111101000;
        weights1[46026] <= 16'b1111111111001101;
        weights1[46027] <= 16'b1111111111000111;
        weights1[46028] <= 16'b1111111111101000;
        weights1[46029] <= 16'b1111111111101011;
        weights1[46030] <= 16'b1111111111110100;
        weights1[46031] <= 16'b1111111111111000;
        weights1[46032] <= 16'b1111111111111011;
        weights1[46033] <= 16'b1111111111110101;
        weights1[46034] <= 16'b1111111111110110;
        weights1[46035] <= 16'b1111111111100000;
        weights1[46036] <= 16'b1111111111110101;
        weights1[46037] <= 16'b1111111111101101;
        weights1[46038] <= 16'b0000000000000010;
        weights1[46039] <= 16'b1111111111110100;
        weights1[46040] <= 16'b1111111111111110;
        weights1[46041] <= 16'b1111111111111001;
        weights1[46042] <= 16'b0000000000000101;
        weights1[46043] <= 16'b1111111111111111;
        weights1[46044] <= 16'b1111111111011000;
        weights1[46045] <= 16'b1111111111110110;
        weights1[46046] <= 16'b1111111111111001;
        weights1[46047] <= 16'b1111111111101101;
        weights1[46048] <= 16'b1111111111101010;
        weights1[46049] <= 16'b0000000000001000;
        weights1[46050] <= 16'b1111111111110100;
        weights1[46051] <= 16'b1111111111111001;
        weights1[46052] <= 16'b0000000000000101;
        weights1[46053] <= 16'b1111111111110000;
        weights1[46054] <= 16'b1111111110111110;
        weights1[46055] <= 16'b1111111111011010;
        weights1[46056] <= 16'b1111111111101111;
        weights1[46057] <= 16'b1111111111110110;
        weights1[46058] <= 16'b1111111111111000;
        weights1[46059] <= 16'b1111111111110110;
        weights1[46060] <= 16'b0000000000000010;
        weights1[46061] <= 16'b1111111111111100;
        weights1[46062] <= 16'b1111111111111010;
        weights1[46063] <= 16'b1111111111100001;
        weights1[46064] <= 16'b1111111111111010;
        weights1[46065] <= 16'b1111111111100110;
        weights1[46066] <= 16'b1111111111111000;
        weights1[46067] <= 16'b1111111111101010;
        weights1[46068] <= 16'b0000000000000111;
        weights1[46069] <= 16'b1111111111110110;
        weights1[46070] <= 16'b1111111111111101;
        weights1[46071] <= 16'b0000000000000000;
        weights1[46072] <= 16'b1111111111111000;
        weights1[46073] <= 16'b1111111111110111;
        weights1[46074] <= 16'b1111111111110100;
        weights1[46075] <= 16'b0000000000000001;
        weights1[46076] <= 16'b1111111111101001;
        weights1[46077] <= 16'b1111111111111001;
        weights1[46078] <= 16'b0000000000000001;
        weights1[46079] <= 16'b1111111111100011;
        weights1[46080] <= 16'b0000000000000100;
        weights1[46081] <= 16'b1111111111000111;
        weights1[46082] <= 16'b1111111110111110;
        weights1[46083] <= 16'b1111111111010110;
        weights1[46084] <= 16'b1111111111110011;
        weights1[46085] <= 16'b1111111111110100;
        weights1[46086] <= 16'b1111111111111101;
        weights1[46087] <= 16'b1111111111111011;
        weights1[46088] <= 16'b1111111111111100;
        weights1[46089] <= 16'b1111111111111100;
        weights1[46090] <= 16'b1111111111110010;
        weights1[46091] <= 16'b1111111111101111;
        weights1[46092] <= 16'b1111111111100011;
        weights1[46093] <= 16'b1111111111111010;
        weights1[46094] <= 16'b1111111111101000;
        weights1[46095] <= 16'b1111111111110111;
        weights1[46096] <= 16'b1111111111101111;
        weights1[46097] <= 16'b1111111111100110;
        weights1[46098] <= 16'b1111111111111011;
        weights1[46099] <= 16'b1111111111111111;
        weights1[46100] <= 16'b1111111111101011;
        weights1[46101] <= 16'b0000000000000000;
        weights1[46102] <= 16'b1111111111101110;
        weights1[46103] <= 16'b0000000000000001;
        weights1[46104] <= 16'b1111111111110000;
        weights1[46105] <= 16'b0000000000010101;
        weights1[46106] <= 16'b1111111111101010;
        weights1[46107] <= 16'b1111111111010111;
        weights1[46108] <= 16'b1111111111000111;
        weights1[46109] <= 16'b1111111111001100;
        weights1[46110] <= 16'b1111111111100001;
        weights1[46111] <= 16'b1111111111101111;
        weights1[46112] <= 16'b1111111111110101;
        weights1[46113] <= 16'b1111111111111011;
        weights1[46114] <= 16'b1111111111111111;
        weights1[46115] <= 16'b1111111111111111;
        weights1[46116] <= 16'b1111111111111100;
        weights1[46117] <= 16'b1111111111111110;
        weights1[46118] <= 16'b1111111111110011;
        weights1[46119] <= 16'b1111111111111101;
        weights1[46120] <= 16'b1111111111100010;
        weights1[46121] <= 16'b1111111111100111;
        weights1[46122] <= 16'b1111111111100010;
        weights1[46123] <= 16'b1111111111101111;
        weights1[46124] <= 16'b0000000000000010;
        weights1[46125] <= 16'b1111111111110011;
        weights1[46126] <= 16'b1111111111111000;
        weights1[46127] <= 16'b1111111111111110;
        weights1[46128] <= 16'b0000000000001001;
        weights1[46129] <= 16'b0000000000000111;
        weights1[46130] <= 16'b1111111111110000;
        weights1[46131] <= 16'b1111111111111000;
        weights1[46132] <= 16'b1111111111110011;
        weights1[46133] <= 16'b0000000000000110;
        weights1[46134] <= 16'b1111111111101010;
        weights1[46135] <= 16'b1111111111100101;
        weights1[46136] <= 16'b1111111111011110;
        weights1[46137] <= 16'b1111111111010010;
        weights1[46138] <= 16'b1111111111100111;
        weights1[46139] <= 16'b1111111111111011;
        weights1[46140] <= 16'b1111111111110110;
        weights1[46141] <= 16'b1111111111111100;
        weights1[46142] <= 16'b1111111111111101;
        weights1[46143] <= 16'b0000000000000000;
        weights1[46144] <= 16'b0000000000000000;
        weights1[46145] <= 16'b1111111111111111;
        weights1[46146] <= 16'b1111111111111101;
        weights1[46147] <= 16'b1111111111111110;
        weights1[46148] <= 16'b0000000000000011;
        weights1[46149] <= 16'b1111111111110000;
        weights1[46150] <= 16'b1111111111010111;
        weights1[46151] <= 16'b0000000000010101;
        weights1[46152] <= 16'b1111111111111010;
        weights1[46153] <= 16'b1111111111111001;
        weights1[46154] <= 16'b1111111111111101;
        weights1[46155] <= 16'b1111111111100111;
        weights1[46156] <= 16'b1111111111111110;
        weights1[46157] <= 16'b0000000000010001;
        weights1[46158] <= 16'b1111111111010010;
        weights1[46159] <= 16'b0000000000010100;
        weights1[46160] <= 16'b0000000000001001;
        weights1[46161] <= 16'b1111111111101000;
        weights1[46162] <= 16'b1111111111010101;
        weights1[46163] <= 16'b1111111111100000;
        weights1[46164] <= 16'b1111111111011001;
        weights1[46165] <= 16'b1111111111100001;
        weights1[46166] <= 16'b1111111111101101;
        weights1[46167] <= 16'b0000000000000000;
        weights1[46168] <= 16'b0000000000000010;
        weights1[46169] <= 16'b0000000000000011;
        weights1[46170] <= 16'b1111111111111111;
        weights1[46171] <= 16'b1111111111111111;
        weights1[46172] <= 16'b0000000000000000;
        weights1[46173] <= 16'b1111111111111110;
        weights1[46174] <= 16'b0000000000000011;
        weights1[46175] <= 16'b0000000000000000;
        weights1[46176] <= 16'b0000000000000011;
        weights1[46177] <= 16'b1111111111110100;
        weights1[46178] <= 16'b1111111111110101;
        weights1[46179] <= 16'b1111111111101111;
        weights1[46180] <= 16'b1111111111100000;
        weights1[46181] <= 16'b1111111111101001;
        weights1[46182] <= 16'b1111111111011100;
        weights1[46183] <= 16'b1111111111010111;
        weights1[46184] <= 16'b1111111111110001;
        weights1[46185] <= 16'b1111111111111110;
        weights1[46186] <= 16'b1111111111101011;
        weights1[46187] <= 16'b1111111111101111;
        weights1[46188] <= 16'b1111111111100001;
        weights1[46189] <= 16'b1111111111100111;
        weights1[46190] <= 16'b1111111111110001;
        weights1[46191] <= 16'b1111111111101100;
        weights1[46192] <= 16'b1111111111110011;
        weights1[46193] <= 16'b1111111111111000;
        weights1[46194] <= 16'b1111111111111110;
        weights1[46195] <= 16'b0000000000000000;
        weights1[46196] <= 16'b0000000000000001;
        weights1[46197] <= 16'b0000000000000000;
        weights1[46198] <= 16'b1111111111111101;
        weights1[46199] <= 16'b1111111111111111;
        weights1[46200] <= 16'b0000000000000000;
        weights1[46201] <= 16'b1111111111111111;
        weights1[46202] <= 16'b0000000000000100;
        weights1[46203] <= 16'b0000000000001000;
        weights1[46204] <= 16'b0000000000000110;
        weights1[46205] <= 16'b0000000000000000;
        weights1[46206] <= 16'b0000000000000000;
        weights1[46207] <= 16'b1111111111111000;
        weights1[46208] <= 16'b1111111111111010;
        weights1[46209] <= 16'b1111111111101111;
        weights1[46210] <= 16'b1111111111110101;
        weights1[46211] <= 16'b1111111111100001;
        weights1[46212] <= 16'b1111111111110101;
        weights1[46213] <= 16'b1111111111111001;
        weights1[46214] <= 16'b1111111111110000;
        weights1[46215] <= 16'b1111111111110100;
        weights1[46216] <= 16'b1111111111111111;
        weights1[46217] <= 16'b1111111111110010;
        weights1[46218] <= 16'b1111111111110101;
        weights1[46219] <= 16'b1111111111111011;
        weights1[46220] <= 16'b1111111111111101;
        weights1[46221] <= 16'b1111111111111001;
        weights1[46222] <= 16'b1111111111111000;
        weights1[46223] <= 16'b1111111111111100;
        weights1[46224] <= 16'b1111111111111011;
        weights1[46225] <= 16'b1111111111111101;
        weights1[46226] <= 16'b0000000000000000;
        weights1[46227] <= 16'b0000000000000000;
        weights1[46228] <= 16'b0000000000000000;
        weights1[46229] <= 16'b0000000000000001;
        weights1[46230] <= 16'b0000000000000011;
        weights1[46231] <= 16'b0000000000000110;
        weights1[46232] <= 16'b0000000000001001;
        weights1[46233] <= 16'b0000000000000000;
        weights1[46234] <= 16'b0000000000000110;
        weights1[46235] <= 16'b0000000000001010;
        weights1[46236] <= 16'b0000000000000000;
        weights1[46237] <= 16'b0000000000000100;
        weights1[46238] <= 16'b1111111111110110;
        weights1[46239] <= 16'b1111111111111011;
        weights1[46240] <= 16'b0000000000000100;
        weights1[46241] <= 16'b1111111111110101;
        weights1[46242] <= 16'b1111111111110110;
        weights1[46243] <= 16'b1111111111111010;
        weights1[46244] <= 16'b1111111111101111;
        weights1[46245] <= 16'b1111111111101001;
        weights1[46246] <= 16'b1111111111111010;
        weights1[46247] <= 16'b1111111111111100;
        weights1[46248] <= 16'b1111111111111010;
        weights1[46249] <= 16'b1111111111111001;
        weights1[46250] <= 16'b1111111111111111;
        weights1[46251] <= 16'b1111111111111110;
        weights1[46252] <= 16'b1111111111111100;
        weights1[46253] <= 16'b1111111111111101;
        weights1[46254] <= 16'b1111111111111110;
        weights1[46255] <= 16'b0000000000000000;
        weights1[46256] <= 16'b0000000000000001;
        weights1[46257] <= 16'b0000000000000000;
        weights1[46258] <= 16'b1111111111111111;
        weights1[46259] <= 16'b1111111111111100;
        weights1[46260] <= 16'b1111111111111101;
        weights1[46261] <= 16'b1111111111111000;
        weights1[46262] <= 16'b1111111111110111;
        weights1[46263] <= 16'b1111111111110011;
        weights1[46264] <= 16'b1111111111111001;
        weights1[46265] <= 16'b1111111111111100;
        weights1[46266] <= 16'b1111111111111011;
        weights1[46267] <= 16'b1111111111110100;
        weights1[46268] <= 16'b0000000000000000;
        weights1[46269] <= 16'b1111111111111110;
        weights1[46270] <= 16'b1111111111111001;
        weights1[46271] <= 16'b0000000000000001;
        weights1[46272] <= 16'b1111111111110001;
        weights1[46273] <= 16'b0000000000001101;
        weights1[46274] <= 16'b0000000000001110;
        weights1[46275] <= 16'b0000000000010000;
        weights1[46276] <= 16'b0000000000011110;
        weights1[46277] <= 16'b0000000000001101;
        weights1[46278] <= 16'b0000000000010011;
        weights1[46279] <= 16'b0000000000001000;
        weights1[46280] <= 16'b0000000000000011;
        weights1[46281] <= 16'b0000000000000010;
        weights1[46282] <= 16'b0000000000000001;
        weights1[46283] <= 16'b0000000000000110;
        weights1[46284] <= 16'b0000000000000000;
        weights1[46285] <= 16'b1111111111111111;
        weights1[46286] <= 16'b1111111111111010;
        weights1[46287] <= 16'b1111111111111100;
        weights1[46288] <= 16'b1111111111111001;
        weights1[46289] <= 16'b0000000000001000;
        weights1[46290] <= 16'b1111111111110110;
        weights1[46291] <= 16'b1111111111111101;
        weights1[46292] <= 16'b0000000000000010;
        weights1[46293] <= 16'b1111111111111011;
        weights1[46294] <= 16'b1111111111100010;
        weights1[46295] <= 16'b0000000000000110;
        weights1[46296] <= 16'b0000000000001100;
        weights1[46297] <= 16'b0000000000010000;
        weights1[46298] <= 16'b0000000000001101;
        weights1[46299] <= 16'b0000000000000111;
        weights1[46300] <= 16'b1111111111110111;
        weights1[46301] <= 16'b0000000000010001;
        weights1[46302] <= 16'b0000000000010110;
        weights1[46303] <= 16'b0000000000001100;
        weights1[46304] <= 16'b0000000000001101;
        weights1[46305] <= 16'b0000000000011001;
        weights1[46306] <= 16'b0000000000011100;
        weights1[46307] <= 16'b0000000000001000;
        weights1[46308] <= 16'b0000000000000010;
        weights1[46309] <= 16'b0000000000001010;
        weights1[46310] <= 16'b0000000000001111;
        weights1[46311] <= 16'b0000000000000110;
        weights1[46312] <= 16'b0000000000000000;
        weights1[46313] <= 16'b1111111111111100;
        weights1[46314] <= 16'b1111111111111110;
        weights1[46315] <= 16'b0000000000000100;
        weights1[46316] <= 16'b0000000000001001;
        weights1[46317] <= 16'b0000000000001100;
        weights1[46318] <= 16'b0000000000001000;
        weights1[46319] <= 16'b1111111111111000;
        weights1[46320] <= 16'b0000000000000101;
        weights1[46321] <= 16'b0000000000000110;
        weights1[46322] <= 16'b0000000000000000;
        weights1[46323] <= 16'b0000000000000110;
        weights1[46324] <= 16'b0000000000001010;
        weights1[46325] <= 16'b0000000000000110;
        weights1[46326] <= 16'b1111111111110110;
        weights1[46327] <= 16'b1111111111110110;
        weights1[46328] <= 16'b0000000000010000;
        weights1[46329] <= 16'b0000000000010010;
        weights1[46330] <= 16'b0000000000010010;
        weights1[46331] <= 16'b0000000000011010;
        weights1[46332] <= 16'b0000000000001111;
        weights1[46333] <= 16'b0000000000010100;
        weights1[46334] <= 16'b0000000000011100;
        weights1[46335] <= 16'b0000000000100001;
        weights1[46336] <= 16'b0000000000011001;
        weights1[46337] <= 16'b0000000000100111;
        weights1[46338] <= 16'b0000000000011100;
        weights1[46339] <= 16'b0000000000001011;
        weights1[46340] <= 16'b1111111111111101;
        weights1[46341] <= 16'b1111111111110110;
        weights1[46342] <= 16'b1111111111111111;
        weights1[46343] <= 16'b0000000000001101;
        weights1[46344] <= 16'b0000000000010101;
        weights1[46345] <= 16'b0000000000011011;
        weights1[46346] <= 16'b0000000000100100;
        weights1[46347] <= 16'b0000000000010110;
        weights1[46348] <= 16'b0000000000011111;
        weights1[46349] <= 16'b0000000000011001;
        weights1[46350] <= 16'b0000000000010010;
        weights1[46351] <= 16'b0000000000010010;
        weights1[46352] <= 16'b0000000000010010;
        weights1[46353] <= 16'b0000000000010100;
        weights1[46354] <= 16'b0000000000010010;
        weights1[46355] <= 16'b0000000000010111;
        weights1[46356] <= 16'b0000000000010111;
        weights1[46357] <= 16'b0000000000011101;
        weights1[46358] <= 16'b0000000000101110;
        weights1[46359] <= 16'b0000000000001010;
        weights1[46360] <= 16'b0000000000010011;
        weights1[46361] <= 16'b0000000000101001;
        weights1[46362] <= 16'b0000000000100000;
        weights1[46363] <= 16'b0000000000011011;
        weights1[46364] <= 16'b0000000000101010;
        weights1[46365] <= 16'b0000000000100100;
        weights1[46366] <= 16'b0000000000010111;
        weights1[46367] <= 16'b0000000000010001;
        weights1[46368] <= 16'b1111111111111110;
        weights1[46369] <= 16'b1111111111111001;
        weights1[46370] <= 16'b0000000000000100;
        weights1[46371] <= 16'b0000000000010001;
        weights1[46372] <= 16'b0000000000100010;
        weights1[46373] <= 16'b0000000000100001;
        weights1[46374] <= 16'b0000000000100001;
        weights1[46375] <= 16'b0000000000100111;
        weights1[46376] <= 16'b0000000000110001;
        weights1[46377] <= 16'b0000000000111011;
        weights1[46378] <= 16'b0000000000101000;
        weights1[46379] <= 16'b0000000000100001;
        weights1[46380] <= 16'b0000000000101010;
        weights1[46381] <= 16'b0000000000100001;
        weights1[46382] <= 16'b0000000000011001;
        weights1[46383] <= 16'b0000000000001110;
        weights1[46384] <= 16'b0000000000111001;
        weights1[46385] <= 16'b0000000000010011;
        weights1[46386] <= 16'b0000000000010101;
        weights1[46387] <= 16'b0000000000101000;
        weights1[46388] <= 16'b0000000000101000;
        weights1[46389] <= 16'b0000000000100101;
        weights1[46390] <= 16'b0000000000110001;
        weights1[46391] <= 16'b0000000000100101;
        weights1[46392] <= 16'b0000000000100011;
        weights1[46393] <= 16'b0000000000010101;
        weights1[46394] <= 16'b0000000000010100;
        weights1[46395] <= 16'b0000000000010110;
        weights1[46396] <= 16'b0000000000001001;
        weights1[46397] <= 16'b0000000000001001;
        weights1[46398] <= 16'b0000000000010110;
        weights1[46399] <= 16'b0000000000010010;
        weights1[46400] <= 16'b0000000000101010;
        weights1[46401] <= 16'b0000000001000010;
        weights1[46402] <= 16'b0000000000100110;
        weights1[46403] <= 16'b0000000000101101;
        weights1[46404] <= 16'b0000000001000001;
        weights1[46405] <= 16'b0000000001000011;
        weights1[46406] <= 16'b0000000000111001;
        weights1[46407] <= 16'b0000000000110001;
        weights1[46408] <= 16'b0000000000100110;
        weights1[46409] <= 16'b0000000000001010;
        weights1[46410] <= 16'b0000000000101111;
        weights1[46411] <= 16'b0000000000100100;
        weights1[46412] <= 16'b0000000000011101;
        weights1[46413] <= 16'b0000000000010010;
        weights1[46414] <= 16'b0000000000101010;
        weights1[46415] <= 16'b0000000000100111;
        weights1[46416] <= 16'b0000000000100001;
        weights1[46417] <= 16'b0000000000011100;
        weights1[46418] <= 16'b0000000000110110;
        weights1[46419] <= 16'b0000000000010001;
        weights1[46420] <= 16'b0000000000001110;
        weights1[46421] <= 16'b0000000000001001;
        weights1[46422] <= 16'b0000000000011001;
        weights1[46423] <= 16'b0000000000001110;
        weights1[46424] <= 16'b0000000000010010;
        weights1[46425] <= 16'b0000000000011010;
        weights1[46426] <= 16'b0000000000011000;
        weights1[46427] <= 16'b0000000000101011;
        weights1[46428] <= 16'b0000000000101001;
        weights1[46429] <= 16'b0000000000110010;
        weights1[46430] <= 16'b0000000000101110;
        weights1[46431] <= 16'b0000000001000111;
        weights1[46432] <= 16'b0000000000101100;
        weights1[46433] <= 16'b0000000000111011;
        weights1[46434] <= 16'b0000000000111110;
        weights1[46435] <= 16'b0000000001000001;
        weights1[46436] <= 16'b0000000000100011;
        weights1[46437] <= 16'b0000000000100010;
        weights1[46438] <= 16'b0000000000111011;
        weights1[46439] <= 16'b0000000000011100;
        weights1[46440] <= 16'b0000000001000000;
        weights1[46441] <= 16'b0000000000011010;
        weights1[46442] <= 16'b0000000000011100;
        weights1[46443] <= 16'b0000000000011110;
        weights1[46444] <= 16'b0000000000010001;
        weights1[46445] <= 16'b0000000000110111;
        weights1[46446] <= 16'b0000000000011011;
        weights1[46447] <= 16'b0000000000101100;
        weights1[46448] <= 16'b0000000000010101;
        weights1[46449] <= 16'b0000000000000011;
        weights1[46450] <= 16'b0000000000011010;
        weights1[46451] <= 16'b0000000000010111;
        weights1[46452] <= 16'b0000000000011011;
        weights1[46453] <= 16'b0000000000101101;
        weights1[46454] <= 16'b0000000000011101;
        weights1[46455] <= 16'b0000000000100010;
        weights1[46456] <= 16'b0000000000100011;
        weights1[46457] <= 16'b0000000000011111;
        weights1[46458] <= 16'b0000000000100000;
        weights1[46459] <= 16'b0000000000100011;
        weights1[46460] <= 16'b0000000000011010;
        weights1[46461] <= 16'b0000000001010010;
        weights1[46462] <= 16'b0000000001010101;
        weights1[46463] <= 16'b0000000001000101;
        weights1[46464] <= 16'b0000000001000010;
        weights1[46465] <= 16'b0000000000111011;
        weights1[46466] <= 16'b0000000001001101;
        weights1[46467] <= 16'b0000000000110000;
        weights1[46468] <= 16'b0000000000100101;
        weights1[46469] <= 16'b0000000000110110;
        weights1[46470] <= 16'b0000000000100000;
        weights1[46471] <= 16'b0000000000010010;
        weights1[46472] <= 16'b0000000000001110;
        weights1[46473] <= 16'b0000000000001110;
        weights1[46474] <= 16'b0000000000101100;
        weights1[46475] <= 16'b0000000001000011;
        weights1[46476] <= 16'b0000000000110011;
        weights1[46477] <= 16'b0000000000010110;
        weights1[46478] <= 16'b0000000000010000;
        weights1[46479] <= 16'b0000000000010101;
        weights1[46480] <= 16'b0000000000100110;
        weights1[46481] <= 16'b0000000000101111;
        weights1[46482] <= 16'b0000000000011111;
        weights1[46483] <= 16'b0000000000011011;
        weights1[46484] <= 16'b0000000000010001;
        weights1[46485] <= 16'b0000000000101110;
        weights1[46486] <= 16'b0000000000100111;
        weights1[46487] <= 16'b0000000000011011;
        weights1[46488] <= 16'b0000000000101110;
        weights1[46489] <= 16'b0000000000110011;
        weights1[46490] <= 16'b0000000000101001;
        weights1[46491] <= 16'b0000000000011101;
        weights1[46492] <= 16'b0000000000011000;
        weights1[46493] <= 16'b0000000000101101;
        weights1[46494] <= 16'b0000000000101111;
        weights1[46495] <= 16'b0000000000100001;
        weights1[46496] <= 16'b0000000000100111;
        weights1[46497] <= 16'b0000000000010110;
        weights1[46498] <= 16'b0000000000010110;
        weights1[46499] <= 16'b0000000000100001;
        weights1[46500] <= 16'b0000000000001001;
        weights1[46501] <= 16'b0000000000001101;
        weights1[46502] <= 16'b0000000000011001;
        weights1[46503] <= 16'b0000000000101110;
        weights1[46504] <= 16'b0000000000110100;
        weights1[46505] <= 16'b0000000000101001;
        weights1[46506] <= 16'b0000000000010000;
        weights1[46507] <= 16'b0000000000011010;
        weights1[46508] <= 16'b0000000000100110;
        weights1[46509] <= 16'b0000000000101011;
        weights1[46510] <= 16'b0000000000100000;
        weights1[46511] <= 16'b0000000000010101;
        weights1[46512] <= 16'b0000000000001011;
        weights1[46513] <= 16'b0000000000010011;
        weights1[46514] <= 16'b0000000000010001;
        weights1[46515] <= 16'b0000000000001100;
        weights1[46516] <= 16'b0000000000010101;
        weights1[46517] <= 16'b0000000000111101;
        weights1[46518] <= 16'b0000000000000111;
        weights1[46519] <= 16'b1111111111010100;
        weights1[46520] <= 16'b1111111111010111;
        weights1[46521] <= 16'b0000000000000010;
        weights1[46522] <= 16'b1111111111111010;
        weights1[46523] <= 16'b1111111111100000;
        weights1[46524] <= 16'b1111111111101010;
        weights1[46525] <= 16'b1111111111110110;
        weights1[46526] <= 16'b1111111111011101;
        weights1[46527] <= 16'b1111111111111010;
        weights1[46528] <= 16'b1111111111110010;
        weights1[46529] <= 16'b0000000000000101;
        weights1[46530] <= 16'b0000000000010001;
        weights1[46531] <= 16'b0000000000101101;
        weights1[46532] <= 16'b0000000000101001;
        weights1[46533] <= 16'b0000000000100011;
        weights1[46534] <= 16'b0000000000100111;
        weights1[46535] <= 16'b0000000000010000;
        weights1[46536] <= 16'b0000000000100111;
        weights1[46537] <= 16'b0000000000101011;
        weights1[46538] <= 16'b0000000000010010;
        weights1[46539] <= 16'b0000000000010101;
        weights1[46540] <= 16'b0000000000001001;
        weights1[46541] <= 16'b0000000000010010;
        weights1[46542] <= 16'b1111111111110110;
        weights1[46543] <= 16'b0000000000010101;
        weights1[46544] <= 16'b0000000000010010;
        weights1[46545] <= 16'b0000000000001101;
        weights1[46546] <= 16'b1111111110111100;
        weights1[46547] <= 16'b1111111101111101;
        weights1[46548] <= 16'b1111111110101011;
        weights1[46549] <= 16'b1111111110111011;
        weights1[46550] <= 16'b1111111110111011;
        weights1[46551] <= 16'b1111111110111011;
        weights1[46552] <= 16'b1111111111010111;
        weights1[46553] <= 16'b1111111111010001;
        weights1[46554] <= 16'b1111111111111000;
        weights1[46555] <= 16'b1111111111111110;
        weights1[46556] <= 16'b1111111111110010;
        weights1[46557] <= 16'b0000000000000000;
        weights1[46558] <= 16'b0000000000011010;
        weights1[46559] <= 16'b0000000000101010;
        weights1[46560] <= 16'b0000000000011110;
        weights1[46561] <= 16'b0000000000101110;
        weights1[46562] <= 16'b0000000000101001;
        weights1[46563] <= 16'b0000000000001110;
        weights1[46564] <= 16'b0000000000100011;
        weights1[46565] <= 16'b0000000000101001;
        weights1[46566] <= 16'b0000000000011111;
        weights1[46567] <= 16'b0000000000001111;
        weights1[46568] <= 16'b0000000000000110;
        weights1[46569] <= 16'b0000000000000010;
        weights1[46570] <= 16'b0000000000000101;
        weights1[46571] <= 16'b0000000000010000;
        weights1[46572] <= 16'b0000000000001101;
        weights1[46573] <= 16'b1111111111100100;
        weights1[46574] <= 16'b1111111101111101;
        weights1[46575] <= 16'b1111111101111110;
        weights1[46576] <= 16'b1111111110111001;
        weights1[46577] <= 16'b1111111111010111;
        weights1[46578] <= 16'b1111111111100001;
        weights1[46579] <= 16'b1111111111010010;
        weights1[46580] <= 16'b1111111111001111;
        weights1[46581] <= 16'b1111111111001110;
        weights1[46582] <= 16'b1111111111000100;
        weights1[46583] <= 16'b1111111111011010;
        weights1[46584] <= 16'b1111111111101010;
        weights1[46585] <= 16'b1111111111101011;
        weights1[46586] <= 16'b1111111111111101;
        weights1[46587] <= 16'b0000000000101000;
        weights1[46588] <= 16'b0000000000100000;
        weights1[46589] <= 16'b0000000000100100;
        weights1[46590] <= 16'b0000000000110101;
        weights1[46591] <= 16'b0000000000010011;
        weights1[46592] <= 16'b0000000000011110;
        weights1[46593] <= 16'b0000000000100011;
        weights1[46594] <= 16'b0000000000011011;
        weights1[46595] <= 16'b0000000000000111;
        weights1[46596] <= 16'b1111111111111110;
        weights1[46597] <= 16'b1111111111111011;
        weights1[46598] <= 16'b0000000000010001;
        weights1[46599] <= 16'b1111111111101001;
        weights1[46600] <= 16'b1111111111111000;
        weights1[46601] <= 16'b1111111110110101;
        weights1[46602] <= 16'b1111111110011100;
        weights1[46603] <= 16'b1111111110111110;
        weights1[46604] <= 16'b1111111111101011;
        weights1[46605] <= 16'b1111111111101001;
        weights1[46606] <= 16'b1111111111001110;
        weights1[46607] <= 16'b1111111111010010;
        weights1[46608] <= 16'b1111111111100100;
        weights1[46609] <= 16'b1111111111001101;
        weights1[46610] <= 16'b1111111111011010;
        weights1[46611] <= 16'b1111111111010100;
        weights1[46612] <= 16'b1111111111101001;
        weights1[46613] <= 16'b1111111111101011;
        weights1[46614] <= 16'b1111111111100111;
        weights1[46615] <= 16'b0000000000010110;
        weights1[46616] <= 16'b0000000000010010;
        weights1[46617] <= 16'b0000000000010001;
        weights1[46618] <= 16'b0000000000010001;
        weights1[46619] <= 16'b0000000000001100;
        weights1[46620] <= 16'b0000000000010010;
        weights1[46621] <= 16'b0000000000011110;
        weights1[46622] <= 16'b0000000000011100;
        weights1[46623] <= 16'b0000000000001010;
        weights1[46624] <= 16'b1111111111111101;
        weights1[46625] <= 16'b1111111111111001;
        weights1[46626] <= 16'b1111111111111001;
        weights1[46627] <= 16'b1111111111101101;
        weights1[46628] <= 16'b1111111111011001;
        weights1[46629] <= 16'b1111111110111011;
        weights1[46630] <= 16'b1111111110011101;
        weights1[46631] <= 16'b1111111111010101;
        weights1[46632] <= 16'b1111111111110101;
        weights1[46633] <= 16'b1111111111011001;
        weights1[46634] <= 16'b1111111111001010;
        weights1[46635] <= 16'b1111111111101101;
        weights1[46636] <= 16'b1111111111011111;
        weights1[46637] <= 16'b1111111111001101;
        weights1[46638] <= 16'b1111111111101010;
        weights1[46639] <= 16'b1111111111001101;
        weights1[46640] <= 16'b1111111111011011;
        weights1[46641] <= 16'b1111111111010000;
        weights1[46642] <= 16'b1111111111110001;
        weights1[46643] <= 16'b0000000000000010;
        weights1[46644] <= 16'b0000000000000011;
        weights1[46645] <= 16'b0000000000000111;
        weights1[46646] <= 16'b0000000000000110;
        weights1[46647] <= 16'b0000000000000010;
        weights1[46648] <= 16'b0000000000001101;
        weights1[46649] <= 16'b0000000000001001;
        weights1[46650] <= 16'b0000000000010100;
        weights1[46651] <= 16'b0000000000001000;
        weights1[46652] <= 16'b1111111111111110;
        weights1[46653] <= 16'b0000000000001000;
        weights1[46654] <= 16'b1111111111101000;
        weights1[46655] <= 16'b1111111111111001;
        weights1[46656] <= 16'b1111111111100011;
        weights1[46657] <= 16'b1111111111011101;
        weights1[46658] <= 16'b1111111110111111;
        weights1[46659] <= 16'b1111111111101101;
        weights1[46660] <= 16'b1111111111111011;
        weights1[46661] <= 16'b1111111111101100;
        weights1[46662] <= 16'b1111111111111001;
        weights1[46663] <= 16'b0000000000010000;
        weights1[46664] <= 16'b1111111111011001;
        weights1[46665] <= 16'b1111111111111000;
        weights1[46666] <= 16'b1111111111110110;
        weights1[46667] <= 16'b1111111111011111;
        weights1[46668] <= 16'b1111111111100100;
        weights1[46669] <= 16'b1111111111110011;
        weights1[46670] <= 16'b0000000000000111;
        weights1[46671] <= 16'b1111111111110110;
        weights1[46672] <= 16'b1111111111111001;
        weights1[46673] <= 16'b1111111111111100;
        weights1[46674] <= 16'b1111111111111111;
        weights1[46675] <= 16'b0000000000000100;
        weights1[46676] <= 16'b1111111111111000;
        weights1[46677] <= 16'b0000000000000010;
        weights1[46678] <= 16'b0000000000000010;
        weights1[46679] <= 16'b0000000000001110;
        weights1[46680] <= 16'b1111111111111101;
        weights1[46681] <= 16'b1111111111111011;
        weights1[46682] <= 16'b0000000000000011;
        weights1[46683] <= 16'b1111111111101101;
        weights1[46684] <= 16'b1111111111110001;
        weights1[46685] <= 16'b1111111111010000;
        weights1[46686] <= 16'b1111111111100000;
        weights1[46687] <= 16'b1111111111011111;
        weights1[46688] <= 16'b1111111111101101;
        weights1[46689] <= 16'b1111111111100101;
        weights1[46690] <= 16'b1111111111101111;
        weights1[46691] <= 16'b1111111111101001;
        weights1[46692] <= 16'b1111111111110111;
        weights1[46693] <= 16'b1111111111011110;
        weights1[46694] <= 16'b1111111111100101;
        weights1[46695] <= 16'b1111111111111001;
        weights1[46696] <= 16'b1111111111110000;
        weights1[46697] <= 16'b1111111111111010;
        weights1[46698] <= 16'b1111111111101011;
        weights1[46699] <= 16'b1111111111110111;
        weights1[46700] <= 16'b1111111111100010;
        weights1[46701] <= 16'b1111111111111100;
        weights1[46702] <= 16'b1111111111111100;
        weights1[46703] <= 16'b1111111111110110;
        weights1[46704] <= 16'b1111111111101101;
        weights1[46705] <= 16'b1111111111111011;
        weights1[46706] <= 16'b1111111111101111;
        weights1[46707] <= 16'b1111111111111110;
        weights1[46708] <= 16'b0000000000000001;
        weights1[46709] <= 16'b0000000000000000;
        weights1[46710] <= 16'b1111111111101101;
        weights1[46711] <= 16'b1111111111110110;
        weights1[46712] <= 16'b1111111111011111;
        weights1[46713] <= 16'b1111111111100000;
        weights1[46714] <= 16'b1111111111010100;
        weights1[46715] <= 16'b1111111111110001;
        weights1[46716] <= 16'b1111111111110011;
        weights1[46717] <= 16'b0000000000001000;
        weights1[46718] <= 16'b1111111111110100;
        weights1[46719] <= 16'b0000000000000101;
        weights1[46720] <= 16'b1111111111111110;
        weights1[46721] <= 16'b1111111111101010;
        weights1[46722] <= 16'b0000000000001000;
        weights1[46723] <= 16'b1111111111101011;
        weights1[46724] <= 16'b1111111111001110;
        weights1[46725] <= 16'b1111111111110111;
        weights1[46726] <= 16'b1111111111101010;
        weights1[46727] <= 16'b1111111111111001;
        weights1[46728] <= 16'b1111111111101010;
        weights1[46729] <= 16'b1111111111101001;
        weights1[46730] <= 16'b1111111111100110;
        weights1[46731] <= 16'b1111111111100111;
        weights1[46732] <= 16'b1111111111110000;
        weights1[46733] <= 16'b1111111111101101;
        weights1[46734] <= 16'b1111111111110000;
        weights1[46735] <= 16'b1111111111110000;
        weights1[46736] <= 16'b1111111111101110;
        weights1[46737] <= 16'b1111111111111000;
        weights1[46738] <= 16'b1111111111101010;
        weights1[46739] <= 16'b1111111111111100;
        weights1[46740] <= 16'b1111111111110000;
        weights1[46741] <= 16'b1111111111110100;
        weights1[46742] <= 16'b1111111111100111;
        weights1[46743] <= 16'b0000000000000111;
        weights1[46744] <= 16'b0000000000000100;
        weights1[46745] <= 16'b1111111111110111;
        weights1[46746] <= 16'b1111111111111111;
        weights1[46747] <= 16'b0000000000000001;
        weights1[46748] <= 16'b1111111111110011;
        weights1[46749] <= 16'b1111111111011000;
        weights1[46750] <= 16'b1111111111100101;
        weights1[46751] <= 16'b1111111111011111;
        weights1[46752] <= 16'b1111111111110000;
        weights1[46753] <= 16'b1111111111111000;
        weights1[46754] <= 16'b1111111111101111;
        weights1[46755] <= 16'b1111111111110001;
        weights1[46756] <= 16'b1111111111010110;
        weights1[46757] <= 16'b1111111111100011;
        weights1[46758] <= 16'b1111111111011111;
        weights1[46759] <= 16'b1111111111100101;
        weights1[46760] <= 16'b1111111111111011;
        weights1[46761] <= 16'b1111111111111010;
        weights1[46762] <= 16'b1111111111110111;
        weights1[46763] <= 16'b1111111111111010;
        weights1[46764] <= 16'b1111111111011111;
        weights1[46765] <= 16'b1111111111111101;
        weights1[46766] <= 16'b1111111111110100;
        weights1[46767] <= 16'b1111111111110101;
        weights1[46768] <= 16'b1111111111100000;
        weights1[46769] <= 16'b1111111111110111;
        weights1[46770] <= 16'b1111111111100000;
        weights1[46771] <= 16'b1111111111100001;
        weights1[46772] <= 16'b0000000000000111;
        weights1[46773] <= 16'b0000000000000011;
        weights1[46774] <= 16'b1111111111110001;
        weights1[46775] <= 16'b0000000000000110;
        weights1[46776] <= 16'b1111111111101001;
        weights1[46777] <= 16'b1111111111100100;
        weights1[46778] <= 16'b1111111111011010;
        weights1[46779] <= 16'b1111111111101110;
        weights1[46780] <= 16'b1111111111110110;
        weights1[46781] <= 16'b1111111111100100;
        weights1[46782] <= 16'b1111111111111001;
        weights1[46783] <= 16'b1111111111101001;
        weights1[46784] <= 16'b1111111111110000;
        weights1[46785] <= 16'b1111111111100100;
        weights1[46786] <= 16'b1111111111100001;
        weights1[46787] <= 16'b1111111111101000;
        weights1[46788] <= 16'b1111111111111010;
        weights1[46789] <= 16'b1111111111111111;
        weights1[46790] <= 16'b0000000000000011;
        weights1[46791] <= 16'b1111111111110010;
        weights1[46792] <= 16'b1111111111110010;
        weights1[46793] <= 16'b1111111111100111;
        weights1[46794] <= 16'b1111111111100010;
        weights1[46795] <= 16'b1111111111111000;
        weights1[46796] <= 16'b1111111111101100;
        weights1[46797] <= 16'b1111111111110110;
        weights1[46798] <= 16'b0000000000000001;
        weights1[46799] <= 16'b1111111111100011;
        weights1[46800] <= 16'b1111111111110110;
        weights1[46801] <= 16'b1111111111101111;
        weights1[46802] <= 16'b1111111111101111;
        weights1[46803] <= 16'b1111111111111010;
        weights1[46804] <= 16'b1111111111100101;
        weights1[46805] <= 16'b1111111111101001;
        weights1[46806] <= 16'b1111111111101100;
        weights1[46807] <= 16'b1111111111100101;
        weights1[46808] <= 16'b1111111111101111;
        weights1[46809] <= 16'b1111111111111000;
        weights1[46810] <= 16'b1111111111110110;
        weights1[46811] <= 16'b1111111111101101;
        weights1[46812] <= 16'b1111111111100000;
        weights1[46813] <= 16'b1111111111101010;
        weights1[46814] <= 16'b1111111111101110;
        weights1[46815] <= 16'b1111111111110010;
        weights1[46816] <= 16'b1111111111111000;
        weights1[46817] <= 16'b1111111111111000;
        weights1[46818] <= 16'b1111111111110101;
        weights1[46819] <= 16'b0000000000001000;
        weights1[46820] <= 16'b1111111111100000;
        weights1[46821] <= 16'b0000000000000011;
        weights1[46822] <= 16'b0000000000001011;
        weights1[46823] <= 16'b1111111111110100;
        weights1[46824] <= 16'b1111111111111101;
        weights1[46825] <= 16'b1111111111111010;
        weights1[46826] <= 16'b1111111111011001;
        weights1[46827] <= 16'b1111111111111111;
        weights1[46828] <= 16'b1111111111110010;
        weights1[46829] <= 16'b0000000000000111;
        weights1[46830] <= 16'b1111111111110100;
        weights1[46831] <= 16'b1111111111100101;
        weights1[46832] <= 16'b1111111111101111;
        weights1[46833] <= 16'b1111111111111010;
        weights1[46834] <= 16'b1111111111100101;
        weights1[46835] <= 16'b1111111111100111;
        weights1[46836] <= 16'b1111111111111011;
        weights1[46837] <= 16'b1111111111111000;
        weights1[46838] <= 16'b1111111111101111;
        weights1[46839] <= 16'b1111111111011001;
        weights1[46840] <= 16'b1111111111001011;
        weights1[46841] <= 16'b1111111111100010;
        weights1[46842] <= 16'b1111111111101111;
        weights1[46843] <= 16'b1111111111111001;
        weights1[46844] <= 16'b1111111111111011;
        weights1[46845] <= 16'b0000000000000000;
        weights1[46846] <= 16'b1111111111111011;
        weights1[46847] <= 16'b1111111111111011;
        weights1[46848] <= 16'b1111111111101111;
        weights1[46849] <= 16'b1111111111101000;
        weights1[46850] <= 16'b1111111111111001;
        weights1[46851] <= 16'b1111111111110100;
        weights1[46852] <= 16'b1111111111011111;
        weights1[46853] <= 16'b1111111111111001;
        weights1[46854] <= 16'b0000000000000001;
        weights1[46855] <= 16'b0000000000000111;
        weights1[46856] <= 16'b0000000000000010;
        weights1[46857] <= 16'b0000000000001110;
        weights1[46858] <= 16'b1111111111100100;
        weights1[46859] <= 16'b1111111111001111;
        weights1[46860] <= 16'b1111111111011111;
        weights1[46861] <= 16'b1111111111100110;
        weights1[46862] <= 16'b1111111111010100;
        weights1[46863] <= 16'b0000000000000010;
        weights1[46864] <= 16'b1111111111111100;
        weights1[46865] <= 16'b1111111111100000;
        weights1[46866] <= 16'b1111111111011011;
        weights1[46867] <= 16'b1111111111010000;
        weights1[46868] <= 16'b1111111111100001;
        weights1[46869] <= 16'b1111111111101100;
        weights1[46870] <= 16'b1111111111110101;
        weights1[46871] <= 16'b1111111111111000;
        weights1[46872] <= 16'b1111111111111110;
        weights1[46873] <= 16'b1111111111111011;
        weights1[46874] <= 16'b1111111111111110;
        weights1[46875] <= 16'b1111111111101110;
        weights1[46876] <= 16'b1111111111110001;
        weights1[46877] <= 16'b1111111111110101;
        weights1[46878] <= 16'b1111111111100010;
        weights1[46879] <= 16'b1111111111101010;
        weights1[46880] <= 16'b1111111111111011;
        weights1[46881] <= 16'b1111111111110001;
        weights1[46882] <= 16'b1111111111110011;
        weights1[46883] <= 16'b1111111111111010;
        weights1[46884] <= 16'b0000000000000010;
        weights1[46885] <= 16'b0000000000001001;
        weights1[46886] <= 16'b1111111111101011;
        weights1[46887] <= 16'b1111111111101101;
        weights1[46888] <= 16'b1111111111111010;
        weights1[46889] <= 16'b1111111111100111;
        weights1[46890] <= 16'b1111111111110101;
        weights1[46891] <= 16'b1111111111110001;
        weights1[46892] <= 16'b1111111111100100;
        weights1[46893] <= 16'b1111111111010100;
        weights1[46894] <= 16'b1111111111010101;
        weights1[46895] <= 16'b1111111111011110;
        weights1[46896] <= 16'b1111111111100010;
        weights1[46897] <= 16'b1111111111101110;
        weights1[46898] <= 16'b1111111111111001;
        weights1[46899] <= 16'b1111111111111011;
        weights1[46900] <= 16'b1111111111111011;
        weights1[46901] <= 16'b1111111111111011;
        weights1[46902] <= 16'b1111111111110101;
        weights1[46903] <= 16'b1111111111111001;
        weights1[46904] <= 16'b1111111111110000;
        weights1[46905] <= 16'b1111111111100110;
        weights1[46906] <= 16'b0000000000001001;
        weights1[46907] <= 16'b1111111111101110;
        weights1[46908] <= 16'b1111111111110010;
        weights1[46909] <= 16'b1111111111110100;
        weights1[46910] <= 16'b0000000000001001;
        weights1[46911] <= 16'b1111111111001101;
        weights1[46912] <= 16'b1111111111101111;
        weights1[46913] <= 16'b1111111111101110;
        weights1[46914] <= 16'b1111111111101101;
        weights1[46915] <= 16'b1111111111010001;
        weights1[46916] <= 16'b1111111111101001;
        weights1[46917] <= 16'b1111111111011000;
        weights1[46918] <= 16'b1111111111010101;
        weights1[46919] <= 16'b1111111111010100;
        weights1[46920] <= 16'b1111111111001111;
        weights1[46921] <= 16'b1111111111010111;
        weights1[46922] <= 16'b1111111111011111;
        weights1[46923] <= 16'b1111111111011011;
        weights1[46924] <= 16'b1111111111100100;
        weights1[46925] <= 16'b1111111111110101;
        weights1[46926] <= 16'b1111111111111101;
        weights1[46927] <= 16'b1111111111111110;
        weights1[46928] <= 16'b1111111111111101;
        weights1[46929] <= 16'b0000000000000010;
        weights1[46930] <= 16'b1111111111111100;
        weights1[46931] <= 16'b1111111111110100;
        weights1[46932] <= 16'b1111111111101001;
        weights1[46933] <= 16'b1111111111110100;
        weights1[46934] <= 16'b1111111111110001;
        weights1[46935] <= 16'b1111111111110100;
        weights1[46936] <= 16'b0000000000000010;
        weights1[46937] <= 16'b1111111111110111;
        weights1[46938] <= 16'b1111111111111101;
        weights1[46939] <= 16'b1111111111111010;
        weights1[46940] <= 16'b1111111111101011;
        weights1[46941] <= 16'b1111111111111100;
        weights1[46942] <= 16'b1111111111010110;
        weights1[46943] <= 16'b1111111111100110;
        weights1[46944] <= 16'b1111111111001001;
        weights1[46945] <= 16'b1111111111001011;
        weights1[46946] <= 16'b1111111110111011;
        weights1[46947] <= 16'b1111111111000101;
        weights1[46948] <= 16'b1111111111010100;
        weights1[46949] <= 16'b1111111111010011;
        weights1[46950] <= 16'b1111111111011111;
        weights1[46951] <= 16'b1111111111101110;
        weights1[46952] <= 16'b1111111111110010;
        weights1[46953] <= 16'b1111111111111010;
        weights1[46954] <= 16'b1111111111111111;
        weights1[46955] <= 16'b1111111111111111;
        weights1[46956] <= 16'b1111111111111110;
        weights1[46957] <= 16'b1111111111111111;
        weights1[46958] <= 16'b1111111111111111;
        weights1[46959] <= 16'b1111111111111001;
        weights1[46960] <= 16'b1111111111110110;
        weights1[46961] <= 16'b1111111111110011;
        weights1[46962] <= 16'b0000000000000011;
        weights1[46963] <= 16'b1111111111111111;
        weights1[46964] <= 16'b0000000000000100;
        weights1[46965] <= 16'b0000000000010100;
        weights1[46966] <= 16'b0000000000001010;
        weights1[46967] <= 16'b1111111111111101;
        weights1[46968] <= 16'b1111111111101110;
        weights1[46969] <= 16'b1111111111111001;
        weights1[46970] <= 16'b1111111111101001;
        weights1[46971] <= 16'b1111111111101101;
        weights1[46972] <= 16'b1111111111010101;
        weights1[46973] <= 16'b1111111110111100;
        weights1[46974] <= 16'b1111111111010110;
        weights1[46975] <= 16'b1111111111010100;
        weights1[46976] <= 16'b1111111111100110;
        weights1[46977] <= 16'b1111111111110000;
        weights1[46978] <= 16'b1111111111101110;
        weights1[46979] <= 16'b1111111111110100;
        weights1[46980] <= 16'b1111111111110111;
        weights1[46981] <= 16'b1111111111111010;
        weights1[46982] <= 16'b1111111111111100;
        weights1[46983] <= 16'b0000000000000000;
        weights1[46984] <= 16'b0000000000000000;
        weights1[46985] <= 16'b1111111111111110;
        weights1[46986] <= 16'b0000000000000001;
        weights1[46987] <= 16'b1111111111111110;
        weights1[46988] <= 16'b1111111111111101;
        weights1[46989] <= 16'b1111111111110000;
        weights1[46990] <= 16'b1111111111111001;
        weights1[46991] <= 16'b1111111111111111;
        weights1[46992] <= 16'b1111111111111001;
        weights1[46993] <= 16'b1111111111111010;
        weights1[46994] <= 16'b1111111111111111;
        weights1[46995] <= 16'b0000000000000100;
        weights1[46996] <= 16'b1111111111111111;
        weights1[46997] <= 16'b0000000000000100;
        weights1[46998] <= 16'b1111111111111001;
        weights1[46999] <= 16'b1111111111111011;
        weights1[47000] <= 16'b1111111111110011;
        weights1[47001] <= 16'b1111111111101011;
        weights1[47002] <= 16'b1111111111100101;
        weights1[47003] <= 16'b1111111111110000;
        weights1[47004] <= 16'b1111111111110100;
        weights1[47005] <= 16'b1111111111110101;
        weights1[47006] <= 16'b1111111111110011;
        weights1[47007] <= 16'b1111111111110111;
        weights1[47008] <= 16'b1111111111111001;
        weights1[47009] <= 16'b1111111111111101;
        weights1[47010] <= 16'b1111111111111111;
        weights1[47011] <= 16'b0000000000000000;
        weights1[47012] <= 16'b0000000000000000;
        weights1[47013] <= 16'b0000000000000000;
        weights1[47014] <= 16'b0000000000000000;
        weights1[47015] <= 16'b1111111111111110;
        weights1[47016] <= 16'b1111111111111100;
        weights1[47017] <= 16'b1111111111111001;
        weights1[47018] <= 16'b1111111111111110;
        weights1[47019] <= 16'b0000000000001000;
        weights1[47020] <= 16'b1111111111111100;
        weights1[47021] <= 16'b0000000000000010;
        weights1[47022] <= 16'b1111111111111101;
        weights1[47023] <= 16'b1111111111111110;
        weights1[47024] <= 16'b1111111111111110;
        weights1[47025] <= 16'b0000000000000100;
        weights1[47026] <= 16'b1111111111111101;
        weights1[47027] <= 16'b1111111111110111;
        weights1[47028] <= 16'b1111111111110011;
        weights1[47029] <= 16'b1111111111110111;
        weights1[47030] <= 16'b1111111111110111;
        weights1[47031] <= 16'b1111111111110111;
        weights1[47032] <= 16'b1111111111110111;
        weights1[47033] <= 16'b1111111111110110;
        weights1[47034] <= 16'b1111111111111000;
        weights1[47035] <= 16'b1111111111111101;
        weights1[47036] <= 16'b1111111111111110;
        weights1[47037] <= 16'b1111111111111110;
        weights1[47038] <= 16'b1111111111111110;
        weights1[47039] <= 16'b1111111111111111;
        weights1[47040] <= 16'b0000000000000000;
        weights1[47041] <= 16'b0000000000000000;
        weights1[47042] <= 16'b1111111111111110;
        weights1[47043] <= 16'b1111111111111011;
        weights1[47044] <= 16'b1111111111111000;
        weights1[47045] <= 16'b1111111111110110;
        weights1[47046] <= 16'b1111111111110010;
        weights1[47047] <= 16'b1111111111110000;
        weights1[47048] <= 16'b1111111111101111;
        weights1[47049] <= 16'b1111111111101100;
        weights1[47050] <= 16'b1111111111101011;
        weights1[47051] <= 16'b1111111111110111;
        weights1[47052] <= 16'b1111111111110111;
        weights1[47053] <= 16'b1111111111110101;
        weights1[47054] <= 16'b1111111111110111;
        weights1[47055] <= 16'b1111111111110111;
        weights1[47056] <= 16'b1111111111110110;
        weights1[47057] <= 16'b1111111111110110;
        weights1[47058] <= 16'b1111111111110101;
        weights1[47059] <= 16'b1111111111110111;
        weights1[47060] <= 16'b1111111111111001;
        weights1[47061] <= 16'b1111111111111101;
        weights1[47062] <= 16'b0000000000000010;
        weights1[47063] <= 16'b1111111111111111;
        weights1[47064] <= 16'b0000000000000001;
        weights1[47065] <= 16'b1111111111111111;
        weights1[47066] <= 16'b1111111111111111;
        weights1[47067] <= 16'b0000000000000000;
        weights1[47068] <= 16'b0000000000000000;
        weights1[47069] <= 16'b0000000000000000;
        weights1[47070] <= 16'b1111111111111100;
        weights1[47071] <= 16'b1111111111111001;
        weights1[47072] <= 16'b1111111111110010;
        weights1[47073] <= 16'b1111111111101101;
        weights1[47074] <= 16'b1111111111101001;
        weights1[47075] <= 16'b1111111111100100;
        weights1[47076] <= 16'b1111111111100111;
        weights1[47077] <= 16'b1111111111100000;
        weights1[47078] <= 16'b1111111111100001;
        weights1[47079] <= 16'b1111111111101110;
        weights1[47080] <= 16'b1111111111100110;
        weights1[47081] <= 16'b1111111111100101;
        weights1[47082] <= 16'b1111111111101001;
        weights1[47083] <= 16'b1111111111101110;
        weights1[47084] <= 16'b1111111111110100;
        weights1[47085] <= 16'b1111111111100110;
        weights1[47086] <= 16'b1111111111110000;
        weights1[47087] <= 16'b1111111111110100;
        weights1[47088] <= 16'b1111111111111001;
        weights1[47089] <= 16'b1111111111110110;
        weights1[47090] <= 16'b1111111111111001;
        weights1[47091] <= 16'b1111111111111010;
        weights1[47092] <= 16'b1111111111111100;
        weights1[47093] <= 16'b1111111111111101;
        weights1[47094] <= 16'b1111111111111101;
        weights1[47095] <= 16'b0000000000000000;
        weights1[47096] <= 16'b1111111111111110;
        weights1[47097] <= 16'b1111111111111110;
        weights1[47098] <= 16'b1111111111111001;
        weights1[47099] <= 16'b1111111111110000;
        weights1[47100] <= 16'b1111111111100101;
        weights1[47101] <= 16'b1111111111100011;
        weights1[47102] <= 16'b1111111111011010;
        weights1[47103] <= 16'b1111111111010111;
        weights1[47104] <= 16'b1111111111011100;
        weights1[47105] <= 16'b1111111111001110;
        weights1[47106] <= 16'b1111111111010011;
        weights1[47107] <= 16'b1111111111001110;
        weights1[47108] <= 16'b1111111111010101;
        weights1[47109] <= 16'b1111111111011001;
        weights1[47110] <= 16'b1111111111011010;
        weights1[47111] <= 16'b1111111111011011;
        weights1[47112] <= 16'b1111111111100001;
        weights1[47113] <= 16'b1111111111011111;
        weights1[47114] <= 16'b1111111111010111;
        weights1[47115] <= 16'b1111111111101001;
        weights1[47116] <= 16'b1111111111101001;
        weights1[47117] <= 16'b1111111111101010;
        weights1[47118] <= 16'b1111111111110011;
        weights1[47119] <= 16'b1111111111110111;
        weights1[47120] <= 16'b1111111111110110;
        weights1[47121] <= 16'b1111111111111000;
        weights1[47122] <= 16'b1111111111111100;
        weights1[47123] <= 16'b1111111111111101;
        weights1[47124] <= 16'b1111111111111111;
        weights1[47125] <= 16'b1111111111111011;
        weights1[47126] <= 16'b1111111111110101;
        weights1[47127] <= 16'b1111111111100101;
        weights1[47128] <= 16'b1111111111010111;
        weights1[47129] <= 16'b1111111111001110;
        weights1[47130] <= 16'b1111111110111100;
        weights1[47131] <= 16'b1111111110111110;
        weights1[47132] <= 16'b1111111110111111;
        weights1[47133] <= 16'b1111111110101101;
        weights1[47134] <= 16'b1111111110011010;
        weights1[47135] <= 16'b1111111110110000;
        weights1[47136] <= 16'b1111111110111101;
        weights1[47137] <= 16'b1111111110110100;
        weights1[47138] <= 16'b1111111110110001;
        weights1[47139] <= 16'b1111111110111100;
        weights1[47140] <= 16'b1111111111000100;
        weights1[47141] <= 16'b1111111111000110;
        weights1[47142] <= 16'b1111111111001100;
        weights1[47143] <= 16'b1111111111010000;
        weights1[47144] <= 16'b1111111111010111;
        weights1[47145] <= 16'b1111111111010100;
        weights1[47146] <= 16'b1111111111101101;
        weights1[47147] <= 16'b1111111111101001;
        weights1[47148] <= 16'b1111111111101101;
        weights1[47149] <= 16'b1111111111111000;
        weights1[47150] <= 16'b1111111111111010;
        weights1[47151] <= 16'b1111111111111010;
        weights1[47152] <= 16'b1111111111111110;
        weights1[47153] <= 16'b1111111111110010;
        weights1[47154] <= 16'b1111111111101010;
        weights1[47155] <= 16'b1111111111100000;
        weights1[47156] <= 16'b1111111111010000;
        weights1[47157] <= 16'b1111111110111010;
        weights1[47158] <= 16'b1111111110101110;
        weights1[47159] <= 16'b1111111110100000;
        weights1[47160] <= 16'b1111111110100011;
        weights1[47161] <= 16'b1111111110010110;
        weights1[47162] <= 16'b1111111110000100;
        weights1[47163] <= 16'b1111111110001010;
        weights1[47164] <= 16'b1111111110010100;
        weights1[47165] <= 16'b1111111110010010;
        weights1[47166] <= 16'b1111111110011011;
        weights1[47167] <= 16'b1111111110100110;
        weights1[47168] <= 16'b1111111110110011;
        weights1[47169] <= 16'b1111111110101110;
        weights1[47170] <= 16'b1111111110101010;
        weights1[47171] <= 16'b1111111110110111;
        weights1[47172] <= 16'b1111111110111110;
        weights1[47173] <= 16'b1111111111001010;
        weights1[47174] <= 16'b1111111111001010;
        weights1[47175] <= 16'b1111111111011000;
        weights1[47176] <= 16'b1111111111011111;
        weights1[47177] <= 16'b1111111111100001;
        weights1[47178] <= 16'b1111111111110000;
        weights1[47179] <= 16'b1111111111110001;
        weights1[47180] <= 16'b1111111111111011;
        weights1[47181] <= 16'b1111111111110111;
        weights1[47182] <= 16'b1111111111100111;
        weights1[47183] <= 16'b1111111111011100;
        weights1[47184] <= 16'b1111111111010100;
        weights1[47185] <= 16'b1111111110111001;
        weights1[47186] <= 16'b1111111110100110;
        weights1[47187] <= 16'b1111111110101101;
        weights1[47188] <= 16'b1111111110101011;
        weights1[47189] <= 16'b1111111110010010;
        weights1[47190] <= 16'b1111111110000000;
        weights1[47191] <= 16'b1111111110000011;
        weights1[47192] <= 16'b1111111110011101;
        weights1[47193] <= 16'b1111111110010010;
        weights1[47194] <= 16'b1111111110010111;
        weights1[47195] <= 16'b1111111111000010;
        weights1[47196] <= 16'b1111111110000110;
        weights1[47197] <= 16'b1111111110010100;
        weights1[47198] <= 16'b1111111110100000;
        weights1[47199] <= 16'b1111111110011001;
        weights1[47200] <= 16'b1111111110001011;
        weights1[47201] <= 16'b1111111110100010;
        weights1[47202] <= 16'b1111111110111000;
        weights1[47203] <= 16'b1111111110101100;
        weights1[47204] <= 16'b1111111110111110;
        weights1[47205] <= 16'b1111111111010110;
        weights1[47206] <= 16'b1111111111011010;
        weights1[47207] <= 16'b1111111111101011;
        weights1[47208] <= 16'b1111111111111011;
        weights1[47209] <= 16'b1111111111111010;
        weights1[47210] <= 16'b1111111111110011;
        weights1[47211] <= 16'b1111111111110110;
        weights1[47212] <= 16'b1111111111111010;
        weights1[47213] <= 16'b1111111111101011;
        weights1[47214] <= 16'b1111111111101111;
        weights1[47215] <= 16'b1111111111001001;
        weights1[47216] <= 16'b1111111111010000;
        weights1[47217] <= 16'b1111111111011101;
        weights1[47218] <= 16'b1111111111011101;
        weights1[47219] <= 16'b1111111111011110;
        weights1[47220] <= 16'b1111111111000101;
        weights1[47221] <= 16'b1111111110111101;
        weights1[47222] <= 16'b1111111111000100;
        weights1[47223] <= 16'b1111111110101101;
        weights1[47224] <= 16'b1111111110110111;
        weights1[47225] <= 16'b1111111111100011;
        weights1[47226] <= 16'b1111111110111100;
        weights1[47227] <= 16'b1111111110110100;
        weights1[47228] <= 16'b1111111110101010;
        weights1[47229] <= 16'b1111111111010110;
        weights1[47230] <= 16'b1111111111000111;
        weights1[47231] <= 16'b1111111110111001;
        weights1[47232] <= 16'b1111111111001011;
        weights1[47233] <= 16'b1111111111011000;
        weights1[47234] <= 16'b1111111111011110;
        weights1[47235] <= 16'b1111111111101011;
        weights1[47236] <= 16'b0000000000000001;
        weights1[47237] <= 16'b1111111111111110;
        weights1[47238] <= 16'b1111111111111101;
        weights1[47239] <= 16'b1111111111110100;
        weights1[47240] <= 16'b0000000000001100;
        weights1[47241] <= 16'b0000000000001110;
        weights1[47242] <= 16'b0000000000011111;
        weights1[47243] <= 16'b0000000000100101;
        weights1[47244] <= 16'b0000000000011001;
        weights1[47245] <= 16'b0000000000011101;
        weights1[47246] <= 16'b0000000000001000;
        weights1[47247] <= 16'b0000000000000001;
        weights1[47248] <= 16'b1111111111111001;
        weights1[47249] <= 16'b1111111111101111;
        weights1[47250] <= 16'b0000000000001111;
        weights1[47251] <= 16'b1111111111100000;
        weights1[47252] <= 16'b1111111111101100;
        weights1[47253] <= 16'b1111111111110110;
        weights1[47254] <= 16'b1111111111100111;
        weights1[47255] <= 16'b1111111111110110;
        weights1[47256] <= 16'b1111111111101011;
        weights1[47257] <= 16'b1111111111101100;
        weights1[47258] <= 16'b1111111111111001;
        weights1[47259] <= 16'b0000000000001010;
        weights1[47260] <= 16'b0000000000000010;
        weights1[47261] <= 16'b1111111111100100;
        weights1[47262] <= 16'b1111111111110111;
        weights1[47263] <= 16'b1111111111111011;
        weights1[47264] <= 16'b1111111111111100;
        weights1[47265] <= 16'b1111111111111110;
        weights1[47266] <= 16'b1111111111111101;
        weights1[47267] <= 16'b0000000000000000;
        weights1[47268] <= 16'b0000000000000101;
        weights1[47269] <= 16'b0000000000100011;
        weights1[47270] <= 16'b0000000000001001;
        weights1[47271] <= 16'b0000000000110110;
        weights1[47272] <= 16'b0000000000110000;
        weights1[47273] <= 16'b0000000000100100;
        weights1[47274] <= 16'b0000000000101100;
        weights1[47275] <= 16'b0000000000100111;
        weights1[47276] <= 16'b0000000000110001;
        weights1[47277] <= 16'b0000000000010111;
        weights1[47278] <= 16'b0000000000010000;
        weights1[47279] <= 16'b0000000000001110;
        weights1[47280] <= 16'b1111111111111110;
        weights1[47281] <= 16'b0000000000010101;
        weights1[47282] <= 16'b0000000000010101;
        weights1[47283] <= 16'b0000000000010101;
        weights1[47284] <= 16'b0000000000100010;
        weights1[47285] <= 16'b0000000000011001;
        weights1[47286] <= 16'b0000000000001110;
        weights1[47287] <= 16'b0000000000100000;
        weights1[47288] <= 16'b0000000000011100;
        weights1[47289] <= 16'b0000000000100000;
        weights1[47290] <= 16'b0000000000001111;
        weights1[47291] <= 16'b0000000000001110;
        weights1[47292] <= 16'b0000000000000011;
        weights1[47293] <= 16'b0000000000000100;
        weights1[47294] <= 16'b0000000000000111;
        weights1[47295] <= 16'b0000000000000101;
        weights1[47296] <= 16'b0000000000000001;
        weights1[47297] <= 16'b0000000000010011;
        weights1[47298] <= 16'b0000000000010111;
        weights1[47299] <= 16'b0000000000010101;
        weights1[47300] <= 16'b0000000000101101;
        weights1[47301] <= 16'b0000000000111100;
        weights1[47302] <= 16'b0000000000110101;
        weights1[47303] <= 16'b0000000000101110;
        weights1[47304] <= 16'b0000000001000010;
        weights1[47305] <= 16'b0000000000011111;
        weights1[47306] <= 16'b0000000000100101;
        weights1[47307] <= 16'b0000000000010001;
        weights1[47308] <= 16'b0000000000100101;
        weights1[47309] <= 16'b0000000000011001;
        weights1[47310] <= 16'b0000000000010001;
        weights1[47311] <= 16'b0000000000010100;
        weights1[47312] <= 16'b0000000000010111;
        weights1[47313] <= 16'b0000000000001110;
        weights1[47314] <= 16'b0000000000011010;
        weights1[47315] <= 16'b1111111111111110;
        weights1[47316] <= 16'b0000000000100100;
        weights1[47317] <= 16'b0000000000011101;
        weights1[47318] <= 16'b0000000000000100;
        weights1[47319] <= 16'b0000000000010100;
        weights1[47320] <= 16'b0000000000001000;
        weights1[47321] <= 16'b0000000000000100;
        weights1[47322] <= 16'b0000000000000100;
        weights1[47323] <= 16'b1111111111111110;
        weights1[47324] <= 16'b0000000000000110;
        weights1[47325] <= 16'b1111111111111110;
        weights1[47326] <= 16'b0000000000010010;
        weights1[47327] <= 16'b0000000000001001;
        weights1[47328] <= 16'b0000000000001111;
        weights1[47329] <= 16'b0000000000011111;
        weights1[47330] <= 16'b0000000000011101;
        weights1[47331] <= 16'b0000000000101010;
        weights1[47332] <= 16'b0000000000101001;
        weights1[47333] <= 16'b0000000001011001;
        weights1[47334] <= 16'b0000000000111100;
        weights1[47335] <= 16'b0000000001000101;
        weights1[47336] <= 16'b0000000000111010;
        weights1[47337] <= 16'b0000000000100010;
        weights1[47338] <= 16'b0000000000110001;
        weights1[47339] <= 16'b0000000000101100;
        weights1[47340] <= 16'b0000000000001001;
        weights1[47341] <= 16'b0000000000010110;
        weights1[47342] <= 16'b0000000000001000;
        weights1[47343] <= 16'b0000000000010101;
        weights1[47344] <= 16'b0000000000001110;
        weights1[47345] <= 16'b0000000000001110;
        weights1[47346] <= 16'b0000000000001110;
        weights1[47347] <= 16'b0000000000001100;
        weights1[47348] <= 16'b0000000000000111;
        weights1[47349] <= 16'b0000000000000011;
        weights1[47350] <= 16'b0000000000001010;
        weights1[47351] <= 16'b1111111111110111;
        weights1[47352] <= 16'b1111111111110110;
        weights1[47353] <= 16'b1111111111100110;
        weights1[47354] <= 16'b0000000000000111;
        weights1[47355] <= 16'b0000000000000101;
        weights1[47356] <= 16'b1111111111101110;
        weights1[47357] <= 16'b0000000000001000;
        weights1[47358] <= 16'b1111111111110100;
        weights1[47359] <= 16'b0000000000100000;
        weights1[47360] <= 16'b0000000000011100;
        weights1[47361] <= 16'b0000000000100110;
        weights1[47362] <= 16'b0000000000111000;
        weights1[47363] <= 16'b0000000000111011;
        weights1[47364] <= 16'b0000000000111010;
        weights1[47365] <= 16'b0000000000111010;
        weights1[47366] <= 16'b0000000000011100;
        weights1[47367] <= 16'b0000000000111000;
        weights1[47368] <= 16'b0000000000100000;
        weights1[47369] <= 16'b0000000000001010;
        weights1[47370] <= 16'b0000000000011010;
        weights1[47371] <= 16'b0000000000000100;
        weights1[47372] <= 16'b1111111111111111;
        weights1[47373] <= 16'b0000000000001010;
        weights1[47374] <= 16'b1111111111111101;
        weights1[47375] <= 16'b0000000000001000;
        weights1[47376] <= 16'b0000000000000011;
        weights1[47377] <= 16'b1111111111110111;
        weights1[47378] <= 16'b0000000000000010;
        weights1[47379] <= 16'b1111111111110111;
        weights1[47380] <= 16'b1111111111110110;
        weights1[47381] <= 16'b1111111111101110;
        weights1[47382] <= 16'b0000000000001101;
        weights1[47383] <= 16'b1111111111110001;
        weights1[47384] <= 16'b1111111111111001;
        weights1[47385] <= 16'b1111111111110000;
        weights1[47386] <= 16'b1111111111101110;
        weights1[47387] <= 16'b1111111111101101;
        weights1[47388] <= 16'b1111111111011100;
        weights1[47389] <= 16'b1111111111110110;
        weights1[47390] <= 16'b0000000000001100;
        weights1[47391] <= 16'b0000000000010010;
        weights1[47392] <= 16'b0000000000011011;
        weights1[47393] <= 16'b1111111111111101;
        weights1[47394] <= 16'b1111111111111101;
        weights1[47395] <= 16'b0000000000010110;
        weights1[47396] <= 16'b0000000000000001;
        weights1[47397] <= 16'b1111111111101101;
        weights1[47398] <= 16'b0000000000000000;
        weights1[47399] <= 16'b1111111111111001;
        weights1[47400] <= 16'b1111111111111001;
        weights1[47401] <= 16'b0000000000010010;
        weights1[47402] <= 16'b1111111111110000;
        weights1[47403] <= 16'b1111111111111101;
        weights1[47404] <= 16'b0000000000000111;
        weights1[47405] <= 16'b1111111111110001;
        weights1[47406] <= 16'b0000000000001110;
        weights1[47407] <= 16'b1111111111110100;
        weights1[47408] <= 16'b1111111111110011;
        weights1[47409] <= 16'b1111111111111010;
        weights1[47410] <= 16'b1111111111111111;
        weights1[47411] <= 16'b1111111111111001;
        weights1[47412] <= 16'b1111111111111101;
        weights1[47413] <= 16'b1111111111111111;
        weights1[47414] <= 16'b1111111111101110;
        weights1[47415] <= 16'b1111111111101110;
        weights1[47416] <= 16'b1111111111101010;
        weights1[47417] <= 16'b1111111111100100;
        weights1[47418] <= 16'b1111111111010100;
        weights1[47419] <= 16'b1111111111100110;
        weights1[47420] <= 16'b1111111111101011;
        weights1[47421] <= 16'b1111111111110100;
        weights1[47422] <= 16'b1111111111111001;
        weights1[47423] <= 16'b1111111111101000;
        weights1[47424] <= 16'b1111111111101010;
        weights1[47425] <= 16'b0000000000001101;
        weights1[47426] <= 16'b0000000000001001;
        weights1[47427] <= 16'b1111111111111101;
        weights1[47428] <= 16'b1111111111101000;
        weights1[47429] <= 16'b0000000000000010;
        weights1[47430] <= 16'b1111111111111101;
        weights1[47431] <= 16'b1111111111111101;
        weights1[47432] <= 16'b0000000000000000;
        weights1[47433] <= 16'b1111111111110111;
        weights1[47434] <= 16'b0000000000000000;
        weights1[47435] <= 16'b0000000000011010;
        weights1[47436] <= 16'b0000000000000000;
        weights1[47437] <= 16'b1111111111111010;
        weights1[47438] <= 16'b1111111111111111;
        weights1[47439] <= 16'b1111111111111111;
        weights1[47440] <= 16'b1111111111111110;
        weights1[47441] <= 16'b1111111111110101;
        weights1[47442] <= 16'b0000000000000100;
        weights1[47443] <= 16'b0000000000000010;
        weights1[47444] <= 16'b1111111111101011;
        weights1[47445] <= 16'b1111111111101101;
        weights1[47446] <= 16'b1111111111100111;
        weights1[47447] <= 16'b1111111111010010;
        weights1[47448] <= 16'b1111111111100101;
        weights1[47449] <= 16'b0000000000001101;
        weights1[47450] <= 16'b1111111111101111;
        weights1[47451] <= 16'b1111111111111010;
        weights1[47452] <= 16'b0000000000000000;
        weights1[47453] <= 16'b1111111111110110;
        weights1[47454] <= 16'b1111111111111111;
        weights1[47455] <= 16'b0000000000001001;
        weights1[47456] <= 16'b0000000000010011;
        weights1[47457] <= 16'b1111111111101111;
        weights1[47458] <= 16'b1111111111111010;
        weights1[47459] <= 16'b1111111111111011;
        weights1[47460] <= 16'b0000000000000010;
        weights1[47461] <= 16'b0000000000000011;
        weights1[47462] <= 16'b1111111111111111;
        weights1[47463] <= 16'b0000000000100000;
        weights1[47464] <= 16'b0000000000100000;
        weights1[47465] <= 16'b1111111111111001;
        weights1[47466] <= 16'b0000000000011110;
        weights1[47467] <= 16'b0000000000010101;
        weights1[47468] <= 16'b1111111111110111;
        weights1[47469] <= 16'b0000000000000100;
        weights1[47470] <= 16'b0000000000000100;
        weights1[47471] <= 16'b1111111111110101;
        weights1[47472] <= 16'b1111111111110001;
        weights1[47473] <= 16'b1111111111101000;
        weights1[47474] <= 16'b1111111111100000;
        weights1[47475] <= 16'b1111111111111000;
        weights1[47476] <= 16'b1111111111011101;
        weights1[47477] <= 16'b1111111111100110;
        weights1[47478] <= 16'b1111111111111011;
        weights1[47479] <= 16'b0000000000000001;
        weights1[47480] <= 16'b0000000000000101;
        weights1[47481] <= 16'b0000000000100011;
        weights1[47482] <= 16'b1111111111101001;
        weights1[47483] <= 16'b0000000000001001;
        weights1[47484] <= 16'b0000000000100110;
        weights1[47485] <= 16'b0000000000000000;
        weights1[47486] <= 16'b1111111111101100;
        weights1[47487] <= 16'b0000000000000110;
        weights1[47488] <= 16'b0000000000000101;
        weights1[47489] <= 16'b0000000000001100;
        weights1[47490] <= 16'b0000000000010100;
        weights1[47491] <= 16'b0000000000010001;
        weights1[47492] <= 16'b0000000000000110;
        weights1[47493] <= 16'b1111111111100011;
        weights1[47494] <= 16'b0000000000000011;
        weights1[47495] <= 16'b1111111111110100;
        weights1[47496] <= 16'b1111111111111010;
        weights1[47497] <= 16'b1111111111111000;
        weights1[47498] <= 16'b1111111111110001;
        weights1[47499] <= 16'b1111111111011000;
        weights1[47500] <= 16'b1111111111110101;
        weights1[47501] <= 16'b1111111111101001;
        weights1[47502] <= 16'b1111111111101111;
        weights1[47503] <= 16'b1111111111111001;
        weights1[47504] <= 16'b1111111111110110;
        weights1[47505] <= 16'b0000000000000111;
        weights1[47506] <= 16'b1111111111110111;
        weights1[47507] <= 16'b1111111111110111;
        weights1[47508] <= 16'b0000000000001011;
        weights1[47509] <= 16'b0000000000000010;
        weights1[47510] <= 16'b0000000000001101;
        weights1[47511] <= 16'b1111111111111011;
        weights1[47512] <= 16'b1111111111111000;
        weights1[47513] <= 16'b1111111111111000;
        weights1[47514] <= 16'b0000000000000010;
        weights1[47515] <= 16'b0000000000010001;
        weights1[47516] <= 16'b1111111111110110;
        weights1[47517] <= 16'b0000000000000011;
        weights1[47518] <= 16'b0000000000010111;
        weights1[47519] <= 16'b0000000000010111;
        weights1[47520] <= 16'b0000000000010010;
        weights1[47521] <= 16'b0000000000010111;
        weights1[47522] <= 16'b0000000000000100;
        weights1[47523] <= 16'b1111111111111100;
        weights1[47524] <= 16'b1111111111111100;
        weights1[47525] <= 16'b1111111111110001;
        weights1[47526] <= 16'b0000000000000011;
        weights1[47527] <= 16'b0000000000000011;
        weights1[47528] <= 16'b1111111111111100;
        weights1[47529] <= 16'b0000000000000001;
        weights1[47530] <= 16'b0000000000000000;
        weights1[47531] <= 16'b1111111111110101;
        weights1[47532] <= 16'b1111111111110101;
        weights1[47533] <= 16'b1111111111111111;
        weights1[47534] <= 16'b0000000000000010;
        weights1[47535] <= 16'b1111111111111010;
        weights1[47536] <= 16'b1111111111111111;
        weights1[47537] <= 16'b0000000000000001;
        weights1[47538] <= 16'b0000000000000101;
        weights1[47539] <= 16'b0000000000010010;
        weights1[47540] <= 16'b0000000000000100;
        weights1[47541] <= 16'b0000000000000000;
        weights1[47542] <= 16'b0000000000000011;
        weights1[47543] <= 16'b0000000000000011;
        weights1[47544] <= 16'b1111111111110110;
        weights1[47545] <= 16'b0000000000000101;
        weights1[47546] <= 16'b0000000000010000;
        weights1[47547] <= 16'b1111111111111100;
        weights1[47548] <= 16'b0000000000000011;
        weights1[47549] <= 16'b0000000000000000;
        weights1[47550] <= 16'b0000000000001010;
        weights1[47551] <= 16'b1111111111110111;
        weights1[47552] <= 16'b1111111111110111;
        weights1[47553] <= 16'b1111111111111001;
        weights1[47554] <= 16'b1111111111111100;
        weights1[47555] <= 16'b0000000000010011;
        weights1[47556] <= 16'b0000000000001110;
        weights1[47557] <= 16'b1111111111110010;
        weights1[47558] <= 16'b0000000000010100;
        weights1[47559] <= 16'b1111111111110000;
        weights1[47560] <= 16'b1111111111101101;
        weights1[47561] <= 16'b1111111111111011;
        weights1[47562] <= 16'b0000000000000000;
        weights1[47563] <= 16'b1111111111110111;
        weights1[47564] <= 16'b1111111111111101;
        weights1[47565] <= 16'b0000000000000100;
        weights1[47566] <= 16'b0000000000001000;
        weights1[47567] <= 16'b0000000000000101;
        weights1[47568] <= 16'b1111111111110101;
        weights1[47569] <= 16'b1111111111110100;
        weights1[47570] <= 16'b1111111111111100;
        weights1[47571] <= 16'b0000000000001010;
        weights1[47572] <= 16'b1111111111101110;
        weights1[47573] <= 16'b1111111111111000;
        weights1[47574] <= 16'b1111111111111100;
        weights1[47575] <= 16'b1111111111101100;
        weights1[47576] <= 16'b1111111111100100;
        weights1[47577] <= 16'b1111111111101110;
        weights1[47578] <= 16'b1111111111110000;
        weights1[47579] <= 16'b0000000000000111;
        weights1[47580] <= 16'b0000000000010011;
        weights1[47581] <= 16'b0000000000001001;
        weights1[47582] <= 16'b1111111111111101;
        weights1[47583] <= 16'b0000000000000000;
        weights1[47584] <= 16'b0000000000010001;
        weights1[47585] <= 16'b1111111111111000;
        weights1[47586] <= 16'b0000000000010001;
        weights1[47587] <= 16'b1111111111111010;
        weights1[47588] <= 16'b1111111111111011;
        weights1[47589] <= 16'b0000000000000100;
        weights1[47590] <= 16'b1111111111110110;
        weights1[47591] <= 16'b1111111111111111;
        weights1[47592] <= 16'b1111111111111111;
        weights1[47593] <= 16'b1111111111110111;
        weights1[47594] <= 16'b1111111111111100;
        weights1[47595] <= 16'b0000000000001001;
        weights1[47596] <= 16'b1111111111111101;
        weights1[47597] <= 16'b0000000000000110;
        weights1[47598] <= 16'b1111111111111000;
        weights1[47599] <= 16'b1111111111111111;
        weights1[47600] <= 16'b1111111111101111;
        weights1[47601] <= 16'b1111111111110001;
        weights1[47602] <= 16'b1111111111110100;
        weights1[47603] <= 16'b1111111111110101;
        weights1[47604] <= 16'b1111111111100100;
        weights1[47605] <= 16'b0000000000000100;
        weights1[47606] <= 16'b0000000000000111;
        weights1[47607] <= 16'b1111111111101001;
        weights1[47608] <= 16'b1111111111111101;
        weights1[47609] <= 16'b0000000000010001;
        weights1[47610] <= 16'b0000000000010001;
        weights1[47611] <= 16'b0000000000010001;
        weights1[47612] <= 16'b0000000000001010;
        weights1[47613] <= 16'b1111111111111000;
        weights1[47614] <= 16'b0000000000000010;
        weights1[47615] <= 16'b0000000000001010;
        weights1[47616] <= 16'b1111111111110001;
        weights1[47617] <= 16'b1111111111111100;
        weights1[47618] <= 16'b1111111111111100;
        weights1[47619] <= 16'b1111111111101110;
        weights1[47620] <= 16'b0000000000000101;
        weights1[47621] <= 16'b1111111111101111;
        weights1[47622] <= 16'b0000000000001001;
        weights1[47623] <= 16'b1111111111110011;
        weights1[47624] <= 16'b1111111111111101;
        weights1[47625] <= 16'b0000000000000010;
        weights1[47626] <= 16'b1111111111110010;
        weights1[47627] <= 16'b1111111111101101;
        weights1[47628] <= 16'b1111111111110011;
        weights1[47629] <= 16'b1111111111101011;
        weights1[47630] <= 16'b1111111111110100;
        weights1[47631] <= 16'b1111111111110111;
        weights1[47632] <= 16'b1111111111110100;
        weights1[47633] <= 16'b1111111111101111;
        weights1[47634] <= 16'b1111111111110011;
        weights1[47635] <= 16'b1111111111011001;
        weights1[47636] <= 16'b1111111111101100;
        weights1[47637] <= 16'b1111111111111011;
        weights1[47638] <= 16'b1111111111011110;
        weights1[47639] <= 16'b1111111111111001;
        weights1[47640] <= 16'b1111111111111011;
        weights1[47641] <= 16'b0000000000000110;
        weights1[47642] <= 16'b1111111111111110;
        weights1[47643] <= 16'b1111111111110111;
        weights1[47644] <= 16'b1111111111110111;
        weights1[47645] <= 16'b0000000000001011;
        weights1[47646] <= 16'b1111111111101101;
        weights1[47647] <= 16'b0000000000000000;
        weights1[47648] <= 16'b1111111111110111;
        weights1[47649] <= 16'b0000000000000111;
        weights1[47650] <= 16'b0000000000001000;
        weights1[47651] <= 16'b1111111111101110;
        weights1[47652] <= 16'b1111111111111000;
        weights1[47653] <= 16'b1111111111110010;
        weights1[47654] <= 16'b1111111111110110;
        weights1[47655] <= 16'b1111111111110101;
        weights1[47656] <= 16'b1111111111101110;
        weights1[47657] <= 16'b1111111111101110;
        weights1[47658] <= 16'b1111111111110110;
        weights1[47659] <= 16'b0000000000001111;
        weights1[47660] <= 16'b1111111111111000;
        weights1[47661] <= 16'b1111111111100011;
        weights1[47662] <= 16'b1111111111111100;
        weights1[47663] <= 16'b1111111111100110;
        weights1[47664] <= 16'b1111111111111111;
        weights1[47665] <= 16'b1111111111111010;
        weights1[47666] <= 16'b1111111111110110;
        weights1[47667] <= 16'b1111111111100010;
        weights1[47668] <= 16'b1111111111110101;
        weights1[47669] <= 16'b1111111111100110;
        weights1[47670] <= 16'b0000000000000010;
        weights1[47671] <= 16'b1111111111111100;
        weights1[47672] <= 16'b1111111111111010;
        weights1[47673] <= 16'b1111111111110100;
        weights1[47674] <= 16'b1111111111111011;
        weights1[47675] <= 16'b1111111111111101;
        weights1[47676] <= 16'b1111111111111110;
        weights1[47677] <= 16'b1111111111111110;
        weights1[47678] <= 16'b0000000000000000;
        weights1[47679] <= 16'b1111111111110010;
        weights1[47680] <= 16'b0000000000000011;
        weights1[47681] <= 16'b1111111111110000;
        weights1[47682] <= 16'b1111111111110011;
        weights1[47683] <= 16'b1111111111110101;
        weights1[47684] <= 16'b1111111111110110;
        weights1[47685] <= 16'b1111111111110101;
        weights1[47686] <= 16'b1111111111110111;
        weights1[47687] <= 16'b1111111111111000;
        weights1[47688] <= 16'b1111111111110111;
        weights1[47689] <= 16'b0000000000000000;
        weights1[47690] <= 16'b1111111111011101;
        weights1[47691] <= 16'b1111111111111001;
        weights1[47692] <= 16'b1111111111111111;
        weights1[47693] <= 16'b1111111111011001;
        weights1[47694] <= 16'b1111111111110001;
        weights1[47695] <= 16'b0000000000000001;
        weights1[47696] <= 16'b1111111111101101;
        weights1[47697] <= 16'b1111111111110010;
        weights1[47698] <= 16'b1111111111111111;
        weights1[47699] <= 16'b1111111111101110;
        weights1[47700] <= 16'b0000000000001000;
        weights1[47701] <= 16'b1111111111111100;
        weights1[47702] <= 16'b1111111111111010;
        weights1[47703] <= 16'b1111111111111100;
        weights1[47704] <= 16'b1111111111110101;
        weights1[47705] <= 16'b0000000000000110;
        weights1[47706] <= 16'b1111111111110110;
        weights1[47707] <= 16'b1111111111111000;
        weights1[47708] <= 16'b1111111111101101;
        weights1[47709] <= 16'b1111111111101100;
        weights1[47710] <= 16'b1111111111111000;
        weights1[47711] <= 16'b1111111111111000;
        weights1[47712] <= 16'b1111111111111010;
        weights1[47713] <= 16'b1111111111111010;
        weights1[47714] <= 16'b1111111111101110;
        weights1[47715] <= 16'b1111111111110101;
        weights1[47716] <= 16'b1111111111101000;
        weights1[47717] <= 16'b1111111111111100;
        weights1[47718] <= 16'b1111111111011000;
        weights1[47719] <= 16'b1111111111101101;
        weights1[47720] <= 16'b1111111111101111;
        weights1[47721] <= 16'b1111111111100110;
        weights1[47722] <= 16'b1111111111110111;
        weights1[47723] <= 16'b1111111111101100;
        weights1[47724] <= 16'b0000000000000011;
        weights1[47725] <= 16'b1111111111111110;
        weights1[47726] <= 16'b1111111111110111;
        weights1[47727] <= 16'b1111111111110001;
        weights1[47728] <= 16'b0000000000000000;
        weights1[47729] <= 16'b1111111111110000;
        weights1[47730] <= 16'b1111111111110011;
        weights1[47731] <= 16'b1111111111110101;
        weights1[47732] <= 16'b1111111111100010;
        weights1[47733] <= 16'b1111111111100111;
        weights1[47734] <= 16'b1111111111111001;
        weights1[47735] <= 16'b1111111111110111;
        weights1[47736] <= 16'b1111111111101011;
        weights1[47737] <= 16'b1111111111100011;
        weights1[47738] <= 16'b1111111111110001;
        weights1[47739] <= 16'b1111111111110111;
        weights1[47740] <= 16'b1111111111111101;
        weights1[47741] <= 16'b1111111111110101;
        weights1[47742] <= 16'b1111111111110100;
        weights1[47743] <= 16'b1111111111101011;
        weights1[47744] <= 16'b1111111111101011;
        weights1[47745] <= 16'b1111111111100001;
        weights1[47746] <= 16'b1111111111101111;
        weights1[47747] <= 16'b0000000000001000;
        weights1[47748] <= 16'b1111111111100111;
        weights1[47749] <= 16'b1111111111101110;
        weights1[47750] <= 16'b1111111111100101;
        weights1[47751] <= 16'b0000000000000010;
        weights1[47752] <= 16'b0000000000000110;
        weights1[47753] <= 16'b1111111111101110;
        weights1[47754] <= 16'b1111111111110100;
        weights1[47755] <= 16'b1111111111110010;
        weights1[47756] <= 16'b0000000000000110;
        weights1[47757] <= 16'b1111111111011001;
        weights1[47758] <= 16'b1111111111111100;
        weights1[47759] <= 16'b0000000000000011;
        weights1[47760] <= 16'b1111111111101010;
        weights1[47761] <= 16'b1111111111101011;
        weights1[47762] <= 16'b1111111111110110;
        weights1[47763] <= 16'b1111111111111100;
        weights1[47764] <= 16'b1111111111110110;
        weights1[47765] <= 16'b1111111111100111;
        weights1[47766] <= 16'b1111111111110101;
        weights1[47767] <= 16'b1111111111111110;
        weights1[47768] <= 16'b1111111111111110;
        weights1[47769] <= 16'b1111111111110101;
        weights1[47770] <= 16'b1111111111110011;
        weights1[47771] <= 16'b1111111111101101;
        weights1[47772] <= 16'b1111111111101010;
        weights1[47773] <= 16'b1111111111011100;
        weights1[47774] <= 16'b1111111111101111;
        weights1[47775] <= 16'b0000000000000001;
        weights1[47776] <= 16'b0000000000001000;
        weights1[47777] <= 16'b0000000000001010;
        weights1[47778] <= 16'b1111111111101111;
        weights1[47779] <= 16'b1111111111110110;
        weights1[47780] <= 16'b1111111111111110;
        weights1[47781] <= 16'b0000000000001011;
        weights1[47782] <= 16'b1111111111101101;
        weights1[47783] <= 16'b1111111111110100;
        weights1[47784] <= 16'b1111111111111111;
        weights1[47785] <= 16'b1111111111111011;
        weights1[47786] <= 16'b1111111111110101;
        weights1[47787] <= 16'b0000000000000000;
        weights1[47788] <= 16'b1111111111101110;
        weights1[47789] <= 16'b1111111111110101;
        weights1[47790] <= 16'b1111111111110100;
        weights1[47791] <= 16'b1111111111101010;
        weights1[47792] <= 16'b0000000000000000;
        weights1[47793] <= 16'b0000000000000000;
        weights1[47794] <= 16'b0000000000000101;
        weights1[47795] <= 16'b0000000000000001;
        weights1[47796] <= 16'b1111111111111101;
        weights1[47797] <= 16'b1111111111111000;
        weights1[47798] <= 16'b1111111111110000;
        weights1[47799] <= 16'b1111111111110100;
        weights1[47800] <= 16'b1111111111110110;
        weights1[47801] <= 16'b1111111111111101;
        weights1[47802] <= 16'b1111111111111011;
        weights1[47803] <= 16'b1111111111110101;
        weights1[47804] <= 16'b1111111111110000;
        weights1[47805] <= 16'b1111111111110001;
        weights1[47806] <= 16'b1111111111110101;
        weights1[47807] <= 16'b1111111111101010;
        weights1[47808] <= 16'b1111111111011100;
        weights1[47809] <= 16'b1111111111110001;
        weights1[47810] <= 16'b1111111111111001;
        weights1[47811] <= 16'b1111111111110001;
        weights1[47812] <= 16'b1111111111101011;
        weights1[47813] <= 16'b1111111111100011;
        weights1[47814] <= 16'b0000000000001101;
        weights1[47815] <= 16'b1111111111110010;
        weights1[47816] <= 16'b1111111111101000;
        weights1[47817] <= 16'b1111111111110000;
        weights1[47818] <= 16'b0000000000000001;
        weights1[47819] <= 16'b1111111111110111;
        weights1[47820] <= 16'b1111111111111101;
        weights1[47821] <= 16'b1111111111111101;
        weights1[47822] <= 16'b0000000000001010;
        weights1[47823] <= 16'b0000000000000101;
        weights1[47824] <= 16'b0000000000000000;
        weights1[47825] <= 16'b0000000000000000;
        weights1[47826] <= 16'b0000000000000000;
        weights1[47827] <= 16'b0000000000000001;
        weights1[47828] <= 16'b0000000000000010;
        weights1[47829] <= 16'b0000000000000010;
        weights1[47830] <= 16'b0000000000000000;
        weights1[47831] <= 16'b0000000000000001;
        weights1[47832] <= 16'b1111111111111110;
        weights1[47833] <= 16'b1111111111110010;
        weights1[47834] <= 16'b1111111111101101;
        weights1[47835] <= 16'b1111111111100101;
        weights1[47836] <= 16'b1111111111100100;
        weights1[47837] <= 16'b1111111111100001;
        weights1[47838] <= 16'b1111111111011101;
        weights1[47839] <= 16'b1111111111011110;
        weights1[47840] <= 16'b1111111111100010;
        weights1[47841] <= 16'b1111111111101001;
        weights1[47842] <= 16'b1111111111111000;
        weights1[47843] <= 16'b1111111111110010;
        weights1[47844] <= 16'b0000000000000100;
        weights1[47845] <= 16'b0000000000000110;
        weights1[47846] <= 16'b0000000000000000;
        weights1[47847] <= 16'b1111111111111010;
        weights1[47848] <= 16'b1111111111111110;
        weights1[47849] <= 16'b0000000000000100;
        weights1[47850] <= 16'b0000000000000111;
        weights1[47851] <= 16'b0000000000000101;
        weights1[47852] <= 16'b0000000000000000;
        weights1[47853] <= 16'b0000000000000000;
        weights1[47854] <= 16'b0000000000000001;
        weights1[47855] <= 16'b0000000000000010;
        weights1[47856] <= 16'b0000000000000100;
        weights1[47857] <= 16'b0000000000000011;
        weights1[47858] <= 16'b1111111111111100;
        weights1[47859] <= 16'b1111111111111010;
        weights1[47860] <= 16'b1111111111110101;
        weights1[47861] <= 16'b1111111111101010;
        weights1[47862] <= 16'b1111111111100011;
        weights1[47863] <= 16'b1111111111100110;
        weights1[47864] <= 16'b1111111111100101;
        weights1[47865] <= 16'b1111111111100011;
        weights1[47866] <= 16'b1111111111101010;
        weights1[47867] <= 16'b1111111111011011;
        weights1[47868] <= 16'b1111111111100011;
        weights1[47869] <= 16'b1111111111100010;
        weights1[47870] <= 16'b1111111111110010;
        weights1[47871] <= 16'b1111111111110101;
        weights1[47872] <= 16'b1111111111110101;
        weights1[47873] <= 16'b1111111111111110;
        weights1[47874] <= 16'b0000000000000101;
        weights1[47875] <= 16'b1111111111111111;
        weights1[47876] <= 16'b0000000000000000;
        weights1[47877] <= 16'b0000000000000111;
        weights1[47878] <= 16'b0000000000001000;
        weights1[47879] <= 16'b0000000000000110;
        weights1[47880] <= 16'b0000000000000000;
        weights1[47881] <= 16'b0000000000000100;
        weights1[47882] <= 16'b0000000000000100;
        weights1[47883] <= 16'b0000000000000011;
        weights1[47884] <= 16'b0000000000000010;
        weights1[47885] <= 16'b1111111111111111;
        weights1[47886] <= 16'b1111111111110111;
        weights1[47887] <= 16'b1111111111111010;
        weights1[47888] <= 16'b1111111111110000;
        weights1[47889] <= 16'b1111111111100100;
        weights1[47890] <= 16'b1111111111011010;
        weights1[47891] <= 16'b1111111111011010;
        weights1[47892] <= 16'b1111111111100011;
        weights1[47893] <= 16'b1111111111101000;
        weights1[47894] <= 16'b1111111111101000;
        weights1[47895] <= 16'b1111111111101111;
        weights1[47896] <= 16'b1111111111101111;
        weights1[47897] <= 16'b1111111111100101;
        weights1[47898] <= 16'b1111111111111101;
        weights1[47899] <= 16'b1111111111111101;
        weights1[47900] <= 16'b1111111111110101;
        weights1[47901] <= 16'b0000000000001001;
        weights1[47902] <= 16'b1111111111111101;
        weights1[47903] <= 16'b0000000000001100;
        weights1[47904] <= 16'b0000000000001011;
        weights1[47905] <= 16'b0000000000001100;
        weights1[47906] <= 16'b0000000000001101;
        weights1[47907] <= 16'b0000000000000110;
        weights1[47908] <= 16'b0000000000000000;
        weights1[47909] <= 16'b0000000000000010;
        weights1[47910] <= 16'b0000000000000011;
        weights1[47911] <= 16'b0000000000000000;
        weights1[47912] <= 16'b1111111111111111;
        weights1[47913] <= 16'b0000000000000000;
        weights1[47914] <= 16'b1111111111111101;
        weights1[47915] <= 16'b1111111111111100;
        weights1[47916] <= 16'b1111111111110000;
        weights1[47917] <= 16'b1111111111100100;
        weights1[47918] <= 16'b1111111111011001;
        weights1[47919] <= 16'b1111111111010111;
        weights1[47920] <= 16'b1111111111100111;
        weights1[47921] <= 16'b1111111111011110;
        weights1[47922] <= 16'b1111111111100001;
        weights1[47923] <= 16'b1111111111101011;
        weights1[47924] <= 16'b1111111111101101;
        weights1[47925] <= 16'b1111111111101001;
        weights1[47926] <= 16'b1111111111111101;
        weights1[47927] <= 16'b0000000000010001;
        weights1[47928] <= 16'b1111111111111101;
        weights1[47929] <= 16'b1111111111111101;
        weights1[47930] <= 16'b0000000000000110;
        weights1[47931] <= 16'b0000000000001101;
        weights1[47932] <= 16'b0000000000011000;
        weights1[47933] <= 16'b0000000000010100;
        weights1[47934] <= 16'b0000000000011011;
        weights1[47935] <= 16'b0000000000001100;
        weights1[47936] <= 16'b0000000000000001;
        weights1[47937] <= 16'b0000000000000001;
        weights1[47938] <= 16'b0000000000000010;
        weights1[47939] <= 16'b1111111111111011;
        weights1[47940] <= 16'b1111111111111000;
        weights1[47941] <= 16'b1111111111111010;
        weights1[47942] <= 16'b0000000000000000;
        weights1[47943] <= 16'b1111111111110010;
        weights1[47944] <= 16'b1111111111100000;
        weights1[47945] <= 16'b1111111111101001;
        weights1[47946] <= 16'b1111111111001000;
        weights1[47947] <= 16'b1111111111001001;
        weights1[47948] <= 16'b1111111110111110;
        weights1[47949] <= 16'b1111111111010100;
        weights1[47950] <= 16'b1111111111010110;
        weights1[47951] <= 16'b1111111111110010;
        weights1[47952] <= 16'b1111111111011101;
        weights1[47953] <= 16'b1111111111111100;
        weights1[47954] <= 16'b0000000000000000;
        weights1[47955] <= 16'b1111111111111101;
        weights1[47956] <= 16'b0000000000000111;
        weights1[47957] <= 16'b0000000000100011;
        weights1[47958] <= 16'b0000000000110111;
        weights1[47959] <= 16'b0000000000101101;
        weights1[47960] <= 16'b0000000000011011;
        weights1[47961] <= 16'b0000000000001011;
        weights1[47962] <= 16'b0000000000010010;
        weights1[47963] <= 16'b0000000000001010;
        weights1[47964] <= 16'b0000000000000001;
        weights1[47965] <= 16'b0000000000000001;
        weights1[47966] <= 16'b1111111111111100;
        weights1[47967] <= 16'b1111111111110101;
        weights1[47968] <= 16'b1111111111110011;
        weights1[47969] <= 16'b1111111111111100;
        weights1[47970] <= 16'b1111111111111011;
        weights1[47971] <= 16'b1111111111001011;
        weights1[47972] <= 16'b1111111111001010;
        weights1[47973] <= 16'b1111111110111111;
        weights1[47974] <= 16'b1111111110111110;
        weights1[47975] <= 16'b1111111111011101;
        weights1[47976] <= 16'b1111111111111111;
        weights1[47977] <= 16'b0000000000001011;
        weights1[47978] <= 16'b1111111111110111;
        weights1[47979] <= 16'b1111111111110000;
        weights1[47980] <= 16'b1111111111101111;
        weights1[47981] <= 16'b0000000000000111;
        weights1[47982] <= 16'b0000000000100000;
        weights1[47983] <= 16'b0000000000000011;
        weights1[47984] <= 16'b0000000000100000;
        weights1[47985] <= 16'b0000000000100100;
        weights1[47986] <= 16'b0000000000010101;
        weights1[47987] <= 16'b0000000000011110;
        weights1[47988] <= 16'b0000000000101011;
        weights1[47989] <= 16'b0000000000100000;
        weights1[47990] <= 16'b0000000000011110;
        weights1[47991] <= 16'b0000000000011001;
        weights1[47992] <= 16'b0000000000000000;
        weights1[47993] <= 16'b1111111111111111;
        weights1[47994] <= 16'b1111111111111010;
        weights1[47995] <= 16'b1111111111111001;
        weights1[47996] <= 16'b1111111111110111;
        weights1[47997] <= 16'b1111111111111101;
        weights1[47998] <= 16'b1111111111111100;
        weights1[47999] <= 16'b1111111111011100;
        weights1[48000] <= 16'b1111111110111001;
        weights1[48001] <= 16'b1111111110111001;
        weights1[48002] <= 16'b1111111111010101;
        weights1[48003] <= 16'b1111111110110101;
        weights1[48004] <= 16'b1111111111110111;
        weights1[48005] <= 16'b0000000000101100;
        weights1[48006] <= 16'b0000000000010111;
        weights1[48007] <= 16'b0000000000010010;
        weights1[48008] <= 16'b1111111111110111;
        weights1[48009] <= 16'b0000000000011100;
        weights1[48010] <= 16'b0000000000001010;
        weights1[48011] <= 16'b0000000000100010;
        weights1[48012] <= 16'b0000000000100011;
        weights1[48013] <= 16'b0000000000011101;
        weights1[48014] <= 16'b0000000000011011;
        weights1[48015] <= 16'b1111111111111011;
        weights1[48016] <= 16'b0000000000101000;
        weights1[48017] <= 16'b0000000000100011;
        weights1[48018] <= 16'b0000000000110111;
        weights1[48019] <= 16'b0000000000101010;
        weights1[48020] <= 16'b1111111111111111;
        weights1[48021] <= 16'b1111111111111110;
        weights1[48022] <= 16'b1111111111111001;
        weights1[48023] <= 16'b1111111111111011;
        weights1[48024] <= 16'b1111111111110111;
        weights1[48025] <= 16'b1111111111111101;
        weights1[48026] <= 16'b1111111111101000;
        weights1[48027] <= 16'b1111111111001101;
        weights1[48028] <= 16'b1111111111001111;
        weights1[48029] <= 16'b1111111110111110;
        weights1[48030] <= 16'b1111111111101000;
        weights1[48031] <= 16'b0000000000101100;
        weights1[48032] <= 16'b0000000000100011;
        weights1[48033] <= 16'b0000000000110100;
        weights1[48034] <= 16'b0000000000001011;
        weights1[48035] <= 16'b0000000000100000;
        weights1[48036] <= 16'b0000000000011010;
        weights1[48037] <= 16'b0000000000011011;
        weights1[48038] <= 16'b0000000000011001;
        weights1[48039] <= 16'b0000000000010001;
        weights1[48040] <= 16'b0000000000010010;
        weights1[48041] <= 16'b0000000000001100;
        weights1[48042] <= 16'b0000000000011111;
        weights1[48043] <= 16'b0000000000010110;
        weights1[48044] <= 16'b0000000000100111;
        weights1[48045] <= 16'b0000000000100001;
        weights1[48046] <= 16'b0000000000100100;
        weights1[48047] <= 16'b0000000000110010;
        weights1[48048] <= 16'b1111111111111110;
        weights1[48049] <= 16'b1111111111111100;
        weights1[48050] <= 16'b0000000000000000;
        weights1[48051] <= 16'b1111111111110100;
        weights1[48052] <= 16'b1111111111101100;
        weights1[48053] <= 16'b1111111111101011;
        weights1[48054] <= 16'b1111111111010011;
        weights1[48055] <= 16'b1111111110101111;
        weights1[48056] <= 16'b1111111110011011;
        weights1[48057] <= 16'b1111111111010110;
        weights1[48058] <= 16'b1111111111101101;
        weights1[48059] <= 16'b0000000000101010;
        weights1[48060] <= 16'b0000000000110111;
        weights1[48061] <= 16'b0000000000011111;
        weights1[48062] <= 16'b0000000000110011;
        weights1[48063] <= 16'b0000000000001111;
        weights1[48064] <= 16'b0000000000101111;
        weights1[48065] <= 16'b0000000000100000;
        weights1[48066] <= 16'b0000000000001011;
        weights1[48067] <= 16'b0000000000011000;
        weights1[48068] <= 16'b0000000000011011;
        weights1[48069] <= 16'b0000000000001111;
        weights1[48070] <= 16'b0000000000001101;
        weights1[48071] <= 16'b0000000001000110;
        weights1[48072] <= 16'b0000000000101010;
        weights1[48073] <= 16'b0000000000100110;
        weights1[48074] <= 16'b0000000000010100;
        weights1[48075] <= 16'b0000000000100111;
        weights1[48076] <= 16'b1111111111111100;
        weights1[48077] <= 16'b1111111111111010;
        weights1[48078] <= 16'b1111111111111010;
        weights1[48079] <= 16'b1111111111110011;
        weights1[48080] <= 16'b1111111111101010;
        weights1[48081] <= 16'b1111111111100011;
        weights1[48082] <= 16'b1111111111000001;
        weights1[48083] <= 16'b1111111110110001;
        weights1[48084] <= 16'b1111111111000100;
        weights1[48085] <= 16'b1111111111101101;
        weights1[48086] <= 16'b0000000000000010;
        weights1[48087] <= 16'b0000000000011110;
        weights1[48088] <= 16'b0000000000101001;
        weights1[48089] <= 16'b0000000001001111;
        weights1[48090] <= 16'b0000000000110110;
        weights1[48091] <= 16'b0000000000001011;
        weights1[48092] <= 16'b1111111111110100;
        weights1[48093] <= 16'b0000000000101001;
        weights1[48094] <= 16'b0000000000110011;
        weights1[48095] <= 16'b0000000000010000;
        weights1[48096] <= 16'b0000000000010100;
        weights1[48097] <= 16'b0000000000011100;
        weights1[48098] <= 16'b1111111111111100;
        weights1[48099] <= 16'b0000000000001011;
        weights1[48100] <= 16'b0000000000010111;
        weights1[48101] <= 16'b0000000000011100;
        weights1[48102] <= 16'b0000000000000111;
        weights1[48103] <= 16'b0000000000101110;
        weights1[48104] <= 16'b1111111111111010;
        weights1[48105] <= 16'b1111111111111011;
        weights1[48106] <= 16'b1111111111111100;
        weights1[48107] <= 16'b1111111111110000;
        weights1[48108] <= 16'b1111111111101100;
        weights1[48109] <= 16'b1111111111010101;
        weights1[48110] <= 16'b1111111110111010;
        weights1[48111] <= 16'b1111111111001001;
        weights1[48112] <= 16'b1111111111100110;
        weights1[48113] <= 16'b0000000000000101;
        weights1[48114] <= 16'b0000000000001010;
        weights1[48115] <= 16'b0000000000111011;
        weights1[48116] <= 16'b0000000000110101;
        weights1[48117] <= 16'b0000000000111011;
        weights1[48118] <= 16'b0000000000001010;
        weights1[48119] <= 16'b1111111111101010;
        weights1[48120] <= 16'b1111111111011110;
        weights1[48121] <= 16'b1111111111101110;
        weights1[48122] <= 16'b1111111111110001;
        weights1[48123] <= 16'b1111111111010001;
        weights1[48124] <= 16'b1111111111110101;
        weights1[48125] <= 16'b1111111111011111;
        weights1[48126] <= 16'b1111111111100111;
        weights1[48127] <= 16'b1111111111100111;
        weights1[48128] <= 16'b1111111111101011;
        weights1[48129] <= 16'b0000000000000011;
        weights1[48130] <= 16'b0000000000001101;
        weights1[48131] <= 16'b0000000000000110;
        weights1[48132] <= 16'b1111111111111010;
        weights1[48133] <= 16'b1111111111111100;
        weights1[48134] <= 16'b1111111111111001;
        weights1[48135] <= 16'b1111111111101110;
        weights1[48136] <= 16'b1111111111100101;
        weights1[48137] <= 16'b1111111111010110;
        weights1[48138] <= 16'b1111111110111111;
        weights1[48139] <= 16'b1111111111001011;
        weights1[48140] <= 16'b1111111111111000;
        weights1[48141] <= 16'b1111111111111110;
        weights1[48142] <= 16'b0000000000010010;
        weights1[48143] <= 16'b0000000000000110;
        weights1[48144] <= 16'b0000000001001000;
        weights1[48145] <= 16'b0000000000111110;
        weights1[48146] <= 16'b1111111111101110;
        weights1[48147] <= 16'b1111111110011111;
        weights1[48148] <= 16'b1111111110100000;
        weights1[48149] <= 16'b1111111111000000;
        weights1[48150] <= 16'b1111111111110101;
        weights1[48151] <= 16'b1111111111110100;
        weights1[48152] <= 16'b1111111111010110;
        weights1[48153] <= 16'b1111111111100010;
        weights1[48154] <= 16'b1111111111101001;
        weights1[48155] <= 16'b1111111111100100;
        weights1[48156] <= 16'b1111111111101010;
        weights1[48157] <= 16'b0000000000000110;
        weights1[48158] <= 16'b0000000000000001;
        weights1[48159] <= 16'b1111111111111101;
        weights1[48160] <= 16'b1111111111111011;
        weights1[48161] <= 16'b1111111111111111;
        weights1[48162] <= 16'b1111111111111101;
        weights1[48163] <= 16'b1111111111100110;
        weights1[48164] <= 16'b1111111111010001;
        weights1[48165] <= 16'b1111111111000111;
        weights1[48166] <= 16'b1111111111010110;
        weights1[48167] <= 16'b1111111111010011;
        weights1[48168] <= 16'b0000000000010000;
        weights1[48169] <= 16'b1111111111111001;
        weights1[48170] <= 16'b0000000000100101;
        weights1[48171] <= 16'b0000000000100111;
        weights1[48172] <= 16'b0000000000100011;
        weights1[48173] <= 16'b0000000001000011;
        weights1[48174] <= 16'b1111111111101001;
        weights1[48175] <= 16'b1111111110010011;
        weights1[48176] <= 16'b1111111110101010;
        weights1[48177] <= 16'b1111111111100111;
        weights1[48178] <= 16'b1111111111110100;
        weights1[48179] <= 16'b1111111111101010;
        weights1[48180] <= 16'b1111111111101100;
        weights1[48181] <= 16'b1111111111011101;
        weights1[48182] <= 16'b1111111111011111;
        weights1[48183] <= 16'b1111111111100010;
        weights1[48184] <= 16'b1111111111111101;
        weights1[48185] <= 16'b1111111111110110;
        weights1[48186] <= 16'b1111111111110100;
        weights1[48187] <= 16'b0000000000000100;
        weights1[48188] <= 16'b1111111111111010;
        weights1[48189] <= 16'b1111111111110111;
        weights1[48190] <= 16'b1111111111110111;
        weights1[48191] <= 16'b1111111111100000;
        weights1[48192] <= 16'b1111111111001101;
        weights1[48193] <= 16'b1111111111101001;
        weights1[48194] <= 16'b0000000000000001;
        weights1[48195] <= 16'b1111111111101110;
        weights1[48196] <= 16'b0000000000001011;
        weights1[48197] <= 16'b1111111111111111;
        weights1[48198] <= 16'b0000000000011111;
        weights1[48199] <= 16'b0000000000010001;
        weights1[48200] <= 16'b0000000000111010;
        weights1[48201] <= 16'b0000000000011111;
        weights1[48202] <= 16'b1111111110111110;
        weights1[48203] <= 16'b1111111110000101;
        weights1[48204] <= 16'b1111111111000110;
        weights1[48205] <= 16'b1111111111011001;
        weights1[48206] <= 16'b1111111111011100;
        weights1[48207] <= 16'b1111111111101011;
        weights1[48208] <= 16'b1111111111101111;
        weights1[48209] <= 16'b1111111111100010;
        weights1[48210] <= 16'b1111111111101011;
        weights1[48211] <= 16'b1111111111110000;
        weights1[48212] <= 16'b0000000000000100;
        weights1[48213] <= 16'b1111111111110100;
        weights1[48214] <= 16'b0000000000010011;
        weights1[48215] <= 16'b0000000000011000;
        weights1[48216] <= 16'b1111111111110111;
        weights1[48217] <= 16'b1111111111110010;
        weights1[48218] <= 16'b1111111111110011;
        weights1[48219] <= 16'b1111111111101111;
        weights1[48220] <= 16'b1111111111001100;
        weights1[48221] <= 16'b1111111111101111;
        weights1[48222] <= 16'b1111111111011110;
        weights1[48223] <= 16'b1111111111111111;
        weights1[48224] <= 16'b0000000000001000;
        weights1[48225] <= 16'b0000000000100110;
        weights1[48226] <= 16'b0000000000101011;
        weights1[48227] <= 16'b0000000000000010;
        weights1[48228] <= 16'b0000000000001110;
        weights1[48229] <= 16'b1111111111101011;
        weights1[48230] <= 16'b1111111110100001;
        weights1[48231] <= 16'b1111111110011110;
        weights1[48232] <= 16'b1111111111000011;
        weights1[48233] <= 16'b1111111111101001;
        weights1[48234] <= 16'b1111111111110011;
        weights1[48235] <= 16'b1111111111100111;
        weights1[48236] <= 16'b1111111111010101;
        weights1[48237] <= 16'b1111111111110010;
        weights1[48238] <= 16'b0000000000000010;
        weights1[48239] <= 16'b1111111111100011;
        weights1[48240] <= 16'b1111111111111101;
        weights1[48241] <= 16'b0000000000010001;
        weights1[48242] <= 16'b0000000000011100;
        weights1[48243] <= 16'b0000000000010011;
        weights1[48244] <= 16'b1111111111110001;
        weights1[48245] <= 16'b1111111111101111;
        weights1[48246] <= 16'b1111111111101111;
        weights1[48247] <= 16'b1111111111101000;
        weights1[48248] <= 16'b1111111111010111;
        weights1[48249] <= 16'b0000000000000011;
        weights1[48250] <= 16'b1111111111101001;
        weights1[48251] <= 16'b0000000000001010;
        weights1[48252] <= 16'b1111111111110100;
        weights1[48253] <= 16'b0000000000010100;
        weights1[48254] <= 16'b0000000000001101;
        weights1[48255] <= 16'b0000000000000000;
        weights1[48256] <= 16'b0000000000000010;
        weights1[48257] <= 16'b1111111111001111;
        weights1[48258] <= 16'b1111111110001001;
        weights1[48259] <= 16'b1111111110110111;
        weights1[48260] <= 16'b1111111111010100;
        weights1[48261] <= 16'b1111111111011101;
        weights1[48262] <= 16'b1111111111101010;
        weights1[48263] <= 16'b1111111111010111;
        weights1[48264] <= 16'b0000000000000000;
        weights1[48265] <= 16'b1111111111110111;
        weights1[48266] <= 16'b1111111111100011;
        weights1[48267] <= 16'b0000000000000000;
        weights1[48268] <= 16'b1111111111101001;
        weights1[48269] <= 16'b0000000000010000;
        weights1[48270] <= 16'b1111111111111010;
        weights1[48271] <= 16'b0000000000001011;
        weights1[48272] <= 16'b1111111111110100;
        weights1[48273] <= 16'b1111111111111010;
        weights1[48274] <= 16'b1111111111101011;
        weights1[48275] <= 16'b1111111111100001;
        weights1[48276] <= 16'b1111111111011111;
        weights1[48277] <= 16'b1111111111111101;
        weights1[48278] <= 16'b1111111111101111;
        weights1[48279] <= 16'b1111111111100101;
        weights1[48280] <= 16'b1111111111111101;
        weights1[48281] <= 16'b0000000000000010;
        weights1[48282] <= 16'b0000000000001000;
        weights1[48283] <= 16'b0000000000001110;
        weights1[48284] <= 16'b1111111111100000;
        weights1[48285] <= 16'b1111111110110010;
        weights1[48286] <= 16'b1111111110110000;
        weights1[48287] <= 16'b1111111111000011;
        weights1[48288] <= 16'b1111111111001111;
        weights1[48289] <= 16'b1111111111100101;
        weights1[48290] <= 16'b1111111111111011;
        weights1[48291] <= 16'b1111111111111011;
        weights1[48292] <= 16'b1111111111101110;
        weights1[48293] <= 16'b0000000000001101;
        weights1[48294] <= 16'b0000000000001000;
        weights1[48295] <= 16'b1111111111111110;
        weights1[48296] <= 16'b0000000000000110;
        weights1[48297] <= 16'b0000000000000001;
        weights1[48298] <= 16'b0000000000000111;
        weights1[48299] <= 16'b0000000000000000;
        weights1[48300] <= 16'b1111111111111010;
        weights1[48301] <= 16'b1111111111110111;
        weights1[48302] <= 16'b1111111111101111;
        weights1[48303] <= 16'b1111111111100011;
        weights1[48304] <= 16'b1111111111011011;
        weights1[48305] <= 16'b1111111111111110;
        weights1[48306] <= 16'b1111111111111100;
        weights1[48307] <= 16'b1111111111110001;
        weights1[48308] <= 16'b1111111111110010;
        weights1[48309] <= 16'b1111111111001111;
        weights1[48310] <= 16'b1111111111110011;
        weights1[48311] <= 16'b0000000000000010;
        weights1[48312] <= 16'b1111111111010100;
        weights1[48313] <= 16'b1111111111001101;
        weights1[48314] <= 16'b1111111110111000;
        weights1[48315] <= 16'b1111111111011111;
        weights1[48316] <= 16'b1111111111101111;
        weights1[48317] <= 16'b1111111111111001;
        weights1[48318] <= 16'b0000000000010110;
        weights1[48319] <= 16'b1111111111111111;
        weights1[48320] <= 16'b0000000000001000;
        weights1[48321] <= 16'b1111111111111010;
        weights1[48322] <= 16'b0000000000000011;
        weights1[48323] <= 16'b0000000000000010;
        weights1[48324] <= 16'b1111111111111001;
        weights1[48325] <= 16'b0000000000000011;
        weights1[48326] <= 16'b0000000000001010;
        weights1[48327] <= 16'b0000000000001010;
        weights1[48328] <= 16'b1111111111111111;
        weights1[48329] <= 16'b0000000000000000;
        weights1[48330] <= 16'b1111111111111100;
        weights1[48331] <= 16'b1111111111110010;
        weights1[48332] <= 16'b1111111111101100;
        weights1[48333] <= 16'b1111111111111000;
        weights1[48334] <= 16'b0000000000010111;
        weights1[48335] <= 16'b1111111111111101;
        weights1[48336] <= 16'b1111111111111000;
        weights1[48337] <= 16'b1111111111111100;
        weights1[48338] <= 16'b1111111111110000;
        weights1[48339] <= 16'b1111111111110101;
        weights1[48340] <= 16'b1111111111001011;
        weights1[48341] <= 16'b1111111111101110;
        weights1[48342] <= 16'b1111111111001010;
        weights1[48343] <= 16'b1111111111110001;
        weights1[48344] <= 16'b0000000000001011;
        weights1[48345] <= 16'b1111111111111111;
        weights1[48346] <= 16'b1111111111101010;
        weights1[48347] <= 16'b1111111111111010;
        weights1[48348] <= 16'b0000000000000001;
        weights1[48349] <= 16'b1111111111100011;
        weights1[48350] <= 16'b0000000000000110;
        weights1[48351] <= 16'b1111111111110111;
        weights1[48352] <= 16'b1111111111110011;
        weights1[48353] <= 16'b0000000000001111;
        weights1[48354] <= 16'b1111111111111101;
        weights1[48355] <= 16'b0000000000000101;
        weights1[48356] <= 16'b0000000000000011;
        weights1[48357] <= 16'b0000000000000111;
        weights1[48358] <= 16'b0000000000000110;
        weights1[48359] <= 16'b1111111111100110;
        weights1[48360] <= 16'b1111111111111010;
        weights1[48361] <= 16'b1111111111111111;
        weights1[48362] <= 16'b0000000000010111;
        weights1[48363] <= 16'b0000000000100111;
        weights1[48364] <= 16'b1111111111101111;
        weights1[48365] <= 16'b0000000000000101;
        weights1[48366] <= 16'b1111111111111111;
        weights1[48367] <= 16'b0000000000001100;
        weights1[48368] <= 16'b1111111111111000;
        weights1[48369] <= 16'b1111111111111100;
        weights1[48370] <= 16'b0000000000010100;
        weights1[48371] <= 16'b1111111111110111;
        weights1[48372] <= 16'b1111111111110101;
        weights1[48373] <= 16'b1111111111110011;
        weights1[48374] <= 16'b0000000000001110;
        weights1[48375] <= 16'b1111111111110111;
        weights1[48376] <= 16'b0000000000010010;
        weights1[48377] <= 16'b1111111111110100;
        weights1[48378] <= 16'b0000000000000001;
        weights1[48379] <= 16'b0000000000000010;
        weights1[48380] <= 16'b0000000000000010;
        weights1[48381] <= 16'b1111111111111111;
        weights1[48382] <= 16'b1111111111110110;
        weights1[48383] <= 16'b1111111111110111;
        weights1[48384] <= 16'b0000000000000000;
        weights1[48385] <= 16'b0000000000001110;
        weights1[48386] <= 16'b0000000000000010;
        weights1[48387] <= 16'b1111111111011011;
        weights1[48388] <= 16'b0000000000000110;
        weights1[48389] <= 16'b0000000000000001;
        weights1[48390] <= 16'b0000000000100000;
        weights1[48391] <= 16'b1111111111110101;
        weights1[48392] <= 16'b0000000000010101;
        weights1[48393] <= 16'b0000000000001010;
        weights1[48394] <= 16'b0000000000010111;
        weights1[48395] <= 16'b0000000000000110;
        weights1[48396] <= 16'b0000000000000010;
        weights1[48397] <= 16'b1111111111111110;
        weights1[48398] <= 16'b1111111111011101;
        weights1[48399] <= 16'b0000000000000101;
        weights1[48400] <= 16'b0000000000000001;
        weights1[48401] <= 16'b1111111111110010;
        weights1[48402] <= 16'b0000000000001101;
        weights1[48403] <= 16'b0000000000001001;
        weights1[48404] <= 16'b1111111111111011;
        weights1[48405] <= 16'b0000000000000100;
        weights1[48406] <= 16'b1111111111110100;
        weights1[48407] <= 16'b1111111111101011;
        weights1[48408] <= 16'b1111111111110110;
        weights1[48409] <= 16'b1111111111110011;
        weights1[48410] <= 16'b1111111111110001;
        weights1[48411] <= 16'b1111111111101111;
        weights1[48412] <= 16'b1111111111111101;
        weights1[48413] <= 16'b0000000000000010;
        weights1[48414] <= 16'b1111111111111101;
        weights1[48415] <= 16'b1111111111101011;
        weights1[48416] <= 16'b1111111111110110;
        weights1[48417] <= 16'b1111111111101000;
        weights1[48418] <= 16'b1111111111100111;
        weights1[48419] <= 16'b1111111111111101;
        weights1[48420] <= 16'b0000000000010100;
        weights1[48421] <= 16'b0000000000000100;
        weights1[48422] <= 16'b1111111111111100;
        weights1[48423] <= 16'b0000000000011000;
        weights1[48424] <= 16'b0000000000000111;
        weights1[48425] <= 16'b0000000000000110;
        weights1[48426] <= 16'b1111111111111010;
        weights1[48427] <= 16'b1111111111111000;
        weights1[48428] <= 16'b1111111111111100;
        weights1[48429] <= 16'b1111111111110000;
        weights1[48430] <= 16'b0000000000010001;
        weights1[48431] <= 16'b0000000000000001;
        weights1[48432] <= 16'b1111111111110011;
        weights1[48433] <= 16'b1111111111111100;
        weights1[48434] <= 16'b1111111111111101;
        weights1[48435] <= 16'b1111111111100100;
        weights1[48436] <= 16'b1111111111110000;
        weights1[48437] <= 16'b1111111111101111;
        weights1[48438] <= 16'b1111111111110110;
        weights1[48439] <= 16'b1111111111101101;
        weights1[48440] <= 16'b1111111111111101;
        weights1[48441] <= 16'b1111111111111101;
        weights1[48442] <= 16'b1111111111110100;
        weights1[48443] <= 16'b1111111111100110;
        weights1[48444] <= 16'b1111111111101000;
        weights1[48445] <= 16'b1111111111011100;
        weights1[48446] <= 16'b1111111111110111;
        weights1[48447] <= 16'b1111111111101111;
        weights1[48448] <= 16'b0000000000001000;
        weights1[48449] <= 16'b0000000000000001;
        weights1[48450] <= 16'b0000000000001000;
        weights1[48451] <= 16'b0000000000001011;
        weights1[48452] <= 16'b0000000000001110;
        weights1[48453] <= 16'b1111111111101100;
        weights1[48454] <= 16'b0000000000000111;
        weights1[48455] <= 16'b0000000000000111;
        weights1[48456] <= 16'b0000000000001010;
        weights1[48457] <= 16'b0000000000001101;
        weights1[48458] <= 16'b0000000000001010;
        weights1[48459] <= 16'b1111111111111001;
        weights1[48460] <= 16'b1111111111111100;
        weights1[48461] <= 16'b1111111111110010;
        weights1[48462] <= 16'b1111111111110011;
        weights1[48463] <= 16'b1111111111011111;
        weights1[48464] <= 16'b1111111111101100;
        weights1[48465] <= 16'b1111111111101100;
        weights1[48466] <= 16'b1111111111110000;
        weights1[48467] <= 16'b1111111111110010;
        weights1[48468] <= 16'b0000000000000000;
        weights1[48469] <= 16'b1111111111111101;
        weights1[48470] <= 16'b1111111111110110;
        weights1[48471] <= 16'b1111111111100110;
        weights1[48472] <= 16'b1111111111110000;
        weights1[48473] <= 16'b1111111111110101;
        weights1[48474] <= 16'b0000000000001101;
        weights1[48475] <= 16'b1111111111110100;
        weights1[48476] <= 16'b1111111111011100;
        weights1[48477] <= 16'b1111111111100100;
        weights1[48478] <= 16'b0000000000100001;
        weights1[48479] <= 16'b0000000000001101;
        weights1[48480] <= 16'b1111111111111101;
        weights1[48481] <= 16'b0000000000001110;
        weights1[48482] <= 16'b0000000000011001;
        weights1[48483] <= 16'b1111111111110010;
        weights1[48484] <= 16'b0000000000010010;
        weights1[48485] <= 16'b1111111111110001;
        weights1[48486] <= 16'b1111111111011111;
        weights1[48487] <= 16'b1111111111110101;
        weights1[48488] <= 16'b1111111111111111;
        weights1[48489] <= 16'b1111111111111001;
        weights1[48490] <= 16'b1111111111101010;
        weights1[48491] <= 16'b1111111111110001;
        weights1[48492] <= 16'b1111111111101001;
        weights1[48493] <= 16'b1111111111101111;
        weights1[48494] <= 16'b1111111111101101;
        weights1[48495] <= 16'b1111111111110001;
        weights1[48496] <= 16'b1111111111111110;
        weights1[48497] <= 16'b1111111111111011;
        weights1[48498] <= 16'b0000000000000001;
        weights1[48499] <= 16'b1111111111110100;
        weights1[48500] <= 16'b1111111111101100;
        weights1[48501] <= 16'b1111111111011110;
        weights1[48502] <= 16'b1111111111110101;
        weights1[48503] <= 16'b1111111111101101;
        weights1[48504] <= 16'b1111111111111001;
        weights1[48505] <= 16'b0000000000000100;
        weights1[48506] <= 16'b1111111111110011;
        weights1[48507] <= 16'b1111111111011111;
        weights1[48508] <= 16'b0000000000001101;
        weights1[48509] <= 16'b1111111111111010;
        weights1[48510] <= 16'b1111111111110110;
        weights1[48511] <= 16'b0000000000010110;
        weights1[48512] <= 16'b1111111111101101;
        weights1[48513] <= 16'b0000000000001111;
        weights1[48514] <= 16'b0000000000000010;
        weights1[48515] <= 16'b1111111111111100;
        weights1[48516] <= 16'b1111111111011100;
        weights1[48517] <= 16'b1111111111101110;
        weights1[48518] <= 16'b1111111111100101;
        weights1[48519] <= 16'b1111111111100100;
        weights1[48520] <= 16'b1111111111100011;
        weights1[48521] <= 16'b1111111111101011;
        weights1[48522] <= 16'b1111111111110001;
        weights1[48523] <= 16'b1111111111110101;
        weights1[48524] <= 16'b1111111111111111;
        weights1[48525] <= 16'b1111111111111101;
        weights1[48526] <= 16'b1111111111111100;
        weights1[48527] <= 16'b1111111111111001;
        weights1[48528] <= 16'b1111111111110101;
        weights1[48529] <= 16'b1111111111100000;
        weights1[48530] <= 16'b0000000000000100;
        weights1[48531] <= 16'b0000000000001011;
        weights1[48532] <= 16'b1111111111111110;
        weights1[48533] <= 16'b0000000000000010;
        weights1[48534] <= 16'b1111111111110010;
        weights1[48535] <= 16'b0000000000010010;
        weights1[48536] <= 16'b0000000000001010;
        weights1[48537] <= 16'b0000000000001001;
        weights1[48538] <= 16'b1111111111011100;
        weights1[48539] <= 16'b1111111111111001;
        weights1[48540] <= 16'b1111111111100011;
        weights1[48541] <= 16'b1111111111110111;
        weights1[48542] <= 16'b1111111111101001;
        weights1[48543] <= 16'b1111111111110010;
        weights1[48544] <= 16'b1111111111011111;
        weights1[48545] <= 16'b1111111111100000;
        weights1[48546] <= 16'b1111111111011000;
        weights1[48547] <= 16'b1111111111101001;
        weights1[48548] <= 16'b1111111111101000;
        weights1[48549] <= 16'b1111111111110000;
        weights1[48550] <= 16'b1111111111110001;
        weights1[48551] <= 16'b1111111111111011;
        weights1[48552] <= 16'b1111111111111111;
        weights1[48553] <= 16'b1111111111111100;
        weights1[48554] <= 16'b1111111111111000;
        weights1[48555] <= 16'b1111111111111010;
        weights1[48556] <= 16'b0000000000000001;
        weights1[48557] <= 16'b1111111111110111;
        weights1[48558] <= 16'b0000000000000001;
        weights1[48559] <= 16'b0000000000011010;
        weights1[48560] <= 16'b0000000000100100;
        weights1[48561] <= 16'b0000000000001100;
        weights1[48562] <= 16'b1111111111110010;
        weights1[48563] <= 16'b0000000000000110;
        weights1[48564] <= 16'b0000000000001010;
        weights1[48565] <= 16'b0000000000000000;
        weights1[48566] <= 16'b0000000000000101;
        weights1[48567] <= 16'b1111111111111010;
        weights1[48568] <= 16'b1111111111101110;
        weights1[48569] <= 16'b1111111111100000;
        weights1[48570] <= 16'b1111111111110000;
        weights1[48571] <= 16'b1111111111100101;
        weights1[48572] <= 16'b1111111111100111;
        weights1[48573] <= 16'b1111111111101000;
        weights1[48574] <= 16'b1111111111101001;
        weights1[48575] <= 16'b1111111111100100;
        weights1[48576] <= 16'b1111111111101101;
        weights1[48577] <= 16'b1111111111110011;
        weights1[48578] <= 16'b1111111111111000;
        weights1[48579] <= 16'b1111111111111100;
        weights1[48580] <= 16'b1111111111111111;
        weights1[48581] <= 16'b1111111111111110;
        weights1[48582] <= 16'b1111111111111010;
        weights1[48583] <= 16'b1111111111111101;
        weights1[48584] <= 16'b1111111111111100;
        weights1[48585] <= 16'b1111111111110100;
        weights1[48586] <= 16'b1111111111110011;
        weights1[48587] <= 16'b1111111111110011;
        weights1[48588] <= 16'b1111111111111100;
        weights1[48589] <= 16'b1111111111100111;
        weights1[48590] <= 16'b1111111111101110;
        weights1[48591] <= 16'b1111111111101111;
        weights1[48592] <= 16'b1111111111111000;
        weights1[48593] <= 16'b1111111111101110;
        weights1[48594] <= 16'b1111111111110011;
        weights1[48595] <= 16'b1111111111000011;
        weights1[48596] <= 16'b1111111111000111;
        weights1[48597] <= 16'b1111111111000111;
        weights1[48598] <= 16'b1111111111001100;
        weights1[48599] <= 16'b1111111111011101;
        weights1[48600] <= 16'b1111111111101001;
        weights1[48601] <= 16'b1111111111011010;
        weights1[48602] <= 16'b1111111111101010;
        weights1[48603] <= 16'b1111111111101111;
        weights1[48604] <= 16'b1111111111110010;
        weights1[48605] <= 16'b1111111111111101;
        weights1[48606] <= 16'b1111111111111110;
        weights1[48607] <= 16'b1111111111111110;
        weights1[48608] <= 16'b0000000000000001;
        weights1[48609] <= 16'b1111111111111111;
        weights1[48610] <= 16'b1111111111111111;
        weights1[48611] <= 16'b1111111111111101;
        weights1[48612] <= 16'b1111111111111011;
        weights1[48613] <= 16'b1111111111111011;
        weights1[48614] <= 16'b0000000000000111;
        weights1[48615] <= 16'b0000000000000100;
        weights1[48616] <= 16'b0000000000000101;
        weights1[48617] <= 16'b0000000000001000;
        weights1[48618] <= 16'b0000000000010001;
        weights1[48619] <= 16'b0000000000001100;
        weights1[48620] <= 16'b0000000000000011;
        weights1[48621] <= 16'b1111111111111110;
        weights1[48622] <= 16'b0000000000000000;
        weights1[48623] <= 16'b1111111111111101;
        weights1[48624] <= 16'b0000000000000000;
        weights1[48625] <= 16'b0000000000001101;
        weights1[48626] <= 16'b1111111111111101;
        weights1[48627] <= 16'b0000000000001011;
        weights1[48628] <= 16'b0000000000010101;
        weights1[48629] <= 16'b0000000000010000;
        weights1[48630] <= 16'b1111111111111111;
        weights1[48631] <= 16'b0000000000000011;
        weights1[48632] <= 16'b1111111111111111;
        weights1[48633] <= 16'b1111111111110011;
        weights1[48634] <= 16'b1111111111111001;
        weights1[48635] <= 16'b0000000000000001;
        weights1[48636] <= 16'b0000000000000001;
        weights1[48637] <= 16'b0000000000000000;
        weights1[48638] <= 16'b1111111111111001;
        weights1[48639] <= 16'b1111111111111100;
        weights1[48640] <= 16'b1111111111111110;
        weights1[48641] <= 16'b1111111111111111;
        weights1[48642] <= 16'b1111111111110001;
        weights1[48643] <= 16'b0000000000000001;
        weights1[48644] <= 16'b1111111111101110;
        weights1[48645] <= 16'b0000000000000010;
        weights1[48646] <= 16'b1111111111111010;
        weights1[48647] <= 16'b1111111111111010;
        weights1[48648] <= 16'b1111111111111101;
        weights1[48649] <= 16'b0000000000000000;
        weights1[48650] <= 16'b1111111111110010;
        weights1[48651] <= 16'b0000000000000111;
        weights1[48652] <= 16'b1111111111110101;
        weights1[48653] <= 16'b1111111111111011;
        weights1[48654] <= 16'b1111111111111101;
        weights1[48655] <= 16'b1111111111110111;
        weights1[48656] <= 16'b0000000000000011;
        weights1[48657] <= 16'b1111111111111011;
        weights1[48658] <= 16'b1111111111110110;
        weights1[48659] <= 16'b1111111111111110;
        weights1[48660] <= 16'b1111111111111110;
        weights1[48661] <= 16'b0000000000000001;
        weights1[48662] <= 16'b1111111111111111;
        weights1[48663] <= 16'b1111111111111110;
        weights1[48664] <= 16'b0000000000000010;
        weights1[48665] <= 16'b1111111111111101;
        weights1[48666] <= 16'b1111111111111001;
        weights1[48667] <= 16'b1111111111110100;
        weights1[48668] <= 16'b1111111111111011;
        weights1[48669] <= 16'b1111111111110010;
        weights1[48670] <= 16'b1111111111110000;
        weights1[48671] <= 16'b1111111111111011;
        weights1[48672] <= 16'b1111111111101110;
        weights1[48673] <= 16'b0000000000000101;
        weights1[48674] <= 16'b1111111111111000;
        weights1[48675] <= 16'b0000000000000000;
        weights1[48676] <= 16'b1111111111111100;
        weights1[48677] <= 16'b1111111111111000;
        weights1[48678] <= 16'b0000000000000001;
        weights1[48679] <= 16'b0000000000010001;
        weights1[48680] <= 16'b1111111111111111;
        weights1[48681] <= 16'b0000000000000100;
        weights1[48682] <= 16'b1111111111110111;
        weights1[48683] <= 16'b0000000000001010;
        weights1[48684] <= 16'b1111111111111101;
        weights1[48685] <= 16'b0000000000000100;
        weights1[48686] <= 16'b1111111111111010;
        weights1[48687] <= 16'b0000000000000111;
        weights1[48688] <= 16'b0000000000001100;
        weights1[48689] <= 16'b0000000000001000;
        weights1[48690] <= 16'b0000000000000101;
        weights1[48691] <= 16'b0000000000000011;
        weights1[48692] <= 16'b0000000000000011;
        weights1[48693] <= 16'b0000000000000011;
        weights1[48694] <= 16'b1111111111110110;
        weights1[48695] <= 16'b1111111111111001;
        weights1[48696] <= 16'b1111111111111111;
        weights1[48697] <= 16'b1111111111110111;
        weights1[48698] <= 16'b1111111111111100;
        weights1[48699] <= 16'b0000000000000001;
        weights1[48700] <= 16'b0000000000001100;
        weights1[48701] <= 16'b1111111111111111;
        weights1[48702] <= 16'b0000000000001001;
        weights1[48703] <= 16'b0000000000000011;
        weights1[48704] <= 16'b1111111111111011;
        weights1[48705] <= 16'b1111111111111110;
        weights1[48706] <= 16'b1111111111110110;
        weights1[48707] <= 16'b1111111111110101;
        weights1[48708] <= 16'b1111111111111110;
        weights1[48709] <= 16'b0000000000000101;
        weights1[48710] <= 16'b1111111111110010;
        weights1[48711] <= 16'b1111111111111100;
        weights1[48712] <= 16'b0000000000000010;
        weights1[48713] <= 16'b0000000000000011;
        weights1[48714] <= 16'b0000000000000001;
        weights1[48715] <= 16'b0000000000001101;
        weights1[48716] <= 16'b0000000000010001;
        weights1[48717] <= 16'b0000000000000101;
        weights1[48718] <= 16'b0000000000001110;
        weights1[48719] <= 16'b0000000000001100;
        weights1[48720] <= 16'b1111111111111110;
        weights1[48721] <= 16'b1111111111111100;
        weights1[48722] <= 16'b1111111111111101;
        weights1[48723] <= 16'b0000000000000001;
        weights1[48724] <= 16'b1111111111111110;
        weights1[48725] <= 16'b1111111111111100;
        weights1[48726] <= 16'b0000000000000000;
        weights1[48727] <= 16'b0000000000001011;
        weights1[48728] <= 16'b1111111111111001;
        weights1[48729] <= 16'b1111111111101111;
        weights1[48730] <= 16'b0000000000000010;
        weights1[48731] <= 16'b0000000000000110;
        weights1[48732] <= 16'b0000000000000001;
        weights1[48733] <= 16'b1111111111111100;
        weights1[48734] <= 16'b0000000000001100;
        weights1[48735] <= 16'b0000000000001110;
        weights1[48736] <= 16'b1111111111110011;
        weights1[48737] <= 16'b0000000000001110;
        weights1[48738] <= 16'b0000000000000000;
        weights1[48739] <= 16'b0000000000001111;
        weights1[48740] <= 16'b1111111111110100;
        weights1[48741] <= 16'b1111111111111000;
        weights1[48742] <= 16'b1111111111100000;
        weights1[48743] <= 16'b0000000000000000;
        weights1[48744] <= 16'b1111111111101101;
        weights1[48745] <= 16'b1111111111110111;
        weights1[48746] <= 16'b1111111111111101;
        weights1[48747] <= 16'b0000000000000000;
        weights1[48748] <= 16'b1111111111111111;
        weights1[48749] <= 16'b1111111111110110;
        weights1[48750] <= 16'b1111111111111110;
        weights1[48751] <= 16'b1111111111111001;
        weights1[48752] <= 16'b1111111111110111;
        weights1[48753] <= 16'b0000000000001101;
        weights1[48754] <= 16'b1111111111110000;
        weights1[48755] <= 16'b0000000000001010;
        weights1[48756] <= 16'b0000000000001101;
        weights1[48757] <= 16'b1111111111111011;
        weights1[48758] <= 16'b1111111111110100;
        weights1[48759] <= 16'b0000000000000111;
        weights1[48760] <= 16'b1111111111110110;
        weights1[48761] <= 16'b0000000000000100;
        weights1[48762] <= 16'b1111111111110011;
        weights1[48763] <= 16'b0000000000000010;
        weights1[48764] <= 16'b1111111111111110;
        weights1[48765] <= 16'b1111111111111000;
        weights1[48766] <= 16'b1111111111110100;
        weights1[48767] <= 16'b0000000000000000;
        weights1[48768] <= 16'b1111111111110110;
        weights1[48769] <= 16'b1111111111111010;
        weights1[48770] <= 16'b1111111111110100;
        weights1[48771] <= 16'b1111111111111100;
        weights1[48772] <= 16'b1111111111110101;
        weights1[48773] <= 16'b0000000000001100;
        weights1[48774] <= 16'b1111111111110100;
        weights1[48775] <= 16'b1111111111110001;
        weights1[48776] <= 16'b0000000000000011;
        weights1[48777] <= 16'b0000000000000011;
        weights1[48778] <= 16'b1111111111111100;
        weights1[48779] <= 16'b0000000000001101;
        weights1[48780] <= 16'b1111111111111100;
        weights1[48781] <= 16'b0000000000001110;
        weights1[48782] <= 16'b0000000000000010;
        weights1[48783] <= 16'b1111111111111101;
        weights1[48784] <= 16'b1111111111111110;
        weights1[48785] <= 16'b0000000000000001;
        weights1[48786] <= 16'b1111111111111001;
        weights1[48787] <= 16'b0000000000000011;
        weights1[48788] <= 16'b1111111111111001;
        weights1[48789] <= 16'b1111111111111011;
        weights1[48790] <= 16'b1111111111110010;
        weights1[48791] <= 16'b1111111111110111;
        weights1[48792] <= 16'b0000000000000101;
        weights1[48793] <= 16'b1111111111111010;
        weights1[48794] <= 16'b0000000000000100;
        weights1[48795] <= 16'b1111111111110110;
        weights1[48796] <= 16'b1111111111110000;
        weights1[48797] <= 16'b1111111111111101;
        weights1[48798] <= 16'b1111111111110110;
        weights1[48799] <= 16'b1111111111110101;
        weights1[48800] <= 16'b1111111111011100;
        weights1[48801] <= 16'b1111111111110000;
        weights1[48802] <= 16'b1111111111111100;
        weights1[48803] <= 16'b1111111111110011;
        weights1[48804] <= 16'b1111111111111111;
        weights1[48805] <= 16'b0000000000000001;
        weights1[48806] <= 16'b0000000000010000;
        weights1[48807] <= 16'b0000000000000001;
        weights1[48808] <= 16'b1111111111111010;
        weights1[48809] <= 16'b1111111111101110;
        weights1[48810] <= 16'b1111111111100111;
        weights1[48811] <= 16'b0000000000000110;
        weights1[48812] <= 16'b1111111111111111;
        weights1[48813] <= 16'b1111111111111001;
        weights1[48814] <= 16'b1111111111111001;
        weights1[48815] <= 16'b0000000000000101;
        weights1[48816] <= 16'b0000000000000001;
        weights1[48817] <= 16'b0000000000000011;
        weights1[48818] <= 16'b1111111111111111;
        weights1[48819] <= 16'b1111111111110010;
        weights1[48820] <= 16'b0000000000001011;
        weights1[48821] <= 16'b1111111111101111;
        weights1[48822] <= 16'b1111111111110100;
        weights1[48823] <= 16'b1111111111111010;
        weights1[48824] <= 16'b1111111111110110;
        weights1[48825] <= 16'b1111111111111101;
        weights1[48826] <= 16'b1111111111101010;
        weights1[48827] <= 16'b1111111111011111;
        weights1[48828] <= 16'b0000000000011110;
        weights1[48829] <= 16'b1111111111111110;
        weights1[48830] <= 16'b1111111111101010;
        weights1[48831] <= 16'b1111111111101110;
        weights1[48832] <= 16'b1111111111111000;
        weights1[48833] <= 16'b1111111111111110;
        weights1[48834] <= 16'b0000000000000010;
        weights1[48835] <= 16'b1111111111111100;
        weights1[48836] <= 16'b1111111111111000;
        weights1[48837] <= 16'b1111111111111011;
        weights1[48838] <= 16'b0000000000000111;
        weights1[48839] <= 16'b1111111111111000;
        weights1[48840] <= 16'b0000000000001001;
        weights1[48841] <= 16'b0000000000000110;
        weights1[48842] <= 16'b1111111111111110;
        weights1[48843] <= 16'b1111111111110111;
        weights1[48844] <= 16'b1111111111111101;
        weights1[48845] <= 16'b1111111111101010;
        weights1[48846] <= 16'b0000000000000001;
        weights1[48847] <= 16'b1111111111110010;
        weights1[48848] <= 16'b1111111111110011;
        weights1[48849] <= 16'b1111111111111001;
        weights1[48850] <= 16'b1111111111101011;
        weights1[48851] <= 16'b1111111111110000;
        weights1[48852] <= 16'b1111111111101110;
        weights1[48853] <= 16'b1111111111111010;
        weights1[48854] <= 16'b1111111111110001;
        weights1[48855] <= 16'b1111111111111000;
        weights1[48856] <= 16'b1111111111100000;
        weights1[48857] <= 16'b1111111111111010;
        weights1[48858] <= 16'b1111111111110001;
        weights1[48859] <= 16'b1111111111101000;
        weights1[48860] <= 16'b1111111111111011;
        weights1[48861] <= 16'b1111111111111110;
        weights1[48862] <= 16'b0000000000001110;
        weights1[48863] <= 16'b0000000000000010;
        weights1[48864] <= 16'b0000000000000011;
        weights1[48865] <= 16'b1111111111111010;
        weights1[48866] <= 16'b1111111111110101;
        weights1[48867] <= 16'b1111111111111101;
        weights1[48868] <= 16'b1111111111111000;
        weights1[48869] <= 16'b1111111111111100;
        weights1[48870] <= 16'b0000000000000010;
        weights1[48871] <= 16'b0000000000001010;
        weights1[48872] <= 16'b1111111111111100;
        weights1[48873] <= 16'b1111111111111001;
        weights1[48874] <= 16'b0000000000001010;
        weights1[48875] <= 16'b1111111111111110;
        weights1[48876] <= 16'b1111111111111111;
        weights1[48877] <= 16'b1111111111111010;
        weights1[48878] <= 16'b0000000000000001;
        weights1[48879] <= 16'b1111111111110111;
        weights1[48880] <= 16'b0000000000001110;
        weights1[48881] <= 16'b1111111111101111;
        weights1[48882] <= 16'b1111111111111100;
        weights1[48883] <= 16'b1111111111100101;
        weights1[48884] <= 16'b1111111111101011;
        weights1[48885] <= 16'b1111111111011011;
        weights1[48886] <= 16'b1111111111011101;
        weights1[48887] <= 16'b1111111111100001;
        weights1[48888] <= 16'b1111111111111110;
        weights1[48889] <= 16'b1111111111111000;
        weights1[48890] <= 16'b1111111111110100;
        weights1[48891] <= 16'b0000000000001011;
        weights1[48892] <= 16'b0000000000000111;
        weights1[48893] <= 16'b0000000000000010;
        weights1[48894] <= 16'b0000000000001000;
        weights1[48895] <= 16'b1111111111110000;
        weights1[48896] <= 16'b0000000000010110;
        weights1[48897] <= 16'b0000000000000010;
        weights1[48898] <= 16'b0000000000001000;
        weights1[48899] <= 16'b0000000000000010;
        weights1[48900] <= 16'b0000000000000010;
        weights1[48901] <= 16'b1111111111111100;
        weights1[48902] <= 16'b0000000000000011;
        weights1[48903] <= 16'b0000000000001001;
        weights1[48904] <= 16'b1111111111111101;
        weights1[48905] <= 16'b0000000000000111;
        weights1[48906] <= 16'b0000000000000100;
        weights1[48907] <= 16'b1111111111111111;
        weights1[48908] <= 16'b1111111111110101;
        weights1[48909] <= 16'b0000000000000111;
        weights1[48910] <= 16'b1111111111111000;
        weights1[48911] <= 16'b0000000000010000;
        weights1[48912] <= 16'b1111111111111111;
        weights1[48913] <= 16'b1111111111101000;
        weights1[48914] <= 16'b1111111111110101;
        weights1[48915] <= 16'b1111111111110000;
        weights1[48916] <= 16'b1111111111111100;
        weights1[48917] <= 16'b1111111111111001;
        weights1[48918] <= 16'b0000000000000110;
        weights1[48919] <= 16'b1111111111111000;
        weights1[48920] <= 16'b1111111111101010;
        weights1[48921] <= 16'b1111111111111000;
        weights1[48922] <= 16'b1111111111111110;
        weights1[48923] <= 16'b1111111111110111;
        weights1[48924] <= 16'b1111111111111001;
        weights1[48925] <= 16'b1111111111110010;
        weights1[48926] <= 16'b1111111111110101;
        weights1[48927] <= 16'b1111111111111101;
        weights1[48928] <= 16'b1111111111110110;
        weights1[48929] <= 16'b1111111111110110;
        weights1[48930] <= 16'b1111111111111011;
        weights1[48931] <= 16'b1111111111111001;
        weights1[48932] <= 16'b1111111111111100;
        weights1[48933] <= 16'b1111111111110011;
        weights1[48934] <= 16'b1111111111111101;
        weights1[48935] <= 16'b0000000000000000;
        weights1[48936] <= 16'b1111111111111011;
        weights1[48937] <= 16'b1111111111111001;
        weights1[48938] <= 16'b1111111111110001;
        weights1[48939] <= 16'b1111111111111111;
        weights1[48940] <= 16'b1111111111100010;
        weights1[48941] <= 16'b1111111111110010;
        weights1[48942] <= 16'b1111111111011010;
        weights1[48943] <= 16'b0000000000000000;
        weights1[48944] <= 16'b1111111111110101;
        weights1[48945] <= 16'b0000000000000100;
        weights1[48946] <= 16'b1111111111110111;
        weights1[48947] <= 16'b0000000000001000;
        weights1[48948] <= 16'b1111111111101100;
        weights1[48949] <= 16'b1111111111110101;
        weights1[48950] <= 16'b0000000000000010;
        weights1[48951] <= 16'b0000000000010010;
        weights1[48952] <= 16'b0000000000000011;
        weights1[48953] <= 16'b1111111111110111;
        weights1[48954] <= 16'b1111111111111100;
        weights1[48955] <= 16'b0000000000000110;
        weights1[48956] <= 16'b1111111111111010;
        weights1[48957] <= 16'b1111111111111110;
        weights1[48958] <= 16'b0000000000000010;
        weights1[48959] <= 16'b0000000000000010;
        weights1[48960] <= 16'b0000000000001000;
        weights1[48961] <= 16'b1111111111111011;
        weights1[48962] <= 16'b0000000000000010;
        weights1[48963] <= 16'b1111111111110101;
        weights1[48964] <= 16'b0000000000001100;
        weights1[48965] <= 16'b1111111111111000;
        weights1[48966] <= 16'b0000000000000100;
        weights1[48967] <= 16'b1111111111110011;
        weights1[48968] <= 16'b0000000000001100;
        weights1[48969] <= 16'b1111111111111001;
        weights1[48970] <= 16'b0000000000001001;
        weights1[48971] <= 16'b0000000000001111;
        weights1[48972] <= 16'b0000000000000111;
        weights1[48973] <= 16'b0000000000001001;
        weights1[48974] <= 16'b0000000000000110;
        weights1[48975] <= 16'b1111111111111110;
        weights1[48976] <= 16'b1111111111111010;
        weights1[48977] <= 16'b0000000000001000;
        weights1[48978] <= 16'b0000000000010000;
        weights1[48979] <= 16'b1111111111111100;
        weights1[48980] <= 16'b1111111111111101;
        weights1[48981] <= 16'b1111111111101110;
        weights1[48982] <= 16'b1111111111110111;
        weights1[48983] <= 16'b0000000000000001;
        weights1[48984] <= 16'b0000000000000010;
        weights1[48985] <= 16'b0000000000000010;
        weights1[48986] <= 16'b1111111111111001;
        weights1[48987] <= 16'b1111111111110001;
        weights1[48988] <= 16'b1111111111111000;
        weights1[48989] <= 16'b1111111111111100;
        weights1[48990] <= 16'b1111111111110111;
        weights1[48991] <= 16'b1111111111111011;
        weights1[48992] <= 16'b1111111111111000;
        weights1[48993] <= 16'b0000000000000101;
        weights1[48994] <= 16'b0000000000000110;
        weights1[48995] <= 16'b0000000000010011;
        weights1[48996] <= 16'b0000000000001101;
        weights1[48997] <= 16'b0000000000011010;
        weights1[48998] <= 16'b0000000000001011;
        weights1[48999] <= 16'b0000000000001001;
        weights1[49000] <= 16'b0000000000001100;
        weights1[49001] <= 16'b1111111111111010;
        weights1[49002] <= 16'b1111111111110000;
        weights1[49003] <= 16'b0000000000000010;
        weights1[49004] <= 16'b1111111111110110;
        weights1[49005] <= 16'b1111111111111110;
        weights1[49006] <= 16'b1111111111110100;
        weights1[49007] <= 16'b1111111111111000;
        weights1[49008] <= 16'b1111111111110100;
        weights1[49009] <= 16'b1111111111110111;
        weights1[49010] <= 16'b1111111111111100;
        weights1[49011] <= 16'b1111111111111101;
        weights1[49012] <= 16'b1111111111101110;
        weights1[49013] <= 16'b1111111111110111;
        weights1[49014] <= 16'b0000000000000100;
        weights1[49015] <= 16'b1111111111110101;
        weights1[49016] <= 16'b0000000000000000;
        weights1[49017] <= 16'b1111111111110111;
        weights1[49018] <= 16'b0000000000000101;
        weights1[49019] <= 16'b1111111111111111;
        weights1[49020] <= 16'b0000000000000010;
        weights1[49021] <= 16'b1111111111111101;
        weights1[49022] <= 16'b0000000000010010;
        weights1[49023] <= 16'b0000000000000110;
        weights1[49024] <= 16'b0000000000001111;
        weights1[49025] <= 16'b0000000000001010;
        weights1[49026] <= 16'b0000000000101011;
        weights1[49027] <= 16'b0000000000001111;
        weights1[49028] <= 16'b0000000000011001;
        weights1[49029] <= 16'b0000000000001011;
        weights1[49030] <= 16'b1111111111111100;
        weights1[49031] <= 16'b1111111111110111;
        weights1[49032] <= 16'b1111111111100101;
        weights1[49033] <= 16'b1111111111101011;
        weights1[49034] <= 16'b0000000000000001;
        weights1[49035] <= 16'b1111111111110001;
        weights1[49036] <= 16'b1111111111111010;
        weights1[49037] <= 16'b1111111111110100;
        weights1[49038] <= 16'b0000000000000111;
        weights1[49039] <= 16'b1111111111110010;
        weights1[49040] <= 16'b1111111111110010;
        weights1[49041] <= 16'b1111111111111111;
        weights1[49042] <= 16'b1111111111101111;
        weights1[49043] <= 16'b1111111111110110;
        weights1[49044] <= 16'b1111111111110000;
        weights1[49045] <= 16'b1111111111110010;
        weights1[49046] <= 16'b1111111111110101;
        weights1[49047] <= 16'b0000000000010000;
        weights1[49048] <= 16'b0000000000010100;
        weights1[49049] <= 16'b0000000000001110;
        weights1[49050] <= 16'b0000000000011010;
        weights1[49051] <= 16'b0000000000000101;
        weights1[49052] <= 16'b0000000000011100;
        weights1[49053] <= 16'b0000000000101000;
        weights1[49054] <= 16'b0000000000011010;
        weights1[49055] <= 16'b0000000000001110;
        weights1[49056] <= 16'b0000000000010110;
        weights1[49057] <= 16'b0000000000010011;
        weights1[49058] <= 16'b0000000000000101;
        weights1[49059] <= 16'b0000000000000111;
        weights1[49060] <= 16'b0000000000001011;
        weights1[49061] <= 16'b1111111111110110;
        weights1[49062] <= 16'b1111111111110110;
        weights1[49063] <= 16'b0000000000000110;
        weights1[49064] <= 16'b1111111111111100;
        weights1[49065] <= 16'b0000000000000000;
        weights1[49066] <= 16'b1111111111111110;
        weights1[49067] <= 16'b1111111111110011;
        weights1[49068] <= 16'b1111111111110001;
        weights1[49069] <= 16'b0000000000000001;
        weights1[49070] <= 16'b1111111111111110;
        weights1[49071] <= 16'b0000000000000000;
        weights1[49072] <= 16'b0000000000000000;
        weights1[49073] <= 16'b0000000000000010;
        weights1[49074] <= 16'b0000000000001110;
        weights1[49075] <= 16'b0000000000010010;
        weights1[49076] <= 16'b0000000000001100;
        weights1[49077] <= 16'b0000000000100101;
        weights1[49078] <= 16'b0000000000010001;
        weights1[49079] <= 16'b0000000000001100;
        weights1[49080] <= 16'b0000000000011010;
        weights1[49081] <= 16'b0000000000011100;
        weights1[49082] <= 16'b0000000000011000;
        weights1[49083] <= 16'b0000000000000110;
        weights1[49084] <= 16'b0000000000011101;
        weights1[49085] <= 16'b0000000000010110;
        weights1[49086] <= 16'b0000000000010110;
        weights1[49087] <= 16'b0000000000001001;
        weights1[49088] <= 16'b0000000000100011;
        weights1[49089] <= 16'b0000000000001100;
        weights1[49090] <= 16'b1111111111111111;
        weights1[49091] <= 16'b1111111111110101;
        weights1[49092] <= 16'b1111111111111100;
        weights1[49093] <= 16'b1111111111110110;
        weights1[49094] <= 16'b0000000000000110;
        weights1[49095] <= 16'b0000000000001010;
        weights1[49096] <= 16'b0000000000000110;
        weights1[49097] <= 16'b0000000000001001;
        weights1[49098] <= 16'b0000000000000010;
        weights1[49099] <= 16'b0000000000001101;
        weights1[49100] <= 16'b0000000000010101;
        weights1[49101] <= 16'b0000000000100011;
        weights1[49102] <= 16'b0000000000011000;
        weights1[49103] <= 16'b0000000000000111;
        weights1[49104] <= 16'b0000000000011010;
        weights1[49105] <= 16'b0000000000001001;
        weights1[49106] <= 16'b0000000000001001;
        weights1[49107] <= 16'b1111111111111111;
        weights1[49108] <= 16'b0000000000000001;
        weights1[49109] <= 16'b0000000000011011;
        weights1[49110] <= 16'b0000000000001101;
        weights1[49111] <= 16'b0000000000001001;
        weights1[49112] <= 16'b0000000000010101;
        weights1[49113] <= 16'b0000000000011001;
        weights1[49114] <= 16'b0000000000100001;
        weights1[49115] <= 16'b0000000000101010;
        weights1[49116] <= 16'b0000000000010101;
        weights1[49117] <= 16'b0000000000011000;
        weights1[49118] <= 16'b0000000000011011;
        weights1[49119] <= 16'b0000000000001111;
        weights1[49120] <= 16'b0000000000010100;
        weights1[49121] <= 16'b0000000000010111;
        weights1[49122] <= 16'b0000000000010110;
        weights1[49123] <= 16'b0000000000010010;
        weights1[49124] <= 16'b0000000000011001;
        weights1[49125] <= 16'b0000000000011000;
        weights1[49126] <= 16'b0000000000101010;
        weights1[49127] <= 16'b0000000000011110;
        weights1[49128] <= 16'b0000000000101001;
        weights1[49129] <= 16'b0000000000010110;
        weights1[49130] <= 16'b0000000000001111;
        weights1[49131] <= 16'b0000000000011101;
        weights1[49132] <= 16'b0000000000001001;
        weights1[49133] <= 16'b0000000000000100;
        weights1[49134] <= 16'b0000000000010010;
        weights1[49135] <= 16'b1111111111111111;
        weights1[49136] <= 16'b0000000000011001;
        weights1[49137] <= 16'b0000000000010010;
        weights1[49138] <= 16'b0000000000001000;
        weights1[49139] <= 16'b1111111111110001;
        weights1[49140] <= 16'b0000000000010101;
        weights1[49141] <= 16'b0000000000001001;
        weights1[49142] <= 16'b0000000000011100;
        weights1[49143] <= 16'b0000000000010101;
        weights1[49144] <= 16'b0000000000111011;
        weights1[49145] <= 16'b0000000000010110;
        weights1[49146] <= 16'b0000000000101000;
        weights1[49147] <= 16'b0000000000100111;
        weights1[49148] <= 16'b0000000000011111;
        weights1[49149] <= 16'b0000000000011101;
        weights1[49150] <= 16'b0000000000100000;
        weights1[49151] <= 16'b0000000000011001;
        weights1[49152] <= 16'b0000000000011100;
        weights1[49153] <= 16'b0000000000100001;
        weights1[49154] <= 16'b0000000000010111;
        weights1[49155] <= 16'b0000000000010000;
        weights1[49156] <= 16'b0000000000010110;
        weights1[49157] <= 16'b0000000000011100;
        weights1[49158] <= 16'b0000000000101001;
        weights1[49159] <= 16'b0000000000010011;
        weights1[49160] <= 16'b0000000000011010;
        weights1[49161] <= 16'b0000000000001100;
        weights1[49162] <= 16'b0000000000100000;
        weights1[49163] <= 16'b1111111111110101;
        weights1[49164] <= 16'b0000000000000000;
        weights1[49165] <= 16'b1111111111101010;
        weights1[49166] <= 16'b1111111111101101;
        weights1[49167] <= 16'b1111111111010111;
        weights1[49168] <= 16'b0000000000011111;
        weights1[49169] <= 16'b0000000000001110;
        weights1[49170] <= 16'b0000000000001110;
        weights1[49171] <= 16'b0000000000010000;
        weights1[49172] <= 16'b0000000000011111;
        weights1[49173] <= 16'b0000000000010001;
        weights1[49174] <= 16'b0000000000010001;
        weights1[49175] <= 16'b0000000000011110;
        weights1[49176] <= 16'b0000000000011111;
        weights1[49177] <= 16'b0000000000001110;
        weights1[49178] <= 16'b0000000000011101;
        weights1[49179] <= 16'b0000000000010111;
        weights1[49180] <= 16'b0000000000010011;
        weights1[49181] <= 16'b0000000000011100;
        weights1[49182] <= 16'b0000000000011010;
        weights1[49183] <= 16'b1111111111111100;
        weights1[49184] <= 16'b0000000000101000;
        weights1[49185] <= 16'b0000000000000010;
        weights1[49186] <= 16'b0000000000011111;
        weights1[49187] <= 16'b0000000000001001;
        weights1[49188] <= 16'b0000000000001100;
        weights1[49189] <= 16'b0000000000011001;
        weights1[49190] <= 16'b0000000000001100;
        weights1[49191] <= 16'b1111111111110100;
        weights1[49192] <= 16'b1111111111100010;
        weights1[49193] <= 16'b1111111111000000;
        weights1[49194] <= 16'b1111111111000011;
        weights1[49195] <= 16'b1111111111001011;
        weights1[49196] <= 16'b0000000000000010;
        weights1[49197] <= 16'b0000000000001101;
        weights1[49198] <= 16'b1111111111111001;
        weights1[49199] <= 16'b1111111111111000;
        weights1[49200] <= 16'b0000000000001100;
        weights1[49201] <= 16'b0000000000010111;
        weights1[49202] <= 16'b1111111111111000;
        weights1[49203] <= 16'b0000000000001001;
        weights1[49204] <= 16'b0000000000000011;
        weights1[49205] <= 16'b0000000000010100;
        weights1[49206] <= 16'b0000000000000101;
        weights1[49207] <= 16'b0000000000001011;
        weights1[49208] <= 16'b0000000000001001;
        weights1[49209] <= 16'b1111111111110101;
        weights1[49210] <= 16'b0000000000001011;
        weights1[49211] <= 16'b0000000000000111;
        weights1[49212] <= 16'b0000000000010100;
        weights1[49213] <= 16'b1111111111111001;
        weights1[49214] <= 16'b1111111111101110;
        weights1[49215] <= 16'b0000000000011000;
        weights1[49216] <= 16'b1111111111110001;
        weights1[49217] <= 16'b1111111111110000;
        weights1[49218] <= 16'b1111111111100000;
        weights1[49219] <= 16'b1111111111000011;
        weights1[49220] <= 16'b1111111110110100;
        weights1[49221] <= 16'b1111111111000110;
        weights1[49222] <= 16'b1111111110111010;
        weights1[49223] <= 16'b1111111111010011;
        weights1[49224] <= 16'b1111111111101110;
        weights1[49225] <= 16'b1111111111101111;
        weights1[49226] <= 16'b1111111111100011;
        weights1[49227] <= 16'b1111111111011111;
        weights1[49228] <= 16'b0000000000000010;
        weights1[49229] <= 16'b1111111111111011;
        weights1[49230] <= 16'b0000000000000000;
        weights1[49231] <= 16'b0000000000000000;
        weights1[49232] <= 16'b1111111111111110;
        weights1[49233] <= 16'b1111111111110010;
        weights1[49234] <= 16'b0000000000001011;
        weights1[49235] <= 16'b1111111111111101;
        weights1[49236] <= 16'b0000000000001001;
        weights1[49237] <= 16'b1111111111111011;
        weights1[49238] <= 16'b0000000000001110;
        weights1[49239] <= 16'b1111111111110100;
        weights1[49240] <= 16'b1111111111100111;
        weights1[49241] <= 16'b1111111111001111;
        weights1[49242] <= 16'b1111111110111110;
        weights1[49243] <= 16'b1111111111000001;
        weights1[49244] <= 16'b1111111110110000;
        weights1[49245] <= 16'b1111111110011101;
        weights1[49246] <= 16'b1111111110011111;
        weights1[49247] <= 16'b1111111110100000;
        weights1[49248] <= 16'b1111111110011100;
        weights1[49249] <= 16'b1111111111000000;
        weights1[49250] <= 16'b1111111111001010;
        weights1[49251] <= 16'b1111111111011010;
        weights1[49252] <= 16'b1111111111101010;
        weights1[49253] <= 16'b1111111111100100;
        weights1[49254] <= 16'b1111111111010001;
        weights1[49255] <= 16'b1111111111010011;
        weights1[49256] <= 16'b1111111110111101;
        weights1[49257] <= 16'b1111111111001011;
        weights1[49258] <= 16'b1111111111011010;
        weights1[49259] <= 16'b1111111111010100;
        weights1[49260] <= 16'b1111111111000100;
        weights1[49261] <= 16'b1111111111001100;
        weights1[49262] <= 16'b1111111111101101;
        weights1[49263] <= 16'b1111111111001011;
        weights1[49264] <= 16'b1111111110110010;
        weights1[49265] <= 16'b1111111110100110;
        weights1[49266] <= 16'b1111111110011000;
        weights1[49267] <= 16'b1111111101111001;
        weights1[49268] <= 16'b1111111100100100;
        weights1[49269] <= 16'b1111111101000011;
        weights1[49270] <= 16'b1111111101101011;
        weights1[49271] <= 16'b1111111101110000;
        weights1[49272] <= 16'b1111111101111000;
        weights1[49273] <= 16'b1111111110011100;
        weights1[49274] <= 16'b1111111110100110;
        weights1[49275] <= 16'b1111111110111000;
        weights1[49276] <= 16'b1111111110101011;
        weights1[49277] <= 16'b1111111111001000;
        weights1[49278] <= 16'b1111111111010100;
        weights1[49279] <= 16'b1111111111100011;
        weights1[49280] <= 16'b1111111111110100;
        weights1[49281] <= 16'b1111111111101000;
        weights1[49282] <= 16'b1111111111011011;
        weights1[49283] <= 16'b1111111111001001;
        weights1[49284] <= 16'b1111111111001000;
        weights1[49285] <= 16'b1111111110110100;
        weights1[49286] <= 16'b1111111110110100;
        weights1[49287] <= 16'b1111111110100001;
        weights1[49288] <= 16'b1111111110010010;
        weights1[49289] <= 16'b1111111101110100;
        weights1[49290] <= 16'b1111111101011011;
        weights1[49291] <= 16'b1111111101011100;
        weights1[49292] <= 16'b1111111101110001;
        weights1[49293] <= 16'b1111111101110011;
        weights1[49294] <= 16'b1111111101100101;
        weights1[49295] <= 16'b1111111101110001;
        weights1[49296] <= 16'b1111111101111110;
        weights1[49297] <= 16'b1111111110011010;
        weights1[49298] <= 16'b1111111110100111;
        weights1[49299] <= 16'b1111111110101000;
        weights1[49300] <= 16'b1111111110001011;
        weights1[49301] <= 16'b1111111110101110;
        weights1[49302] <= 16'b1111111110110100;
        weights1[49303] <= 16'b1111111111000101;
        weights1[49304] <= 16'b1111111111001000;
        weights1[49305] <= 16'b1111111111011010;
        weights1[49306] <= 16'b1111111111100100;
        weights1[49307] <= 16'b1111111111101100;
        weights1[49308] <= 16'b1111111111110110;
        weights1[49309] <= 16'b1111111111110011;
        weights1[49310] <= 16'b1111111111101011;
        weights1[49311] <= 16'b1111111111011101;
        weights1[49312] <= 16'b1111111111010011;
        weights1[49313] <= 16'b1111111110111111;
        weights1[49314] <= 16'b1111111110111101;
        weights1[49315] <= 16'b1111111110110111;
        weights1[49316] <= 16'b1111111110110000;
        weights1[49317] <= 16'b1111111110011011;
        weights1[49318] <= 16'b1111111110110100;
        weights1[49319] <= 16'b1111111110111000;
        weights1[49320] <= 16'b1111111110101111;
        weights1[49321] <= 16'b1111111110110011;
        weights1[49322] <= 16'b1111111110111000;
        weights1[49323] <= 16'b1111111110101011;
        weights1[49324] <= 16'b1111111111000011;
        weights1[49325] <= 16'b1111111110111101;
        weights1[49326] <= 16'b1111111111000100;
        weights1[49327] <= 16'b1111111111001011;
        weights1[49328] <= 16'b1111111110111111;
        weights1[49329] <= 16'b1111111111010010;
        weights1[49330] <= 16'b1111111111011010;
        weights1[49331] <= 16'b1111111111010011;
        weights1[49332] <= 16'b1111111111011010;
        weights1[49333] <= 16'b1111111111101100;
        weights1[49334] <= 16'b1111111111101011;
        weights1[49335] <= 16'b1111111111111000;
        weights1[49336] <= 16'b1111111111111101;
        weights1[49337] <= 16'b0000000000000000;
        weights1[49338] <= 16'b1111111111111000;
        weights1[49339] <= 16'b1111111111110110;
        weights1[49340] <= 16'b1111111111100101;
        weights1[49341] <= 16'b1111111111011100;
        weights1[49342] <= 16'b1111111111011110;
        weights1[49343] <= 16'b1111111111001000;
        weights1[49344] <= 16'b1111111111001011;
        weights1[49345] <= 16'b1111111111010001;
        weights1[49346] <= 16'b1111111111011000;
        weights1[49347] <= 16'b1111111111000101;
        weights1[49348] <= 16'b1111111111001100;
        weights1[49349] <= 16'b1111111111010101;
        weights1[49350] <= 16'b1111111111010111;
        weights1[49351] <= 16'b1111111111010110;
        weights1[49352] <= 16'b1111111111011001;
        weights1[49353] <= 16'b1111111111010111;
        weights1[49354] <= 16'b1111111111001110;
        weights1[49355] <= 16'b1111111111011110;
        weights1[49356] <= 16'b1111111111011010;
        weights1[49357] <= 16'b1111111111100000;
        weights1[49358] <= 16'b1111111111101101;
        weights1[49359] <= 16'b1111111111101001;
        weights1[49360] <= 16'b1111111111101101;
        weights1[49361] <= 16'b1111111111110001;
        weights1[49362] <= 16'b1111111111111001;
        weights1[49363] <= 16'b1111111111111100;
        weights1[49364] <= 16'b1111111111111111;
        weights1[49365] <= 16'b1111111111111101;
        weights1[49366] <= 16'b1111111111111010;
        weights1[49367] <= 16'b1111111111111100;
        weights1[49368] <= 16'b1111111111110111;
        weights1[49369] <= 16'b1111111111110101;
        weights1[49370] <= 16'b1111111111101111;
        weights1[49371] <= 16'b1111111111101010;
        weights1[49372] <= 16'b1111111111101011;
        weights1[49373] <= 16'b1111111111100110;
        weights1[49374] <= 16'b1111111111100111;
        weights1[49375] <= 16'b1111111111101000;
        weights1[49376] <= 16'b1111111111101010;
        weights1[49377] <= 16'b1111111111101011;
        weights1[49378] <= 16'b1111111111100011;
        weights1[49379] <= 16'b1111111111101000;
        weights1[49380] <= 16'b1111111111100100;
        weights1[49381] <= 16'b1111111111100100;
        weights1[49382] <= 16'b1111111111011110;
        weights1[49383] <= 16'b1111111111100000;
        weights1[49384] <= 16'b1111111111110000;
        weights1[49385] <= 16'b1111111111100111;
        weights1[49386] <= 16'b1111111111110110;
        weights1[49387] <= 16'b1111111111110010;
        weights1[49388] <= 16'b1111111111110010;
        weights1[49389] <= 16'b1111111111110100;
        weights1[49390] <= 16'b1111111111111011;
        weights1[49391] <= 16'b1111111111111101;
        weights1[49392] <= 16'b0000000000000001;
        weights1[49393] <= 16'b0000000000000000;
        weights1[49394] <= 16'b0000000000000001;
        weights1[49395] <= 16'b0000000000000100;
        weights1[49396] <= 16'b0000000000000111;
        weights1[49397] <= 16'b0000000000001001;
        weights1[49398] <= 16'b0000000000010000;
        weights1[49399] <= 16'b0000000000011010;
        weights1[49400] <= 16'b0000000000011110;
        weights1[49401] <= 16'b0000000000100001;
        weights1[49402] <= 16'b0000000000110010;
        weights1[49403] <= 16'b0000000000111010;
        weights1[49404] <= 16'b0000000000101110;
        weights1[49405] <= 16'b0000000000110001;
        weights1[49406] <= 16'b0000000000001110;
        weights1[49407] <= 16'b0000000000100111;
        weights1[49408] <= 16'b0000000000110100;
        weights1[49409] <= 16'b0000000000101000;
        weights1[49410] <= 16'b0000000000101011;
        weights1[49411] <= 16'b0000000000100110;
        weights1[49412] <= 16'b0000000000010111;
        weights1[49413] <= 16'b0000000000100010;
        weights1[49414] <= 16'b0000000000010100;
        weights1[49415] <= 16'b0000000000001100;
        weights1[49416] <= 16'b0000000000001011;
        weights1[49417] <= 16'b0000000000000000;
        weights1[49418] <= 16'b0000000000001000;
        weights1[49419] <= 16'b0000000000000010;
        weights1[49420] <= 16'b0000000000000001;
        weights1[49421] <= 16'b1111111111111111;
        weights1[49422] <= 16'b0000000000000101;
        weights1[49423] <= 16'b0000000000000110;
        weights1[49424] <= 16'b0000000000001010;
        weights1[49425] <= 16'b0000000000001011;
        weights1[49426] <= 16'b0000000000010001;
        weights1[49427] <= 16'b0000000000001110;
        weights1[49428] <= 16'b0000000000010011;
        weights1[49429] <= 16'b0000000000001001;
        weights1[49430] <= 16'b0000000000001100;
        weights1[49431] <= 16'b0000000000010011;
        weights1[49432] <= 16'b0000000000000111;
        weights1[49433] <= 16'b1111111111101001;
        weights1[49434] <= 16'b0000000000000101;
        weights1[49435] <= 16'b0000000000010111;
        weights1[49436] <= 16'b0000000000010111;
        weights1[49437] <= 16'b0000000000000001;
        weights1[49438] <= 16'b0000000000010010;
        weights1[49439] <= 16'b0000000000010000;
        weights1[49440] <= 16'b0000000000010010;
        weights1[49441] <= 16'b0000000000001011;
        weights1[49442] <= 16'b0000000000010111;
        weights1[49443] <= 16'b0000000000001001;
        weights1[49444] <= 16'b0000000000001111;
        weights1[49445] <= 16'b0000000000000110;
        weights1[49446] <= 16'b0000000000001011;
        weights1[49447] <= 16'b0000000000000100;
        weights1[49448] <= 16'b0000000000000001;
        weights1[49449] <= 16'b0000000000000011;
        weights1[49450] <= 16'b0000000000001010;
        weights1[49451] <= 16'b0000000000000010;
        weights1[49452] <= 16'b0000000000001010;
        weights1[49453] <= 16'b0000000000001010;
        weights1[49454] <= 16'b0000000000001001;
        weights1[49455] <= 16'b0000000000001011;
        weights1[49456] <= 16'b0000000000000000;
        weights1[49457] <= 16'b0000000000000001;
        weights1[49458] <= 16'b0000000000000101;
        weights1[49459] <= 16'b0000000000010000;
        weights1[49460] <= 16'b1111111111111011;
        weights1[49461] <= 16'b1111111111101111;
        weights1[49462] <= 16'b1111111111111001;
        weights1[49463] <= 16'b1111111111110110;
        weights1[49464] <= 16'b0000000000000000;
        weights1[49465] <= 16'b1111111111110110;
        weights1[49466] <= 16'b0000000000000101;
        weights1[49467] <= 16'b1111111111110100;
        weights1[49468] <= 16'b1111111111111101;
        weights1[49469] <= 16'b0000000000001001;
        weights1[49470] <= 16'b0000000000010101;
        weights1[49471] <= 16'b0000000000001010;
        weights1[49472] <= 16'b0000000000001011;
        weights1[49473] <= 16'b0000000000010011;
        weights1[49474] <= 16'b0000000000010001;
        weights1[49475] <= 16'b0000000000001000;
        weights1[49476] <= 16'b0000000000000010;
        weights1[49477] <= 16'b0000000000000001;
        weights1[49478] <= 16'b1111111111111110;
        weights1[49479] <= 16'b0000000000001101;
        weights1[49480] <= 16'b0000000000000110;
        weights1[49481] <= 16'b0000000000000110;
        weights1[49482] <= 16'b0000000000000000;
        weights1[49483] <= 16'b1111111111111100;
        weights1[49484] <= 16'b1111111111101101;
        weights1[49485] <= 16'b1111111111111000;
        weights1[49486] <= 16'b1111111111111001;
        weights1[49487] <= 16'b1111111111111011;
        weights1[49488] <= 16'b1111111111101101;
        weights1[49489] <= 16'b1111111111111101;
        weights1[49490] <= 16'b0000000000000011;
        weights1[49491] <= 16'b1111111111110001;
        weights1[49492] <= 16'b1111111111100100;
        weights1[49493] <= 16'b1111111111111010;
        weights1[49494] <= 16'b1111111111111111;
        weights1[49495] <= 16'b1111111111101101;
        weights1[49496] <= 16'b1111111111100110;
        weights1[49497] <= 16'b1111111111110011;
        weights1[49498] <= 16'b1111111111111000;
        weights1[49499] <= 16'b1111111111110110;
        weights1[49500] <= 16'b1111111111111101;
        weights1[49501] <= 16'b0000000000001111;
        weights1[49502] <= 16'b0000000000001010;
        weights1[49503] <= 16'b0000000000001001;
        weights1[49504] <= 16'b0000000000000000;
        weights1[49505] <= 16'b0000000000000011;
        weights1[49506] <= 16'b1111111111111110;
        weights1[49507] <= 16'b0000000000000011;
        weights1[49508] <= 16'b0000000000001100;
        weights1[49509] <= 16'b0000000000000011;
        weights1[49510] <= 16'b0000000000000011;
        weights1[49511] <= 16'b1111111111111010;
        weights1[49512] <= 16'b0000000000001100;
        weights1[49513] <= 16'b0000000000000101;
        weights1[49514] <= 16'b1111111111101101;
        weights1[49515] <= 16'b1111111111101101;
        weights1[49516] <= 16'b1111111111100010;
        weights1[49517] <= 16'b1111111111111101;
        weights1[49518] <= 16'b1111111111111000;
        weights1[49519] <= 16'b1111111111111101;
        weights1[49520] <= 16'b1111111111101000;
        weights1[49521] <= 16'b0000000000000000;
        weights1[49522] <= 16'b1111111111111110;
        weights1[49523] <= 16'b1111111111110011;
        weights1[49524] <= 16'b1111111111101100;
        weights1[49525] <= 16'b1111111111111001;
        weights1[49526] <= 16'b1111111111110100;
        weights1[49527] <= 16'b1111111111100000;
        weights1[49528] <= 16'b0000000000000001;
        weights1[49529] <= 16'b0000000000000000;
        weights1[49530] <= 16'b0000000000000010;
        weights1[49531] <= 16'b0000000000000010;
        weights1[49532] <= 16'b1111111111111111;
        weights1[49533] <= 16'b0000000000000011;
        weights1[49534] <= 16'b1111111111111110;
        weights1[49535] <= 16'b0000000000000110;
        weights1[49536] <= 16'b0000000000011000;
        weights1[49537] <= 16'b0000000000011001;
        weights1[49538] <= 16'b0000000000000000;
        weights1[49539] <= 16'b1111111111111011;
        weights1[49540] <= 16'b0000000000011010;
        weights1[49541] <= 16'b1111111111101101;
        weights1[49542] <= 16'b0000000000001010;
        weights1[49543] <= 16'b1111111111101111;
        weights1[49544] <= 16'b1111111111110000;
        weights1[49545] <= 16'b0000000000001001;
        weights1[49546] <= 16'b1111111111111110;
        weights1[49547] <= 16'b0000000000010010;
        weights1[49548] <= 16'b0000000000010010;
        weights1[49549] <= 16'b0000000000011000;
        weights1[49550] <= 16'b1111111111100111;
        weights1[49551] <= 16'b1111111111100011;
        weights1[49552] <= 16'b1111111111110010;
        weights1[49553] <= 16'b1111111111100011;
        weights1[49554] <= 16'b1111111111110101;
        weights1[49555] <= 16'b1111111111110111;
        weights1[49556] <= 16'b0000000000001100;
        weights1[49557] <= 16'b0000000000000000;
        weights1[49558] <= 16'b0000000000000000;
        weights1[49559] <= 16'b0000000000000011;
        weights1[49560] <= 16'b1111111111111110;
        weights1[49561] <= 16'b1111111111111111;
        weights1[49562] <= 16'b1111111111110111;
        weights1[49563] <= 16'b0000000000000001;
        weights1[49564] <= 16'b0000000000001001;
        weights1[49565] <= 16'b0000000000010110;
        weights1[49566] <= 16'b0000000000000011;
        weights1[49567] <= 16'b0000000000010000;
        weights1[49568] <= 16'b0000000000001100;
        weights1[49569] <= 16'b0000000000000001;
        weights1[49570] <= 16'b0000000000000101;
        weights1[49571] <= 16'b0000000000000110;
        weights1[49572] <= 16'b1111111111101111;
        weights1[49573] <= 16'b0000000000001100;
        weights1[49574] <= 16'b1111111111111001;
        weights1[49575] <= 16'b1111111111110010;
        weights1[49576] <= 16'b0000000000001010;
        weights1[49577] <= 16'b1111111111111110;
        weights1[49578] <= 16'b0000000000010101;
        weights1[49579] <= 16'b0000000000000001;
        weights1[49580] <= 16'b1111111111111001;
        weights1[49581] <= 16'b0000000000000100;
        weights1[49582] <= 16'b0000000000000110;
        weights1[49583] <= 16'b1111111111011011;
        weights1[49584] <= 16'b0000000000001100;
        weights1[49585] <= 16'b0000000000000100;
        weights1[49586] <= 16'b0000000000001010;
        weights1[49587] <= 16'b0000000000000000;
        weights1[49588] <= 16'b1111111111111100;
        weights1[49589] <= 16'b1111111111111001;
        weights1[49590] <= 16'b1111111111110100;
        weights1[49591] <= 16'b0000000000001110;
        weights1[49592] <= 16'b0000000000001010;
        weights1[49593] <= 16'b1111111111111101;
        weights1[49594] <= 16'b0000000000000011;
        weights1[49595] <= 16'b0000000000011111;
        weights1[49596] <= 16'b1111111111111110;
        weights1[49597] <= 16'b1111111111100101;
        weights1[49598] <= 16'b0000000000001111;
        weights1[49599] <= 16'b1111111111111000;
        weights1[49600] <= 16'b0000000000001111;
        weights1[49601] <= 16'b0000000000010111;
        weights1[49602] <= 16'b0000000000000110;
        weights1[49603] <= 16'b0000000000001011;
        weights1[49604] <= 16'b0000000000000011;
        weights1[49605] <= 16'b1111111111110111;
        weights1[49606] <= 16'b1111111111101110;
        weights1[49607] <= 16'b1111111111111011;
        weights1[49608] <= 16'b0000000000000100;
        weights1[49609] <= 16'b0000000000001011;
        weights1[49610] <= 16'b0000000000001011;
        weights1[49611] <= 16'b0000000000001011;
        weights1[49612] <= 16'b0000000000001111;
        weights1[49613] <= 16'b0000000000010001;
        weights1[49614] <= 16'b0000000000000011;
        weights1[49615] <= 16'b1111111111111100;
        weights1[49616] <= 16'b0000000000000100;
        weights1[49617] <= 16'b1111111111111000;
        weights1[49618] <= 16'b0000000000001010;
        weights1[49619] <= 16'b0000000000000010;
        weights1[49620] <= 16'b0000000000001111;
        weights1[49621] <= 16'b0000000000010101;
        weights1[49622] <= 16'b0000000000010111;
        weights1[49623] <= 16'b0000000000011111;
        weights1[49624] <= 16'b0000000000011101;
        weights1[49625] <= 16'b0000000000000010;
        weights1[49626] <= 16'b0000000000011000;
        weights1[49627] <= 16'b0000000000001110;
        weights1[49628] <= 16'b1111111111100111;
        weights1[49629] <= 16'b1111111111110100;
        weights1[49630] <= 16'b1111111111110111;
        weights1[49631] <= 16'b0000000000011110;
        weights1[49632] <= 16'b0000000000000000;
        weights1[49633] <= 16'b0000000000001001;
        weights1[49634] <= 16'b1111111111111100;
        weights1[49635] <= 16'b0000000000000001;
        weights1[49636] <= 16'b0000000000010111;
        weights1[49637] <= 16'b0000000000010100;
        weights1[49638] <= 16'b0000000000010010;
        weights1[49639] <= 16'b0000000000001101;
        weights1[49640] <= 16'b0000000000001110;
        weights1[49641] <= 16'b0000000000001110;
        weights1[49642] <= 16'b1111111111111111;
        weights1[49643] <= 16'b0000000000000010;
        weights1[49644] <= 16'b1111111111111110;
        weights1[49645] <= 16'b0000000000001000;
        weights1[49646] <= 16'b0000000000000010;
        weights1[49647] <= 16'b0000000000000000;
        weights1[49648] <= 16'b0000000000010111;
        weights1[49649] <= 16'b0000000000000110;
        weights1[49650] <= 16'b1111111111111111;
        weights1[49651] <= 16'b0000000000011101;
        weights1[49652] <= 16'b0000000000101001;
        weights1[49653] <= 16'b0000000000001100;
        weights1[49654] <= 16'b0000000000001011;
        weights1[49655] <= 16'b0000000000010111;
        weights1[49656] <= 16'b0000000000000000;
        weights1[49657] <= 16'b0000000000000110;
        weights1[49658] <= 16'b0000000000010111;
        weights1[49659] <= 16'b1111111111101011;
        weights1[49660] <= 16'b0000000000001111;
        weights1[49661] <= 16'b0000000000001000;
        weights1[49662] <= 16'b0000000000010001;
        weights1[49663] <= 16'b0000000000000100;
        weights1[49664] <= 16'b0000000000011000;
        weights1[49665] <= 16'b0000000000000100;
        weights1[49666] <= 16'b1111111111111010;
        weights1[49667] <= 16'b0000000000001100;
        weights1[49668] <= 16'b0000000000010011;
        weights1[49669] <= 16'b0000000000001100;
        weights1[49670] <= 16'b0000000000011000;
        weights1[49671] <= 16'b0000000000010001;
        weights1[49672] <= 16'b1111111111111111;
        weights1[49673] <= 16'b0000000000001001;
        weights1[49674] <= 16'b0000000000010101;
        weights1[49675] <= 16'b0000000000010011;
        weights1[49676] <= 16'b0000000000010110;
        weights1[49677] <= 16'b0000000000010001;
        weights1[49678] <= 16'b0000000000000101;
        weights1[49679] <= 16'b0000000000010001;
        weights1[49680] <= 16'b0000000000011110;
        weights1[49681] <= 16'b0000000000001111;
        weights1[49682] <= 16'b0000000000100100;
        weights1[49683] <= 16'b0000000000001011;
        weights1[49684] <= 16'b1111111111111001;
        weights1[49685] <= 16'b0000000000010111;
        weights1[49686] <= 16'b0000000000011001;
        weights1[49687] <= 16'b0000000000011101;
        weights1[49688] <= 16'b0000000000010111;
        weights1[49689] <= 16'b0000000000010001;
        weights1[49690] <= 16'b0000000000000000;
        weights1[49691] <= 16'b0000000000011011;
        weights1[49692] <= 16'b0000000000010111;
        weights1[49693] <= 16'b0000000000011011;
        weights1[49694] <= 16'b0000000000001110;
        weights1[49695] <= 16'b0000000000001101;
        weights1[49696] <= 16'b0000000000001010;
        weights1[49697] <= 16'b0000000000011111;
        weights1[49698] <= 16'b0000000000001101;
        weights1[49699] <= 16'b0000000000001010;
        weights1[49700] <= 16'b0000000000000000;
        weights1[49701] <= 16'b0000000000001100;
        weights1[49702] <= 16'b0000000000011100;
        weights1[49703] <= 16'b0000000000010011;
        weights1[49704] <= 16'b1111111111111101;
        weights1[49705] <= 16'b0000000000001010;
        weights1[49706] <= 16'b0000000000011100;
        weights1[49707] <= 16'b0000000000010110;
        weights1[49708] <= 16'b0000000000101010;
        weights1[49709] <= 16'b0000000000010011;
        weights1[49710] <= 16'b0000000000100100;
        weights1[49711] <= 16'b0000000000101110;
        weights1[49712] <= 16'b0000000000100111;
        weights1[49713] <= 16'b0000000000100001;
        weights1[49714] <= 16'b0000000000011110;
        weights1[49715] <= 16'b0000000000010101;
        weights1[49716] <= 16'b0000000000101001;
        weights1[49717] <= 16'b0000000000100110;
        weights1[49718] <= 16'b0000000000100010;
        weights1[49719] <= 16'b0000000000001110;
        weights1[49720] <= 16'b0000000000101011;
        weights1[49721] <= 16'b0000000000010101;
        weights1[49722] <= 16'b0000000000010101;
        weights1[49723] <= 16'b0000000000101011;
        weights1[49724] <= 16'b0000000000000110;
        weights1[49725] <= 16'b0000000000010110;
        weights1[49726] <= 16'b0000000000001110;
        weights1[49727] <= 16'b0000000000000110;
        weights1[49728] <= 16'b1111111111111111;
        weights1[49729] <= 16'b0000000000000110;
        weights1[49730] <= 16'b0000000000010111;
        weights1[49731] <= 16'b0000000000011010;
        weights1[49732] <= 16'b0000000000010111;
        weights1[49733] <= 16'b1111111111110100;
        weights1[49734] <= 16'b0000000000010011;
        weights1[49735] <= 16'b0000000000010101;
        weights1[49736] <= 16'b1111111111111001;
        weights1[49737] <= 16'b0000000000100101;
        weights1[49738] <= 16'b0000000000100010;
        weights1[49739] <= 16'b0000000000100011;
        weights1[49740] <= 16'b0000000000100110;
        weights1[49741] <= 16'b0000000000011101;
        weights1[49742] <= 16'b0000000000011010;
        weights1[49743] <= 16'b0000000000011100;
        weights1[49744] <= 16'b0000000000100101;
        weights1[49745] <= 16'b0000000000011101;
        weights1[49746] <= 16'b0000000000100001;
        weights1[49747] <= 16'b0000000000101000;
        weights1[49748] <= 16'b0000000000011001;
        weights1[49749] <= 16'b0000000000101100;
        weights1[49750] <= 16'b0000000000001001;
        weights1[49751] <= 16'b0000000000101010;
        weights1[49752] <= 16'b0000000000100100;
        weights1[49753] <= 16'b0000000000100100;
        weights1[49754] <= 16'b0000000000010010;
        weights1[49755] <= 16'b0000000000001110;
        weights1[49756] <= 16'b1111111111111110;
        weights1[49757] <= 16'b0000000000001000;
        weights1[49758] <= 16'b0000000000010010;
        weights1[49759] <= 16'b0000000000100110;
        weights1[49760] <= 16'b0000000000011110;
        weights1[49761] <= 16'b0000000000001101;
        weights1[49762] <= 16'b0000000000001010;
        weights1[49763] <= 16'b0000000000001011;
        weights1[49764] <= 16'b0000000000001100;
        weights1[49765] <= 16'b0000000000001000;
        weights1[49766] <= 16'b0000000000011100;
        weights1[49767] <= 16'b0000000000100110;
        weights1[49768] <= 16'b0000000000110010;
        weights1[49769] <= 16'b0000000000100010;
        weights1[49770] <= 16'b0000000000011011;
        weights1[49771] <= 16'b0000000000010001;
        weights1[49772] <= 16'b0000000000100110;
        weights1[49773] <= 16'b0000000000101000;
        weights1[49774] <= 16'b0000000000001001;
        weights1[49775] <= 16'b0000000000101000;
        weights1[49776] <= 16'b0000000000100000;
        weights1[49777] <= 16'b0000000000010010;
        weights1[49778] <= 16'b0000000000011110;
        weights1[49779] <= 16'b0000000000100000;
        weights1[49780] <= 16'b0000000000100110;
        weights1[49781] <= 16'b0000000000010001;
        weights1[49782] <= 16'b0000000000010001;
        weights1[49783] <= 16'b1111111111111111;
        weights1[49784] <= 16'b1111111111111011;
        weights1[49785] <= 16'b0000000000000000;
        weights1[49786] <= 16'b0000000000001010;
        weights1[49787] <= 16'b1111111111111010;
        weights1[49788] <= 16'b1111111111111000;
        weights1[49789] <= 16'b0000000000011001;
        weights1[49790] <= 16'b0000000000001000;
        weights1[49791] <= 16'b0000000000011011;
        weights1[49792] <= 16'b0000000000100011;
        weights1[49793] <= 16'b0000000000100000;
        weights1[49794] <= 16'b0000000000100110;
        weights1[49795] <= 16'b0000000000110011;
        weights1[49796] <= 16'b0000000000101100;
        weights1[49797] <= 16'b0000000000100001;
        weights1[49798] <= 16'b0000000000100101;
        weights1[49799] <= 16'b0000000000110010;
        weights1[49800] <= 16'b0000000000011010;
        weights1[49801] <= 16'b0000000000011111;
        weights1[49802] <= 16'b0000000000010010;
        weights1[49803] <= 16'b0000000000010000;
        weights1[49804] <= 16'b0000000000100001;
        weights1[49805] <= 16'b0000000000100110;
        weights1[49806] <= 16'b0000000000101110;
        weights1[49807] <= 16'b0000000000001111;
        weights1[49808] <= 16'b0000000000000111;
        weights1[49809] <= 16'b1111111111111011;
        weights1[49810] <= 16'b0000000000000101;
        weights1[49811] <= 16'b0000000000000110;
        weights1[49812] <= 16'b1111111111111110;
        weights1[49813] <= 16'b1111111111101111;
        weights1[49814] <= 16'b1111111111100110;
        weights1[49815] <= 16'b1111111111100010;
        weights1[49816] <= 16'b1111111111101110;
        weights1[49817] <= 16'b1111111111110001;
        weights1[49818] <= 16'b1111111111101001;
        weights1[49819] <= 16'b0000000000000010;
        weights1[49820] <= 16'b1111111111110110;
        weights1[49821] <= 16'b1111111111111101;
        weights1[49822] <= 16'b0000000000001000;
        weights1[49823] <= 16'b0000000000010111;
        weights1[49824] <= 16'b0000000000101100;
        weights1[49825] <= 16'b0000000000111000;
        weights1[49826] <= 16'b0000000000111110;
        weights1[49827] <= 16'b0000000000101110;
        weights1[49828] <= 16'b0000000000101110;
        weights1[49829] <= 16'b0000000000100110;
        weights1[49830] <= 16'b0000000000110011;
        weights1[49831] <= 16'b0000000000101000;
        weights1[49832] <= 16'b0000000000010100;
        weights1[49833] <= 16'b0000000000001100;
        weights1[49834] <= 16'b0000000000000010;
        weights1[49835] <= 16'b0000000000010010;
        weights1[49836] <= 16'b0000000000001001;
        weights1[49837] <= 16'b0000000000000001;
        weights1[49838] <= 16'b0000000000000100;
        weights1[49839] <= 16'b0000000000001100;
        weights1[49840] <= 16'b1111111111110001;
        weights1[49841] <= 16'b1111111111100100;
        weights1[49842] <= 16'b1111111111101011;
        weights1[49843] <= 16'b1111111111011000;
        weights1[49844] <= 16'b1111111111011111;
        weights1[49845] <= 16'b1111111111001010;
        weights1[49846] <= 16'b1111111111101110;
        weights1[49847] <= 16'b1111111111111001;
        weights1[49848] <= 16'b1111111111011100;
        weights1[49849] <= 16'b1111111111101000;
        weights1[49850] <= 16'b1111111111101100;
        weights1[49851] <= 16'b1111111111100010;
        weights1[49852] <= 16'b0000000000000111;
        weights1[49853] <= 16'b0000000000001000;
        weights1[49854] <= 16'b0000000000110010;
        weights1[49855] <= 16'b0000000000010001;
        weights1[49856] <= 16'b0000000000011111;
        weights1[49857] <= 16'b0000000000010000;
        weights1[49858] <= 16'b0000000000010110;
        weights1[49859] <= 16'b1111111111110000;
        weights1[49860] <= 16'b1111111111100110;
        weights1[49861] <= 16'b1111111111111101;
        weights1[49862] <= 16'b1111111111011000;
        weights1[49863] <= 16'b1111111111101011;
        weights1[49864] <= 16'b1111111111111100;
        weights1[49865] <= 16'b1111111111111000;
        weights1[49866] <= 16'b1111111111111011;
        weights1[49867] <= 16'b1111111111111101;
        weights1[49868] <= 16'b1111111111101100;
        weights1[49869] <= 16'b1111111111011111;
        weights1[49870] <= 16'b1111111111001110;
        weights1[49871] <= 16'b1111111111001101;
        weights1[49872] <= 16'b1111111111001101;
        weights1[49873] <= 16'b1111111111010101;
        weights1[49874] <= 16'b1111111111011111;
        weights1[49875] <= 16'b1111111111000110;
        weights1[49876] <= 16'b1111111110111011;
        weights1[49877] <= 16'b1111111110110010;
        weights1[49878] <= 16'b1111111110101110;
        weights1[49879] <= 16'b1111111110101000;
        weights1[49880] <= 16'b1111111110110000;
        weights1[49881] <= 16'b1111111110110111;
        weights1[49882] <= 16'b1111111111001111;
        weights1[49883] <= 16'b1111111111010011;
        weights1[49884] <= 16'b1111111111011010;
        weights1[49885] <= 16'b1111111111100011;
        weights1[49886] <= 16'b1111111111001110;
        weights1[49887] <= 16'b1111111111010101;
        weights1[49888] <= 16'b1111111111001101;
        weights1[49889] <= 16'b1111111111010110;
        weights1[49890] <= 16'b1111111111000110;
        weights1[49891] <= 16'b1111111111001100;
        weights1[49892] <= 16'b1111111111001011;
        weights1[49893] <= 16'b1111111111011110;
        weights1[49894] <= 16'b1111111111100111;
        weights1[49895] <= 16'b1111111111111011;
        weights1[49896] <= 16'b1111111111101111;
        weights1[49897] <= 16'b1111111111011111;
        weights1[49898] <= 16'b1111111111010110;
        weights1[49899] <= 16'b1111111111011110;
        weights1[49900] <= 16'b1111111111010101;
        weights1[49901] <= 16'b1111111111010000;
        weights1[49902] <= 16'b1111111111001001;
        weights1[49903] <= 16'b1111111111010001;
        weights1[49904] <= 16'b1111111111011100;
        weights1[49905] <= 16'b1111111111010101;
        weights1[49906] <= 16'b1111111111000010;
        weights1[49907] <= 16'b1111111110101111;
        weights1[49908] <= 16'b1111111110011001;
        weights1[49909] <= 16'b1111111110010111;
        weights1[49910] <= 16'b1111111101111000;
        weights1[49911] <= 16'b1111111110100011;
        weights1[49912] <= 16'b1111111110100100;
        weights1[49913] <= 16'b1111111110100111;
        weights1[49914] <= 16'b1111111111000011;
        weights1[49915] <= 16'b1111111111011000;
        weights1[49916] <= 16'b1111111110110101;
        weights1[49917] <= 16'b1111111111011010;
        weights1[49918] <= 16'b1111111110110010;
        weights1[49919] <= 16'b1111111110111011;
        weights1[49920] <= 16'b1111111110110010;
        weights1[49921] <= 16'b1111111111001111;
        weights1[49922] <= 16'b1111111111100101;
        weights1[49923] <= 16'b1111111111110000;
        weights1[49924] <= 16'b1111111111101111;
        weights1[49925] <= 16'b1111111111100110;
        weights1[49926] <= 16'b1111111111100011;
        weights1[49927] <= 16'b1111111111100110;
        weights1[49928] <= 16'b1111111111100101;
        weights1[49929] <= 16'b1111111111100101;
        weights1[49930] <= 16'b1111111111011101;
        weights1[49931] <= 16'b1111111111010100;
        weights1[49932] <= 16'b1111111111011001;
        weights1[49933] <= 16'b1111111111010111;
        weights1[49934] <= 16'b1111111111001000;
        weights1[49935] <= 16'b1111111111010001;
        weights1[49936] <= 16'b1111111110111011;
        weights1[49937] <= 16'b1111111110111111;
        weights1[49938] <= 16'b1111111111001101;
        weights1[49939] <= 16'b1111111110111000;
        weights1[49940] <= 16'b1111111111000011;
        weights1[49941] <= 16'b1111111110111011;
        weights1[49942] <= 16'b1111111111000100;
        weights1[49943] <= 16'b1111111111001000;
        weights1[49944] <= 16'b1111111111001010;
        weights1[49945] <= 16'b1111111111010000;
        weights1[49946] <= 16'b1111111110101110;
        weights1[49947] <= 16'b1111111111000011;
        weights1[49948] <= 16'b1111111111000001;
        weights1[49949] <= 16'b1111111111010011;
        weights1[49950] <= 16'b1111111111011100;
        weights1[49951] <= 16'b1111111111110010;
        weights1[49952] <= 16'b1111111111110111;
        weights1[49953] <= 16'b1111111111101011;
        weights1[49954] <= 16'b1111111111100110;
        weights1[49955] <= 16'b1111111111101110;
        weights1[49956] <= 16'b1111111111100101;
        weights1[49957] <= 16'b0000000000000000;
        weights1[49958] <= 16'b1111111111110011;
        weights1[49959] <= 16'b1111111111011110;
        weights1[49960] <= 16'b1111111111010110;
        weights1[49961] <= 16'b1111111111010100;
        weights1[49962] <= 16'b1111111111011110;
        weights1[49963] <= 16'b1111111110111011;
        weights1[49964] <= 16'b1111111111000110;
        weights1[49965] <= 16'b1111111110111000;
        weights1[49966] <= 16'b1111111111001101;
        weights1[49967] <= 16'b1111111111000101;
        weights1[49968] <= 16'b1111111111010010;
        weights1[49969] <= 16'b1111111111000111;
        weights1[49970] <= 16'b1111111111010001;
        weights1[49971] <= 16'b1111111111010001;
        weights1[49972] <= 16'b1111111110111001;
        weights1[49973] <= 16'b1111111111001010;
        weights1[49974] <= 16'b1111111111001000;
        weights1[49975] <= 16'b1111111111010000;
        weights1[49976] <= 16'b1111111111010111;
        weights1[49977] <= 16'b1111111111011011;
        weights1[49978] <= 16'b1111111111100111;
        weights1[49979] <= 16'b1111111111111000;
        weights1[49980] <= 16'b1111111111111000;
        weights1[49981] <= 16'b1111111111111101;
        weights1[49982] <= 16'b1111111111110011;
        weights1[49983] <= 16'b1111111111111010;
        weights1[49984] <= 16'b1111111111111011;
        weights1[49985] <= 16'b1111111111101011;
        weights1[49986] <= 16'b1111111111101101;
        weights1[49987] <= 16'b1111111111010110;
        weights1[49988] <= 16'b1111111111011001;
        weights1[49989] <= 16'b1111111111011110;
        weights1[49990] <= 16'b1111111111110000;
        weights1[49991] <= 16'b1111111111010000;
        weights1[49992] <= 16'b1111111111000001;
        weights1[49993] <= 16'b1111111111000001;
        weights1[49994] <= 16'b1111111111001111;
        weights1[49995] <= 16'b1111111111001110;
        weights1[49996] <= 16'b1111111110111100;
        weights1[49997] <= 16'b1111111111000010;
        weights1[49998] <= 16'b1111111111001111;
        weights1[49999] <= 16'b1111111111010110;
        weights1[50000] <= 16'b1111111111001110;
        weights1[50001] <= 16'b1111111111011100;
        weights1[50002] <= 16'b1111111111011001;
        weights1[50003] <= 16'b1111111111011100;
        weights1[50004] <= 16'b1111111111100010;
        weights1[50005] <= 16'b1111111111011110;
        weights1[50006] <= 16'b1111111111101011;
        weights1[50007] <= 16'b1111111111110110;
        weights1[50008] <= 16'b1111111111111011;
        weights1[50009] <= 16'b1111111111111110;
        weights1[50010] <= 16'b1111111111110101;
        weights1[50011] <= 16'b1111111111111011;
        weights1[50012] <= 16'b1111111111110101;
        weights1[50013] <= 16'b1111111111110000;
        weights1[50014] <= 16'b1111111111101000;
        weights1[50015] <= 16'b1111111111100001;
        weights1[50016] <= 16'b1111111111111010;
        weights1[50017] <= 16'b1111111111011101;
        weights1[50018] <= 16'b1111111111101001;
        weights1[50019] <= 16'b1111111111100010;
        weights1[50020] <= 16'b1111111111000110;
        weights1[50021] <= 16'b1111111111101010;
        weights1[50022] <= 16'b1111111111011111;
        weights1[50023] <= 16'b1111111111011101;
        weights1[50024] <= 16'b1111111111011100;
        weights1[50025] <= 16'b1111111111010010;
        weights1[50026] <= 16'b1111111111100011;
        weights1[50027] <= 16'b1111111111010111;
        weights1[50028] <= 16'b1111111111100001;
        weights1[50029] <= 16'b1111111111110100;
        weights1[50030] <= 16'b1111111111101010;
        weights1[50031] <= 16'b1111111111010101;
        weights1[50032] <= 16'b1111111111101010;
        weights1[50033] <= 16'b1111111111101000;
        weights1[50034] <= 16'b1111111111110010;
        weights1[50035] <= 16'b1111111111110111;
        weights1[50036] <= 16'b1111111111111111;
        weights1[50037] <= 16'b1111111111111110;
        weights1[50038] <= 16'b1111111111110110;
        weights1[50039] <= 16'b1111111111111001;
        weights1[50040] <= 16'b1111111111101110;
        weights1[50041] <= 16'b1111111111100011;
        weights1[50042] <= 16'b1111111111110111;
        weights1[50043] <= 16'b1111111111011011;
        weights1[50044] <= 16'b1111111111011101;
        weights1[50045] <= 16'b1111111111101100;
        weights1[50046] <= 16'b1111111111101000;
        weights1[50047] <= 16'b1111111111101100;
        weights1[50048] <= 16'b0000000000001010;
        weights1[50049] <= 16'b1111111111110001;
        weights1[50050] <= 16'b1111111111011000;
        weights1[50051] <= 16'b1111111111010001;
        weights1[50052] <= 16'b0000000000000011;
        weights1[50053] <= 16'b1111111111101001;
        weights1[50054] <= 16'b1111111111011111;
        weights1[50055] <= 16'b1111111111111010;
        weights1[50056] <= 16'b1111111111011111;
        weights1[50057] <= 16'b1111111111101011;
        weights1[50058] <= 16'b1111111111101110;
        weights1[50059] <= 16'b1111111111101001;
        weights1[50060] <= 16'b1111111111101111;
        weights1[50061] <= 16'b1111111111110100;
        weights1[50062] <= 16'b1111111111110111;
        weights1[50063] <= 16'b1111111111111001;
        weights1[50064] <= 16'b1111111111111110;
        weights1[50065] <= 16'b1111111111111001;
        weights1[50066] <= 16'b1111111111110010;
        weights1[50067] <= 16'b1111111111110111;
        weights1[50068] <= 16'b1111111111110111;
        weights1[50069] <= 16'b1111111111100111;
        weights1[50070] <= 16'b1111111111101100;
        weights1[50071] <= 16'b1111111111001110;
        weights1[50072] <= 16'b1111111111010011;
        weights1[50073] <= 16'b1111111111100110;
        weights1[50074] <= 16'b1111111111101000;
        weights1[50075] <= 16'b1111111111110010;
        weights1[50076] <= 16'b1111111111111000;
        weights1[50077] <= 16'b1111111111101001;
        weights1[50078] <= 16'b1111111111100111;
        weights1[50079] <= 16'b1111111111011101;
        weights1[50080] <= 16'b1111111111101110;
        weights1[50081] <= 16'b1111111111011000;
        weights1[50082] <= 16'b1111111111101101;
        weights1[50083] <= 16'b1111111111100001;
        weights1[50084] <= 16'b0000000000000111;
        weights1[50085] <= 16'b1111111111110110;
        weights1[50086] <= 16'b1111111111110001;
        weights1[50087] <= 16'b1111111111101100;
        weights1[50088] <= 16'b1111111111110001;
        weights1[50089] <= 16'b1111111111111001;
        weights1[50090] <= 16'b0000000000000010;
        weights1[50091] <= 16'b1111111111111110;
        weights1[50092] <= 16'b1111111111111110;
        weights1[50093] <= 16'b1111111111111000;
        weights1[50094] <= 16'b1111111111111001;
        weights1[50095] <= 16'b1111111111110110;
        weights1[50096] <= 16'b1111111111111001;
        weights1[50097] <= 16'b1111111111101101;
        weights1[50098] <= 16'b1111111111010011;
        weights1[50099] <= 16'b1111111111001000;
        weights1[50100] <= 16'b1111111111010100;
        weights1[50101] <= 16'b1111111111100101;
        weights1[50102] <= 16'b1111111111001110;
        weights1[50103] <= 16'b1111111111000110;
        weights1[50104] <= 16'b1111111110011001;
        weights1[50105] <= 16'b1111111111001111;
        weights1[50106] <= 16'b1111111110111110;
        weights1[50107] <= 16'b1111111111100000;
        weights1[50108] <= 16'b1111111111000010;
        weights1[50109] <= 16'b1111111111000110;
        weights1[50110] <= 16'b1111111110101110;
        weights1[50111] <= 16'b1111111110101101;
        weights1[50112] <= 16'b1111111111001101;
        weights1[50113] <= 16'b1111111111010011;
        weights1[50114] <= 16'b1111111111101011;
        weights1[50115] <= 16'b1111111111110100;
        weights1[50116] <= 16'b1111111111110110;
        weights1[50117] <= 16'b1111111111111110;
        weights1[50118] <= 16'b0000000000000000;
        weights1[50119] <= 16'b0000000000000000;
        weights1[50120] <= 16'b1111111111111111;
        weights1[50121] <= 16'b1111111111111011;
        weights1[50122] <= 16'b1111111111111110;
        weights1[50123] <= 16'b1111111111111010;
        weights1[50124] <= 16'b1111111111111011;
        weights1[50125] <= 16'b1111111111111010;
        weights1[50126] <= 16'b1111111111110000;
        weights1[50127] <= 16'b1111111111100001;
        weights1[50128] <= 16'b1111111111001101;
        weights1[50129] <= 16'b1111111111001001;
        weights1[50130] <= 16'b1111111111010110;
        weights1[50131] <= 16'b1111111111001111;
        weights1[50132] <= 16'b1111111111010011;
        weights1[50133] <= 16'b1111111110111001;
        weights1[50134] <= 16'b1111111111001011;
        weights1[50135] <= 16'b1111111111010001;
        weights1[50136] <= 16'b1111111111000001;
        weights1[50137] <= 16'b1111111110111101;
        weights1[50138] <= 16'b1111111111001011;
        weights1[50139] <= 16'b1111111111000011;
        weights1[50140] <= 16'b1111111111010100;
        weights1[50141] <= 16'b1111111111011011;
        weights1[50142] <= 16'b1111111111100101;
        weights1[50143] <= 16'b1111111111110100;
        weights1[50144] <= 16'b1111111111111001;
        weights1[50145] <= 16'b1111111111111111;
        weights1[50146] <= 16'b0000000000000000;
        weights1[50147] <= 16'b0000000000000010;
        weights1[50148] <= 16'b0000000000000000;
        weights1[50149] <= 16'b1111111111111110;
        weights1[50150] <= 16'b0000000000000000;
        weights1[50151] <= 16'b0000000000000000;
        weights1[50152] <= 16'b1111111111111100;
        weights1[50153] <= 16'b1111111111111101;
        weights1[50154] <= 16'b1111111111111100;
        weights1[50155] <= 16'b1111111111110101;
        weights1[50156] <= 16'b1111111111101111;
        weights1[50157] <= 16'b1111111111100111;
        weights1[50158] <= 16'b1111111111100000;
        weights1[50159] <= 16'b1111111111101100;
        weights1[50160] <= 16'b1111111111110100;
        weights1[50161] <= 16'b1111111111101010;
        weights1[50162] <= 16'b1111111111011100;
        weights1[50163] <= 16'b1111111111100110;
        weights1[50164] <= 16'b1111111111011111;
        weights1[50165] <= 16'b1111111111011011;
        weights1[50166] <= 16'b1111111111010111;
        weights1[50167] <= 16'b1111111111100011;
        weights1[50168] <= 16'b1111111111100001;
        weights1[50169] <= 16'b1111111111100010;
        weights1[50170] <= 16'b1111111111110001;
        weights1[50171] <= 16'b1111111111110011;
        weights1[50172] <= 16'b1111111111111000;
        weights1[50173] <= 16'b1111111111111101;
        weights1[50174] <= 16'b1111111111111111;
        weights1[50175] <= 16'b0000000000000010;
        biases1[0] <= 16'b0000000001110011;
        biases1[1] <= 16'b0000000000100101;
        biases1[2] <= 16'b0000000001000000;
        biases1[3] <= 16'b0000000001010010;
        biases1[4] <= 16'b1111111111100000;
        biases1[5] <= 16'b0000000001000110;
        biases1[6] <= 16'b0000000000000000;
        biases1[7] <= 16'b0000000001010000;
        biases1[8] <= 16'b1111111101110101;
        biases1[9] <= 16'b1111111110010110;
        biases1[10] <= 16'b1111111111001111;
        biases1[11] <= 16'b0000000000011100;
        biases1[12] <= 16'b0000000001000100;
        biases1[13] <= 16'b0000000000011010;
        biases1[14] <= 16'b1111111111111001;
        biases1[15] <= 16'b1111111110010111;
        biases1[16] <= 16'b1111111110010011;
        biases1[17] <= 16'b0000000100011101;
        biases1[18] <= 16'b0000000000011001;
        biases1[19] <= 16'b1111111111111010;
        biases1[20] <= 16'b0000000001001100;
        biases1[21] <= 16'b0000000100001110;
        biases1[22] <= 16'b0000000001000101;
        biases1[23] <= 16'b1111111110100000;
        biases1[24] <= 16'b0000000001001101;
        biases1[25] <= 16'b0000000000011000;
        biases1[26] <= 16'b1111111111101101;
        biases1[27] <= 16'b0000000001001010;
        biases1[28] <= 16'b0000000010000110;
        biases1[29] <= 16'b0000000010011001;
        biases1[30] <= 16'b0000000000010111;
        biases1[31] <= 16'b0000000000100101;
        biases1[32] <= 16'b1111111111110100;
        biases1[33] <= 16'b1111111111101000;
        biases1[34] <= 16'b0000000010011111;
        biases1[35] <= 16'b0000000000110111;
        biases1[36] <= 16'b0000000000001001;
        biases1[37] <= 16'b0000000000101001;
        biases1[38] <= 16'b0000000000011000;
        biases1[39] <= 16'b0000000010011101;
        biases1[40] <= 16'b1111111001101000;
        biases1[41] <= 16'b1111111101011000;
        biases1[42] <= 16'b0000000010010111;
        biases1[43] <= 16'b0000000000000001;
        biases1[44] <= 16'b0000000000011001;
        biases1[45] <= 16'b1111111110001111;
        biases1[46] <= 16'b0000000001000110;
        biases1[47] <= 16'b0000000000101110;
        biases1[48] <= 16'b0000000000110100;
        biases1[49] <= 16'b0000000100010011;
        biases1[50] <= 16'b0000000010000101;
        biases1[51] <= 16'b1111111111111000;
        biases1[52] <= 16'b0000000010010001;
        biases1[53] <= 16'b1111111111110110;
        biases1[54] <= 16'b0000000000000000;
        biases1[55] <= 16'b0000000000000010;
        biases1[56] <= 16'b0000000001000000;
        biases1[57] <= 16'b0000000001001100;
        biases1[58] <= 16'b1111111110100001;
        biases1[59] <= 16'b0000000010010101;
        biases1[60] <= 16'b1111111111100010;
        biases1[61] <= 16'b0000000010100000;
        biases1[62] <= 16'b0000000000001000;
        biases1[63] <= 16'b1111111111101010;
        weights2[0] <= 16'b0000000000000001;
        weights2[1] <= 16'b1111111101101100;
        weights2[2] <= 16'b0000000000000100;
        weights2[3] <= 16'b1111111111001101;
        weights2[4] <= 16'b0000000000001001;
        weights2[5] <= 16'b1111111111110101;
        weights2[6] <= 16'b0000000000000000;
        weights2[7] <= 16'b1111111111110101;
        weights2[8] <= 16'b0000000000100011;
        weights2[9] <= 16'b0000000000010001;
        weights2[10] <= 16'b1111111110001011;
        weights2[11] <= 16'b0000000000001000;
        weights2[12] <= 16'b1111111111010001;
        weights2[13] <= 16'b1111111100110001;
        weights2[14] <= 16'b1111111110101110;
        weights2[15] <= 16'b0000000000011101;
        weights2[16] <= 16'b0000000000010111;
        weights2[17] <= 16'b0000000000110010;
        weights2[18] <= 16'b1111111111111001;
        weights2[19] <= 16'b1111111111110011;
        weights2[20] <= 16'b1111111110100001;
        weights2[21] <= 16'b0000000000011000;
        weights2[22] <= 16'b0000000000000011;
        weights2[23] <= 16'b0000000000001010;
        weights2[24] <= 16'b1111111110111010;
        weights2[25] <= 16'b0000000000000101;
        weights2[26] <= 16'b0000000000001111;
        weights2[27] <= 16'b1111111111010001;
        weights2[28] <= 16'b1111111111100111;
        weights2[29] <= 16'b0000000000000100;
        weights2[30] <= 16'b0000000000000111;
        weights2[31] <= 16'b1111111110011001;
        weights2[32] <= 16'b0000000000011001;
        weights2[33] <= 16'b0000000001000110;
        weights2[34] <= 16'b1111111110100111;
        weights2[35] <= 16'b1111111111100010;
        weights2[36] <= 16'b1111111111010101;
        weights2[37] <= 16'b1111111110011101;
        weights2[38] <= 16'b1111111111100100;
        weights2[39] <= 16'b1111111110011010;
        weights2[40] <= 16'b0000000000001000;
        weights2[41] <= 16'b1111111101100100;
        weights2[42] <= 16'b0000000000011101;
        weights2[43] <= 16'b1111111111001101;
        weights2[44] <= 16'b0000000000100011;
        weights2[45] <= 16'b0000000000101101;
        weights2[46] <= 16'b1111111111111010;
        weights2[47] <= 16'b1111111111110100;
        weights2[48] <= 16'b0000000000101011;
        weights2[49] <= 16'b0000000000100001;
        weights2[50] <= 16'b1111111111011100;
        weights2[51] <= 16'b0000000000001010;
        weights2[52] <= 16'b0000000000101111;
        weights2[53] <= 16'b1111111100100011;
        weights2[54] <= 16'b0000000000000000;
        weights2[55] <= 16'b0000000000010101;
        weights2[56] <= 16'b1111111100010100;
        weights2[57] <= 16'b1111111111101100;
        weights2[58] <= 16'b1111111101010011;
        weights2[59] <= 16'b1111111111111000;
        weights2[60] <= 16'b0000000000001000;
        weights2[61] <= 16'b0000000000011010;
        weights2[62] <= 16'b0000000000001111;
        weights2[63] <= 16'b1111111110001111;
        weights2[64] <= 16'b1111111111110101;
        weights2[65] <= 16'b0000000001100001;
        weights2[66] <= 16'b1111111111001110;
        weights2[67] <= 16'b1111111101111111;
        weights2[68] <= 16'b1111111110010110;
        weights2[69] <= 16'b0000000000001110;
        weights2[70] <= 16'b0000000000000000;
        weights2[71] <= 16'b0000000001110100;
        weights2[72] <= 16'b0000000000011010;
        weights2[73] <= 16'b1111111110110001;
        weights2[74] <= 16'b0000000000100100;
        weights2[75] <= 16'b1111111111111110;
        weights2[76] <= 16'b0000000001101100;
        weights2[77] <= 16'b0000000001111000;
        weights2[78] <= 16'b1111111111110100;
        weights2[79] <= 16'b0000000000001000;
        weights2[80] <= 16'b0000000000001000;
        weights2[81] <= 16'b1111111110110110;
        weights2[82] <= 16'b1111111111110001;
        weights2[83] <= 16'b1111111111010111;
        weights2[84] <= 16'b1111111110010000;
        weights2[85] <= 16'b1111111111010110;
        weights2[86] <= 16'b1111111111100101;
        weights2[87] <= 16'b1111111110110111;
        weights2[88] <= 16'b1111111110000001;
        weights2[89] <= 16'b1111111111110001;
        weights2[90] <= 16'b1111111110011011;
        weights2[91] <= 16'b0000000000100100;
        weights2[92] <= 16'b0000000010010011;
        weights2[93] <= 16'b1111111111100001;
        weights2[94] <= 16'b1111111111110001;
        weights2[95] <= 16'b1111111111111101;
        weights2[96] <= 16'b1111111111100101;
        weights2[97] <= 16'b1111111101111111;
        weights2[98] <= 16'b1111111110000111;
        weights2[99] <= 16'b1111111110110101;
        weights2[100] <= 16'b0000000001001110;
        weights2[101] <= 16'b1111111111110010;
        weights2[102] <= 16'b1111111111011011;
        weights2[103] <= 16'b0000000000010010;
        weights2[104] <= 16'b0000000000000000;
        weights2[105] <= 16'b0000000000110001;
        weights2[106] <= 16'b1111111111001100;
        weights2[107] <= 16'b1111111101010110;
        weights2[108] <= 16'b0000000000001000;
        weights2[109] <= 16'b1111111111011101;
        weights2[110] <= 16'b0000000001101101;
        weights2[111] <= 16'b0000000001001000;
        weights2[112] <= 16'b0000000000101100;
        weights2[113] <= 16'b1111111110111011;
        weights2[114] <= 16'b0000000001010011;
        weights2[115] <= 16'b0000000000000011;
        weights2[116] <= 16'b1111111111000011;
        weights2[117] <= 16'b0000000000010110;
        weights2[118] <= 16'b0000000000000000;
        weights2[119] <= 16'b1111111110111100;
        weights2[120] <= 16'b0000000001101100;
        weights2[121] <= 16'b1111111110101000;
        weights2[122] <= 16'b0000000000011111;
        weights2[123] <= 16'b1111111111011111;
        weights2[124] <= 16'b1111111111110010;
        weights2[125] <= 16'b1111111111011100;
        weights2[126] <= 16'b0000000000101111;
        weights2[127] <= 16'b1111111110111110;
        weights2[128] <= 16'b0000000001111111;
        weights2[129] <= 16'b1111111110100010;
        weights2[130] <= 16'b0000000000011100;
        weights2[131] <= 16'b0000000000000110;
        weights2[132] <= 16'b1111111101110100;
        weights2[133] <= 16'b0000000000001100;
        weights2[134] <= 16'b0000000000000000;
        weights2[135] <= 16'b1111111111110001;
        weights2[136] <= 16'b0000000001001000;
        weights2[137] <= 16'b1111111110101000;
        weights2[138] <= 16'b1111111111011001;
        weights2[139] <= 16'b1111111111100011;
        weights2[140] <= 16'b1111111111110100;
        weights2[141] <= 16'b1111111110011011;
        weights2[142] <= 16'b0000000000000101;
        weights2[143] <= 16'b0000000000101010;
        weights2[144] <= 16'b0000000000111101;
        weights2[145] <= 16'b0000000001011100;
        weights2[146] <= 16'b0000000000011010;
        weights2[147] <= 16'b0000000010000000;
        weights2[148] <= 16'b0000000000010000;
        weights2[149] <= 16'b0000000000111001;
        weights2[150] <= 16'b0000000001111111;
        weights2[151] <= 16'b0000000001010001;
        weights2[152] <= 16'b1111111111111011;
        weights2[153] <= 16'b0000000000010110;
        weights2[154] <= 16'b1111111101101000;
        weights2[155] <= 16'b0000000000111110;
        weights2[156] <= 16'b1111111110100100;
        weights2[157] <= 16'b1111111111111011;
        weights2[158] <= 16'b0000000001110101;
        weights2[159] <= 16'b1111111111111101;
        weights2[160] <= 16'b0000000000010111;
        weights2[161] <= 16'b1111111110010000;
        weights2[162] <= 16'b1111111111111110;
        weights2[163] <= 16'b1111111111011100;
        weights2[164] <= 16'b1111111111111010;
        weights2[165] <= 16'b1111111111111101;
        weights2[166] <= 16'b0000000000100000;
        weights2[167] <= 16'b1111111111001010;
        weights2[168] <= 16'b0000000000000000;
        weights2[169] <= 16'b1111111111101001;
        weights2[170] <= 16'b0000000000100111;
        weights2[171] <= 16'b0000000000000011;
        weights2[172] <= 16'b0000000000100001;
        weights2[173] <= 16'b0000000000000010;
        weights2[174] <= 16'b1111111110110000;
        weights2[175] <= 16'b1111111111011011;
        weights2[176] <= 16'b0000000001000110;
        weights2[177] <= 16'b0000000000110001;
        weights2[178] <= 16'b1111111111111011;
        weights2[179] <= 16'b1111111111111100;
        weights2[180] <= 16'b0000000001000101;
        weights2[181] <= 16'b1111111111011101;
        weights2[182] <= 16'b0000000000000000;
        weights2[183] <= 16'b1111111111001000;
        weights2[184] <= 16'b1111111111010001;
        weights2[185] <= 16'b1111111111111010;
        weights2[186] <= 16'b1111111111101111;
        weights2[187] <= 16'b0000000000000000;
        weights2[188] <= 16'b0000000000001001;
        weights2[189] <= 16'b0000000000011001;
        weights2[190] <= 16'b0000000000110001;
        weights2[191] <= 16'b1111111101010000;
        weights2[192] <= 16'b1111111111111111;
        weights2[193] <= 16'b1111111101111101;
        weights2[194] <= 16'b1111111111111011;
        weights2[195] <= 16'b1111111111100101;
        weights2[196] <= 16'b1111111111100100;
        weights2[197] <= 16'b1111111111001011;
        weights2[198] <= 16'b0000000000000000;
        weights2[199] <= 16'b1111111100011010;
        weights2[200] <= 16'b1111111111010111;
        weights2[201] <= 16'b1111111111111111;
        weights2[202] <= 16'b1111111110011101;
        weights2[203] <= 16'b1111111101011010;
        weights2[204] <= 16'b1111111111111111;
        weights2[205] <= 16'b1111111110000011;
        weights2[206] <= 16'b1111111101110010;
        weights2[207] <= 16'b0000000000001000;
        weights2[208] <= 16'b1111111111111100;
        weights2[209] <= 16'b1111111110001111;
        weights2[210] <= 16'b1111111110001000;
        weights2[211] <= 16'b1111111101111010;
        weights2[212] <= 16'b1111111111111111;
        weights2[213] <= 16'b1111111110101100;
        weights2[214] <= 16'b1111111110111001;
        weights2[215] <= 16'b1111111110010111;
        weights2[216] <= 16'b0000000000011110;
        weights2[217] <= 16'b0000000000001001;
        weights2[218] <= 16'b1111111111110011;
        weights2[219] <= 16'b1111111101010011;
        weights2[220] <= 16'b0000000000001111;
        weights2[221] <= 16'b0000000000010100;
        weights2[222] <= 16'b1111111111110000;
        weights2[223] <= 16'b1111111110010100;
        weights2[224] <= 16'b0000000000011000;
        weights2[225] <= 16'b1111111111111110;
        weights2[226] <= 16'b1111111111110100;
        weights2[227] <= 16'b1111111111111001;
        weights2[228] <= 16'b1111111100111110;
        weights2[229] <= 16'b1111111101111010;
        weights2[230] <= 16'b1111111111110110;
        weights2[231] <= 16'b1111111101111110;
        weights2[232] <= 16'b1111111111111010;
        weights2[233] <= 16'b1111111101111000;
        weights2[234] <= 16'b0000000000101111;
        weights2[235] <= 16'b0000000000100100;
        weights2[236] <= 16'b0000000000001010;
        weights2[237] <= 16'b0000000000010111;
        weights2[238] <= 16'b0000000000101011;
        weights2[239] <= 16'b1111111101111110;
        weights2[240] <= 16'b0000000000011010;
        weights2[241] <= 16'b0000000000100001;
        weights2[242] <= 16'b0000000000001011;
        weights2[243] <= 16'b0000000000010100;
        weights2[244] <= 16'b0000000000100011;
        weights2[245] <= 16'b1111111101100111;
        weights2[246] <= 16'b0000000000000000;
        weights2[247] <= 16'b0000000000010100;
        weights2[248] <= 16'b1111111110111101;
        weights2[249] <= 16'b0000000000110100;
        weights2[250] <= 16'b1111111101101010;
        weights2[251] <= 16'b0000000000011111;
        weights2[252] <= 16'b1111111111111110;
        weights2[253] <= 16'b0000000000011110;
        weights2[254] <= 16'b0000000000001010;
        weights2[255] <= 16'b1111111110001111;
        weights2[256] <= 16'b1111111111101001;
        weights2[257] <= 16'b1111111110011101;
        weights2[258] <= 16'b0000000000111010;
        weights2[259] <= 16'b0000000000100111;
        weights2[260] <= 16'b0000000000010110;
        weights2[261] <= 16'b0000000000011111;
        weights2[262] <= 16'b0000000000000000;
        weights2[263] <= 16'b1111111110000100;
        weights2[264] <= 16'b1111111110100101;
        weights2[265] <= 16'b0000000000000000;
        weights2[266] <= 16'b0000000000000011;
        weights2[267] <= 16'b0000000000001111;
        weights2[268] <= 16'b1111111101011011;
        weights2[269] <= 16'b1111111111000000;
        weights2[270] <= 16'b0000000001101110;
        weights2[271] <= 16'b1111111100111101;
        weights2[272] <= 16'b1111111111110011;
        weights2[273] <= 16'b0000000000011110;
        weights2[274] <= 16'b1111111111111111;
        weights2[275] <= 16'b0000000000010111;
        weights2[276] <= 16'b0000000000110110;
        weights2[277] <= 16'b0000000001000010;
        weights2[278] <= 16'b0000000000000101;
        weights2[279] <= 16'b1111111110111101;
        weights2[280] <= 16'b0000000000110000;
        weights2[281] <= 16'b0000000000001001;
        weights2[282] <= 16'b1111111111111010;
        weights2[283] <= 16'b1111111111100101;
        weights2[284] <= 16'b1111111111111001;
        weights2[285] <= 16'b0000000000000100;
        weights2[286] <= 16'b0000000000100011;
        weights2[287] <= 16'b0000000001011011;
        weights2[288] <= 16'b0000000000001000;
        weights2[289] <= 16'b1111111111011000;
        weights2[290] <= 16'b0000000000101010;
        weights2[291] <= 16'b1111111110001100;
        weights2[292] <= 16'b1111111110101010;
        weights2[293] <= 16'b0000000001100101;
        weights2[294] <= 16'b0000000000100001;
        weights2[295] <= 16'b0000000000101100;
        weights2[296] <= 16'b1111111111001001;
        weights2[297] <= 16'b0000000000011000;
        weights2[298] <= 16'b0000000000110001;
        weights2[299] <= 16'b0000000000101011;
        weights2[300] <= 16'b0000000000000111;
        weights2[301] <= 16'b1111111111100110;
        weights2[302] <= 16'b0000000000010000;
        weights2[303] <= 16'b1111111111010011;
        weights2[304] <= 16'b1111111100000001;
        weights2[305] <= 16'b0000000001000011;
        weights2[306] <= 16'b0000000000000010;
        weights2[307] <= 16'b0000000000000001;
        weights2[308] <= 16'b1111111111101101;
        weights2[309] <= 16'b0000000000111101;
        weights2[310] <= 16'b0000000000000000;
        weights2[311] <= 16'b1111111110001001;
        weights2[312] <= 16'b0000000000010001;
        weights2[313] <= 16'b0000000000101011;
        weights2[314] <= 16'b0000000000101001;
        weights2[315] <= 16'b0000000000000111;
        weights2[316] <= 16'b1111111111111011;
        weights2[317] <= 16'b0000000000011111;
        weights2[318] <= 16'b1111111011111000;
        weights2[319] <= 16'b1111111111111011;
        weights2[320] <= 16'b0000000000001111;
        weights2[321] <= 16'b1111111110101001;
        weights2[322] <= 16'b0000000001000010;
        weights2[323] <= 16'b0000000000110100;
        weights2[324] <= 16'b0000000000110101;
        weights2[325] <= 16'b0000000000010000;
        weights2[326] <= 16'b0000000000000000;
        weights2[327] <= 16'b1111111100001010;
        weights2[328] <= 16'b1111111111001010;
        weights2[329] <= 16'b0000000000001110;
        weights2[330] <= 16'b1111111110110001;
        weights2[331] <= 16'b0000000000010010;
        weights2[332] <= 16'b1111111110000001;
        weights2[333] <= 16'b1111111110101101;
        weights2[334] <= 16'b0000000001110000;
        weights2[335] <= 16'b1111111101101011;
        weights2[336] <= 16'b0000000000100001;
        weights2[337] <= 16'b1111111111110001;
        weights2[338] <= 16'b0000000000001001;
        weights2[339] <= 16'b0000000000100010;
        weights2[340] <= 16'b0000000000101110;
        weights2[341] <= 16'b0000000000111011;
        weights2[342] <= 16'b0000000000100000;
        weights2[343] <= 16'b1111111110100100;
        weights2[344] <= 16'b0000000000000001;
        weights2[345] <= 16'b0000000000010101;
        weights2[346] <= 16'b0000000000010100;
        weights2[347] <= 16'b1111111111011100;
        weights2[348] <= 16'b1111111100010110;
        weights2[349] <= 16'b1111111111011111;
        weights2[350] <= 16'b1111111111110101;
        weights2[351] <= 16'b0000000001011110;
        weights2[352] <= 16'b0000000000110110;
        weights2[353] <= 16'b0000000000001100;
        weights2[354] <= 16'b0000000000010010;
        weights2[355] <= 16'b1111111111101011;
        weights2[356] <= 16'b1111111100110001;
        weights2[357] <= 16'b0000000001110101;
        weights2[358] <= 16'b1111111111101000;
        weights2[359] <= 16'b0000000000010110;
        weights2[360] <= 16'b1111111111101110;
        weights2[361] <= 16'b0000000000000101;
        weights2[362] <= 16'b0000000001101000;
        weights2[363] <= 16'b1111111111110000;
        weights2[364] <= 16'b0000000000101100;
        weights2[365] <= 16'b0000000000000000;
        weights2[366] <= 16'b1111111101101101;
        weights2[367] <= 16'b1111111111011110;
        weights2[368] <= 16'b1111111111001110;
        weights2[369] <= 16'b0000000001011011;
        weights2[370] <= 16'b1111111110101110;
        weights2[371] <= 16'b0000000000000101;
        weights2[372] <= 16'b0000000000110010;
        weights2[373] <= 16'b0000000000110100;
        weights2[374] <= 16'b0000000000000000;
        weights2[375] <= 16'b1111111111111100;
        weights2[376] <= 16'b0000000000011010;
        weights2[377] <= 16'b1111111111111111;
        weights2[378] <= 16'b1111111111111101;
        weights2[379] <= 16'b0000000000010100;
        weights2[380] <= 16'b0000000000101101;
        weights2[381] <= 16'b0000000001000110;
        weights2[382] <= 16'b1111111111100100;
        weights2[383] <= 16'b0000000000001101;
        weights2[384] <= 16'b0000000000000110;
        weights2[385] <= 16'b0000000001000101;
        weights2[386] <= 16'b1111111111000010;
        weights2[387] <= 16'b0000000000000100;
        weights2[388] <= 16'b1111111111110001;
        weights2[389] <= 16'b1111111111010001;
        weights2[390] <= 16'b0000000000000000;
        weights2[391] <= 16'b1111111100101010;
        weights2[392] <= 16'b1111111101111110;
        weights2[393] <= 16'b0000000000100101;
        weights2[394] <= 16'b1111111110011010;
        weights2[395] <= 16'b1111111100010100;
        weights2[396] <= 16'b0000000000111010;
        weights2[397] <= 16'b0000000000111101;
        weights2[398] <= 16'b1111111111111111;
        weights2[399] <= 16'b1111111110111000;
        weights2[400] <= 16'b0000000000001111;
        weights2[401] <= 16'b1111111100111010;
        weights2[402] <= 16'b1111111101000111;
        weights2[403] <= 16'b1111111101000011;
        weights2[404] <= 16'b1111111111011001;
        weights2[405] <= 16'b1111111101101010;
        weights2[406] <= 16'b1111111110011010;
        weights2[407] <= 16'b1111111101010000;
        weights2[408] <= 16'b0000000000000101;
        weights2[409] <= 16'b1111111111110011;
        weights2[410] <= 16'b1111111111011010;
        weights2[411] <= 16'b1111111111000001;
        weights2[412] <= 16'b1111111101101110;
        weights2[413] <= 16'b0000000000000111;
        weights2[414] <= 16'b1111111110011111;
        weights2[415] <= 16'b1111111111111100;
        weights2[416] <= 16'b0000000000101010;
        weights2[417] <= 16'b1111111111110001;
        weights2[418] <= 16'b1111111111111001;
        weights2[419] <= 16'b1111111111111100;
        weights2[420] <= 16'b1111111110000001;
        weights2[421] <= 16'b0000000000000001;
        weights2[422] <= 16'b1111111111011000;
        weights2[423] <= 16'b1111111110011100;
        weights2[424] <= 16'b1111111111101100;
        weights2[425] <= 16'b1111111111110011;
        weights2[426] <= 16'b1111111111010111;
        weights2[427] <= 16'b0000000000010010;
        weights2[428] <= 16'b0000000000011100;
        weights2[429] <= 16'b0000000000011001;
        weights2[430] <= 16'b1111111111101000;
        weights2[431] <= 16'b1111111110100111;
        weights2[432] <= 16'b1111111111110011;
        weights2[433] <= 16'b1111111110100110;
        weights2[434] <= 16'b1111111111110101;
        weights2[435] <= 16'b0000000000001111;
        weights2[436] <= 16'b1111111110100001;
        weights2[437] <= 16'b0000000000001100;
        weights2[438] <= 16'b0000000000000000;
        weights2[439] <= 16'b0000000001000000;
        weights2[440] <= 16'b0000000000101010;
        weights2[441] <= 16'b0000000000001100;
        weights2[442] <= 16'b1111111101110101;
        weights2[443] <= 16'b0000000000010110;
        weights2[444] <= 16'b1111111111110011;
        weights2[445] <= 16'b1111111111111010;
        weights2[446] <= 16'b0000000000001100;
        weights2[447] <= 16'b0000000000101000;
        weights2[448] <= 16'b0000000000010101;
        weights2[449] <= 16'b1111111101011000;
        weights2[450] <= 16'b0000000000011000;
        weights2[451] <= 16'b1111111111111111;
        weights2[452] <= 16'b1111111100000011;
        weights2[453] <= 16'b1111111111101010;
        weights2[454] <= 16'b0000000000000000;
        weights2[455] <= 16'b1111111111011111;
        weights2[456] <= 16'b0000000001000001;
        weights2[457] <= 16'b1111111100110111;
        weights2[458] <= 16'b0000000000001011;
        weights2[459] <= 16'b1111111111100010;
        weights2[460] <= 16'b1111111101000110;
        weights2[461] <= 16'b1111111101101110;
        weights2[462] <= 16'b0000000000010010;
        weights2[463] <= 16'b1111111111100001;
        weights2[464] <= 16'b0000000000011101;
        weights2[465] <= 16'b0000000000110000;
        weights2[466] <= 16'b0000000000001101;
        weights2[467] <= 16'b0000000000000111;
        weights2[468] <= 16'b1111111111110001;
        weights2[469] <= 16'b0000000000101110;
        weights2[470] <= 16'b0000000000100101;
        weights2[471] <= 16'b0000000001000000;
        weights2[472] <= 16'b0000000000001011;
        weights2[473] <= 16'b0000000000001111;
        weights2[474] <= 16'b1111111100111101;
        weights2[475] <= 16'b1111111111001101;
        weights2[476] <= 16'b1111111110110101;
        weights2[477] <= 16'b1111111111111111;
        weights2[478] <= 16'b1111111111111111;
        weights2[479] <= 16'b0000000000001001;
        weights2[480] <= 16'b1111111111111010;
        weights2[481] <= 16'b1111111110010110;
        weights2[482] <= 16'b0000000000000000;
        weights2[483] <= 16'b1111111110101110;
        weights2[484] <= 16'b0000000000010001;
        weights2[485] <= 16'b0000000000010110;
        weights2[486] <= 16'b0000000000100001;
        weights2[487] <= 16'b1111111111100100;
        weights2[488] <= 16'b1111111111110011;
        weights2[489] <= 16'b1111111111101110;
        weights2[490] <= 16'b0000000000100110;
        weights2[491] <= 16'b0000000000001100;
        weights2[492] <= 16'b1111111111110001;
        weights2[493] <= 16'b0000000000000110;
        weights2[494] <= 16'b1111111111110010;
        weights2[495] <= 16'b1111111110000111;
        weights2[496] <= 16'b1111111111001101;
        weights2[497] <= 16'b0000000000100000;
        weights2[498] <= 16'b0000000000011110;
        weights2[499] <= 16'b0000000000000100;
        weights2[500] <= 16'b0000000000010000;
        weights2[501] <= 16'b1111111111111001;
        weights2[502] <= 16'b0000000000000000;
        weights2[503] <= 16'b1111111100011111;
        weights2[504] <= 16'b1111111110100111;
        weights2[505] <= 16'b0000000000001011;
        weights2[506] <= 16'b0000000000001110;
        weights2[507] <= 16'b0000000000010010;
        weights2[508] <= 16'b0000000000100001;
        weights2[509] <= 16'b0000000000011010;
        weights2[510] <= 16'b1111111111001110;
        weights2[511] <= 16'b1111111110011000;
        weights2[512] <= 16'b1111111111000101;
        weights2[513] <= 16'b0000000000011101;
        weights2[514] <= 16'b1111111111011000;
        weights2[515] <= 16'b1111111111000011;
        weights2[516] <= 16'b1111111111010101;
        weights2[517] <= 16'b1111111111001111;
        weights2[518] <= 16'b0000000000000000;
        weights2[519] <= 16'b0000000010110011;
        weights2[520] <= 16'b0000000000111001;
        weights2[521] <= 16'b1111111111110010;
        weights2[522] <= 16'b0000000001011111;
        weights2[523] <= 16'b0000000000000010;
        weights2[524] <= 16'b0000000000101111;
        weights2[525] <= 16'b0000000000011110;
        weights2[526] <= 16'b1111111110011111;
        weights2[527] <= 16'b0000000000001100;
        weights2[528] <= 16'b1111111111111111;
        weights2[529] <= 16'b0000000000011111;
        weights2[530] <= 16'b0000000000000011;
        weights2[531] <= 16'b0000000000010000;
        weights2[532] <= 16'b1111111101111111;
        weights2[533] <= 16'b1111111111011011;
        weights2[534] <= 16'b0000000000001000;
        weights2[535] <= 16'b0000000000010111;
        weights2[536] <= 16'b0000000000010010;
        weights2[537] <= 16'b1111111111011000;
        weights2[538] <= 16'b1111111111101000;
        weights2[539] <= 16'b0000000000011011;
        weights2[540] <= 16'b0000000010011100;
        weights2[541] <= 16'b0000000000011100;
        weights2[542] <= 16'b0000000000001000;
        weights2[543] <= 16'b1111111111000001;
        weights2[544] <= 16'b1111111110101111;
        weights2[545] <= 16'b0000000000010100;
        weights2[546] <= 16'b1111111110110010;
        weights2[547] <= 16'b1111111111110100;
        weights2[548] <= 16'b0000000001000100;
        weights2[549] <= 16'b1111111101100110;
        weights2[550] <= 16'b1111111111111010;
        weights2[551] <= 16'b1111111110101100;
        weights2[552] <= 16'b0000000000000000;
        weights2[553] <= 16'b0000000000101111;
        weights2[554] <= 16'b1111111110101011;
        weights2[555] <= 16'b0000000000010100;
        weights2[556] <= 16'b1111111111001000;
        weights2[557] <= 16'b0000000000000101;
        weights2[558] <= 16'b0000000010001111;
        weights2[559] <= 16'b0000000000001011;
        weights2[560] <= 16'b0000000000010010;
        weights2[561] <= 16'b1111111111000000;
        weights2[562] <= 16'b0000000010011100;
        weights2[563] <= 16'b1111111111110010;
        weights2[564] <= 16'b1111111110101110;
        weights2[565] <= 16'b1111111110110111;
        weights2[566] <= 16'b1111111111111111;
        weights2[567] <= 16'b1111111111001011;
        weights2[568] <= 16'b0000000000000010;
        weights2[569] <= 16'b0000000000001011;
        weights2[570] <= 16'b0000000000011110;
        weights2[571] <= 16'b1111111111001000;
        weights2[572] <= 16'b1111111111100100;
        weights2[573] <= 16'b1111111111011011;
        weights2[574] <= 16'b0000000000010101;
        weights2[575] <= 16'b1111111101000011;
        weights2[576] <= 16'b0000000000001100;
        weights2[577] <= 16'b1111111110010101;
        weights2[578] <= 16'b0000000001001001;
        weights2[579] <= 16'b0000000000111010;
        weights2[580] <= 16'b0000000000110111;
        weights2[581] <= 16'b0000000000010110;
        weights2[582] <= 16'b0000000000000000;
        weights2[583] <= 16'b0000000000111000;
        weights2[584] <= 16'b0000000000100111;
        weights2[585] <= 16'b0000000000010111;
        weights2[586] <= 16'b1111111111100011;
        weights2[587] <= 16'b0000000001001001;
        weights2[588] <= 16'b1111111110001001;
        weights2[589] <= 16'b1111111110101111;
        weights2[590] <= 16'b0000000000101010;
        weights2[591] <= 16'b1111111111100111;
        weights2[592] <= 16'b1111111111111011;
        weights2[593] <= 16'b0000000010001011;
        weights2[594] <= 16'b0000000000110111;
        weights2[595] <= 16'b0000000000111110;
        weights2[596] <= 16'b1111111101011110;
        weights2[597] <= 16'b0000000001111100;
        weights2[598] <= 16'b0000000001001110;
        weights2[599] <= 16'b0000000000101111;
        weights2[600] <= 16'b0000000000101001;
        weights2[601] <= 16'b1111111111111101;
        weights2[602] <= 16'b0000000001001001;
        weights2[603] <= 16'b0000000000000010;
        weights2[604] <= 16'b0000000000010111;
        weights2[605] <= 16'b1111111111111001;
        weights2[606] <= 16'b0000000000101011;
        weights2[607] <= 16'b0000000000100100;
        weights2[608] <= 16'b1111111111111110;
        weights2[609] <= 16'b0000000010100010;
        weights2[610] <= 16'b0000000000011000;
        weights2[611] <= 16'b1111111111000001;
        weights2[612] <= 16'b0000000000001100;
        weights2[613] <= 16'b0000000000110000;
        weights2[614] <= 16'b0000000000110100;
        weights2[615] <= 16'b0000000000110011;
        weights2[616] <= 16'b1111111111011001;
        weights2[617] <= 16'b1111111111001110;
        weights2[618] <= 16'b0000000000100100;
        weights2[619] <= 16'b0000000000111110;
        weights2[620] <= 16'b0000000000000010;
        weights2[621] <= 16'b0000000000001101;
        weights2[622] <= 16'b0000000000001010;
        weights2[623] <= 16'b0000000000000001;
        weights2[624] <= 16'b1111111111101001;
        weights2[625] <= 16'b0000000000011001;
        weights2[626] <= 16'b0000000000001011;
        weights2[627] <= 16'b1111111111010001;
        weights2[628] <= 16'b0000000001001001;
        weights2[629] <= 16'b0000000000110010;
        weights2[630] <= 16'b0000000000000000;
        weights2[631] <= 16'b0000000000101111;
        weights2[632] <= 16'b1111111110111001;
        weights2[633] <= 16'b0000000000100001;
        weights2[634] <= 16'b1111111111001111;
        weights2[635] <= 16'b0000000000000111;
        weights2[636] <= 16'b1111111111100010;
        weights2[637] <= 16'b0000000000011001;
        weights2[638] <= 16'b1111111111110111;
        weights2[639] <= 16'b0000000001000111;
        weights2[640] <= 16'b0000000000011011;
        weights2[641] <= 16'b0000000001101000;
        weights2[642] <= 16'b1111111111010110;
        weights2[643] <= 16'b1111111110010100;
        weights2[644] <= 16'b1111111111110011;
        weights2[645] <= 16'b0000000000001001;
        weights2[646] <= 16'b0000000000000000;
        weights2[647] <= 16'b0000000000010011;
        weights2[648] <= 16'b0000000000011011;
        weights2[649] <= 16'b0000000000001000;
        weights2[650] <= 16'b0000000000010100;
        weights2[651] <= 16'b0000000001111100;
        weights2[652] <= 16'b0000000001000001;
        weights2[653] <= 16'b0000000001101101;
        weights2[654] <= 16'b0000000000111000;
        weights2[655] <= 16'b1111111111111101;
        weights2[656] <= 16'b0000000000110101;
        weights2[657] <= 16'b0000000000111110;
        weights2[658] <= 16'b0000000001110101;
        weights2[659] <= 16'b0000000001010111;
        weights2[660] <= 16'b0000000000100000;
        weights2[661] <= 16'b0000000000111100;
        weights2[662] <= 16'b0000000001111011;
        weights2[663] <= 16'b0000000000101101;
        weights2[664] <= 16'b1111111101011010;
        weights2[665] <= 16'b1111111111110000;
        weights2[666] <= 16'b0000000000000100;
        weights2[667] <= 16'b0000000010111001;
        weights2[668] <= 16'b1111111111100111;
        weights2[669] <= 16'b1111111110110110;
        weights2[670] <= 16'b1111111111110001;
        weights2[671] <= 16'b0000000000110110;
        weights2[672] <= 16'b0000000000000100;
        weights2[673] <= 16'b1111111111100000;
        weights2[674] <= 16'b1111111110100000;
        weights2[675] <= 16'b1111111110101001;
        weights2[676] <= 16'b0000000000100101;
        weights2[677] <= 16'b0000000000110001;
        weights2[678] <= 16'b1111111111100000;
        weights2[679] <= 16'b1111111111111101;
        weights2[680] <= 16'b1111111111111001;
        weights2[681] <= 16'b0000000000011011;
        weights2[682] <= 16'b1111111111100110;
        weights2[683] <= 16'b1111111101101111;
        weights2[684] <= 16'b1111111111111011;
        weights2[685] <= 16'b1111111111010101;
        weights2[686] <= 16'b0000000000011100;
        weights2[687] <= 16'b0000000001110000;
        weights2[688] <= 16'b1111111111110000;
        weights2[689] <= 16'b1111111111110010;
        weights2[690] <= 16'b0000000000100110;
        weights2[691] <= 16'b1111111111100101;
        weights2[692] <= 16'b1111111111111101;
        weights2[693] <= 16'b0000000000010110;
        weights2[694] <= 16'b0000000000000000;
        weights2[695] <= 16'b1111111111110110;
        weights2[696] <= 16'b0000000000110100;
        weights2[697] <= 16'b1111111110001101;
        weights2[698] <= 16'b0000000000000010;
        weights2[699] <= 16'b1111111111101001;
        weights2[700] <= 16'b0000000001000001;
        weights2[701] <= 16'b1111111111110000;
        weights2[702] <= 16'b1111111111110001;
        weights2[703] <= 16'b1111111111010101;
        weights2[704] <= 16'b0000000000000100;
        weights2[705] <= 16'b1111111101111111;
        weights2[706] <= 16'b1111111111100000;
        weights2[707] <= 16'b1111111111001001;
        weights2[708] <= 16'b0000000000010101;
        weights2[709] <= 16'b1111111111101111;
        weights2[710] <= 16'b0000000000000000;
        weights2[711] <= 16'b0000000000010010;
        weights2[712] <= 16'b0000000000111111;
        weights2[713] <= 16'b0000000000000100;
        weights2[714] <= 16'b1111111111001101;
        weights2[715] <= 16'b1111111111111011;
        weights2[716] <= 16'b1111111111000011;
        weights2[717] <= 16'b1111111101011101;
        weights2[718] <= 16'b1111111110010001;
        weights2[719] <= 16'b1111111111101010;
        weights2[720] <= 16'b0000000000100101;
        weights2[721] <= 16'b1111111111010110;
        weights2[722] <= 16'b0000000000001000;
        weights2[723] <= 16'b1111111111011111;
        weights2[724] <= 16'b1111111100100011;
        weights2[725] <= 16'b0000000000001011;
        weights2[726] <= 16'b0000000000011110;
        weights2[727] <= 16'b0000000000101110;
        weights2[728] <= 16'b1111111111100000;
        weights2[729] <= 16'b1111111111001110;
        weights2[730] <= 16'b0000000000001010;
        weights2[731] <= 16'b1111111110000111;
        weights2[732] <= 16'b1111111111000001;
        weights2[733] <= 16'b1111111110110000;
        weights2[734] <= 16'b1111111110101011;
        weights2[735] <= 16'b1111111110010001;
        weights2[736] <= 16'b1111111111010111;
        weights2[737] <= 16'b0000000000110100;
        weights2[738] <= 16'b1111111111000111;
        weights2[739] <= 16'b0000000000001010;
        weights2[740] <= 16'b0000000000101100;
        weights2[741] <= 16'b1111111111000101;
        weights2[742] <= 16'b1111111111101000;
        weights2[743] <= 16'b1111111111010111;
        weights2[744] <= 16'b0000000000001001;
        weights2[745] <= 16'b1111111111110110;
        weights2[746] <= 16'b1111111101101100;
        weights2[747] <= 16'b1111111111100010;
        weights2[748] <= 16'b1111111111110010;
        weights2[749] <= 16'b0000000000001100;
        weights2[750] <= 16'b1111111111111000;
        weights2[751] <= 16'b1111111111010100;
        weights2[752] <= 16'b1111111111111010;
        weights2[753] <= 16'b1111111111000011;
        weights2[754] <= 16'b1111111111100101;
        weights2[755] <= 16'b0000000000000000;
        weights2[756] <= 16'b1111111111110101;
        weights2[757] <= 16'b1111111111100001;
        weights2[758] <= 16'b0000000000000000;
        weights2[759] <= 16'b1111111111001000;
        weights2[760] <= 16'b1111111110111111;
        weights2[761] <= 16'b1111111111010111;
        weights2[762] <= 16'b1111111111111010;
        weights2[763] <= 16'b1111111111000010;
        weights2[764] <= 16'b1111111111011101;
        weights2[765] <= 16'b1111111110111110;
        weights2[766] <= 16'b0000000000001111;
        weights2[767] <= 16'b0000000000100011;
        weights2[768] <= 16'b1111111101111001;
        weights2[769] <= 16'b0000000000000101;
        weights2[770] <= 16'b0000000001010011;
        weights2[771] <= 16'b0000000000111001;
        weights2[772] <= 16'b1111111111111111;
        weights2[773] <= 16'b1111111101100000;
        weights2[774] <= 16'b0000000000000000;
        weights2[775] <= 16'b0000000000100001;
        weights2[776] <= 16'b0000000000011000;
        weights2[777] <= 16'b1111111111100100;
        weights2[778] <= 16'b1111111111100001;
        weights2[779] <= 16'b0000000000100001;
        weights2[780] <= 16'b1111111111101111;
        weights2[781] <= 16'b0000000000001100;
        weights2[782] <= 16'b0000000000011011;
        weights2[783] <= 16'b0000000000000100;
        weights2[784] <= 16'b1111111111100100;
        weights2[785] <= 16'b0000000000100111;
        weights2[786] <= 16'b0000000000001000;
        weights2[787] <= 16'b0000000000001001;
        weights2[788] <= 16'b0000000000011111;
        weights2[789] <= 16'b0000000001101011;
        weights2[790] <= 16'b1111111111011010;
        weights2[791] <= 16'b0000000000001010;
        weights2[792] <= 16'b0000000010111111;
        weights2[793] <= 16'b0000000000110101;
        weights2[794] <= 16'b0000000000011110;
        weights2[795] <= 16'b0000000000101011;
        weights2[796] <= 16'b0000000000101010;
        weights2[797] <= 16'b0000000010001110;
        weights2[798] <= 16'b0000000000000000;
        weights2[799] <= 16'b0000000000011011;
        weights2[800] <= 16'b1111111111010100;
        weights2[801] <= 16'b0000000000000001;
        weights2[802] <= 16'b0000000001000000;
        weights2[803] <= 16'b0000000001100101;
        weights2[804] <= 16'b1111111111110110;
        weights2[805] <= 16'b0000000000010111;
        weights2[806] <= 16'b0000000000011011;
        weights2[807] <= 16'b0000000000001110;
        weights2[808] <= 16'b1111111111100010;
        weights2[809] <= 16'b0000000000001001;
        weights2[810] <= 16'b0000000001001100;
        weights2[811] <= 16'b0000000010011011;
        weights2[812] <= 16'b1111111110101011;
        weights2[813] <= 16'b0000000001001111;
        weights2[814] <= 16'b0000000000101111;
        weights2[815] <= 16'b0000000000100101;
        weights2[816] <= 16'b0000000000100100;
        weights2[817] <= 16'b0000000001110111;
        weights2[818] <= 16'b0000000001101101;
        weights2[819] <= 16'b0000000000011001;
        weights2[820] <= 16'b0000000000111011;
        weights2[821] <= 16'b0000000000011000;
        weights2[822] <= 16'b0000000000000000;
        weights2[823] <= 16'b0000000000001000;
        weights2[824] <= 16'b0000000000001100;
        weights2[825] <= 16'b0000000010010111;
        weights2[826] <= 16'b1111111111100011;
        weights2[827] <= 16'b0000000000100000;
        weights2[828] <= 16'b0000000000100000;
        weights2[829] <= 16'b0000000001011111;
        weights2[830] <= 16'b0000000000111001;
        weights2[831] <= 16'b1111111111101101;
        weights2[832] <= 16'b1111111111011100;
        weights2[833] <= 16'b1111111101111111;
        weights2[834] <= 16'b0000000000000111;
        weights2[835] <= 16'b0000000000101001;
        weights2[836] <= 16'b1111111110100011;
        weights2[837] <= 16'b1111111111111100;
        weights2[838] <= 16'b0000000000000000;
        weights2[839] <= 16'b1111111111110110;
        weights2[840] <= 16'b0000000000010000;
        weights2[841] <= 16'b1111111110010010;
        weights2[842] <= 16'b0000000000010111;
        weights2[843] <= 16'b1111111111001110;
        weights2[844] <= 16'b1111111110001011;
        weights2[845] <= 16'b1111111110100100;
        weights2[846] <= 16'b0000000000000110;
        weights2[847] <= 16'b1111111111111101;
        weights2[848] <= 16'b1111111111111110;
        weights2[849] <= 16'b1111111110110111;
        weights2[850] <= 16'b1111111111001011;
        weights2[851] <= 16'b1111111110101101;
        weights2[852] <= 16'b1111111110100011;
        weights2[853] <= 16'b1111111110111111;
        weights2[854] <= 16'b1111111110110111;
        weights2[855] <= 16'b0000000000001001;
        weights2[856] <= 16'b1111111111111111;
        weights2[857] <= 16'b1111111111111110;
        weights2[858] <= 16'b1111111110011100;
        weights2[859] <= 16'b1111111110000100;
        weights2[860] <= 16'b1111111111000101;
        weights2[861] <= 16'b1111111111110111;
        weights2[862] <= 16'b1111111111010110;
        weights2[863] <= 16'b1111111111111111;
        weights2[864] <= 16'b1111111111101111;
        weights2[865] <= 16'b1111111111001001;
        weights2[866] <= 16'b0000000000000111;
        weights2[867] <= 16'b1111111111001000;
        weights2[868] <= 16'b0000000000011101;
        weights2[869] <= 16'b0000000000001100;
        weights2[870] <= 16'b0000000000010111;
        weights2[871] <= 16'b1111111111110111;
        weights2[872] <= 16'b0000000000001011;
        weights2[873] <= 16'b1111111111111111;
        weights2[874] <= 16'b1111111111010101;
        weights2[875] <= 16'b0000000000100110;
        weights2[876] <= 16'b1111111111110010;
        weights2[877] <= 16'b0000000000101011;
        weights2[878] <= 16'b1111111111001010;
        weights2[879] <= 16'b1111111110111001;
        weights2[880] <= 16'b1111111111010010;
        weights2[881] <= 16'b1111111111110100;
        weights2[882] <= 16'b1111111110101001;
        weights2[883] <= 16'b0000000000001101;
        weights2[884] <= 16'b1111111101111011;
        weights2[885] <= 16'b1111111111101001;
        weights2[886] <= 16'b0000000000000000;
        weights2[887] <= 16'b1111111110110101;
        weights2[888] <= 16'b1111111110011101;
        weights2[889] <= 16'b0000000000101011;
        weights2[890] <= 16'b0000000000100110;
        weights2[891] <= 16'b1111111111000101;
        weights2[892] <= 16'b1111111110110111;
        weights2[893] <= 16'b1111111111110101;
        weights2[894] <= 16'b1111111110101101;
        weights2[895] <= 16'b1111111111111010;
        weights2[896] <= 16'b0000000000000111;
        weights2[897] <= 16'b1111111111101000;
        weights2[898] <= 16'b1111111110100011;
        weights2[899] <= 16'b1111111101111000;
        weights2[900] <= 16'b1111111111010010;
        weights2[901] <= 16'b1111111110100010;
        weights2[902] <= 16'b0000000000000000;
        weights2[903] <= 16'b1111111111111100;
        weights2[904] <= 16'b1111111110100110;
        weights2[905] <= 16'b1111111111101100;
        weights2[906] <= 16'b1111111111000100;
        weights2[907] <= 16'b1111111110101010;
        weights2[908] <= 16'b1111111111101010;
        weights2[909] <= 16'b1111111111100100;
        weights2[910] <= 16'b0000000000000110;
        weights2[911] <= 16'b0000000000000010;
        weights2[912] <= 16'b0000000001001101;
        weights2[913] <= 16'b1111111110101100;
        weights2[914] <= 16'b1111111111000011;
        weights2[915] <= 16'b1111111110110001;
        weights2[916] <= 16'b0000000001100011;
        weights2[917] <= 16'b1111111111101100;
        weights2[918] <= 16'b1111111111101110;
        weights2[919] <= 16'b1111111111100110;
        weights2[920] <= 16'b1111111101011011;
        weights2[921] <= 16'b0000000000100011;
        weights2[922] <= 16'b1111111110111111;
        weights2[923] <= 16'b1111111111001110;
        weights2[924] <= 16'b0000000001001100;
        weights2[925] <= 16'b1111111110110010;
        weights2[926] <= 16'b1111111110011101;
        weights2[927] <= 16'b0000000000000111;
        weights2[928] <= 16'b0000000000010100;
        weights2[929] <= 16'b1111111110110011;
        weights2[930] <= 16'b1111111110000111;
        weights2[931] <= 16'b1111111110001100;
        weights2[932] <= 16'b1111111111011001;
        weights2[933] <= 16'b0000000000000010;
        weights2[934] <= 16'b1111111111001000;
        weights2[935] <= 16'b1111111111110011;
        weights2[936] <= 16'b1111111111110111;
        weights2[937] <= 16'b0000000000001101;
        weights2[938] <= 16'b0000000000011111;
        weights2[939] <= 16'b1111111101101100;
        weights2[940] <= 16'b0000000000011100;
        weights2[941] <= 16'b1111111111010010;
        weights2[942] <= 16'b0000000001010000;
        weights2[943] <= 16'b1111111111011101;
        weights2[944] <= 16'b1111111111100011;
        weights2[945] <= 16'b0000000000101010;
        weights2[946] <= 16'b0000000000001100;
        weights2[947] <= 16'b0000000000010110;
        weights2[948] <= 16'b0000000000011111;
        weights2[949] <= 16'b0000000000001011;
        weights2[950] <= 16'b0000000000000000;
        weights2[951] <= 16'b1111111111101101;
        weights2[952] <= 16'b0000000000000011;
        weights2[953] <= 16'b1111111101111110;
        weights2[954] <= 16'b0000000000000010;
        weights2[955] <= 16'b0000000001001011;
        weights2[956] <= 16'b0000000010000010;
        weights2[957] <= 16'b0000000000010110;
        weights2[958] <= 16'b1111111111010000;
        weights2[959] <= 16'b1111111111010110;
        weights2[960] <= 16'b1111111111000101;
        weights2[961] <= 16'b1111111101000011;
        weights2[962] <= 16'b0000000000011101;
        weights2[963] <= 16'b0000000000011110;
        weights2[964] <= 16'b0000000000001000;
        weights2[965] <= 16'b0000000000100000;
        weights2[966] <= 16'b0000000000000000;
        weights2[967] <= 16'b1111111111111010;
        weights2[968] <= 16'b0000000000000011;
        weights2[969] <= 16'b0000000000000001;
        weights2[970] <= 16'b0000000000000101;
        weights2[971] <= 16'b1111111101001010;
        weights2[972] <= 16'b1111111110111111;
        weights2[973] <= 16'b1111111101111001;
        weights2[974] <= 16'b0000000000001001;
        weights2[975] <= 16'b0000000000010101;
        weights2[976] <= 16'b1111111101100111;
        weights2[977] <= 16'b0000000000111001;
        weights2[978] <= 16'b1111111101000101;
        weights2[979] <= 16'b1111111110100110;
        weights2[980] <= 16'b1111111110110111;
        weights2[981] <= 16'b0000000001100000;
        weights2[982] <= 16'b1111111101000111;
        weights2[983] <= 16'b1111111111111111;
        weights2[984] <= 16'b0000000000111001;
        weights2[985] <= 16'b1111111111011010;
        weights2[986] <= 16'b1111111111111010;
        weights2[987] <= 16'b1111111110001101;
        weights2[988] <= 16'b0000000000110000;
        weights2[989] <= 16'b0000000000101111;
        weights2[990] <= 16'b0000000001011101;
        weights2[991] <= 16'b0000000000000010;
        weights2[992] <= 16'b1111111111111100;
        weights2[993] <= 16'b0000000000001011;
        weights2[994] <= 16'b0000000000010011;
        weights2[995] <= 16'b1111111111111001;
        weights2[996] <= 16'b0000000000000101;
        weights2[997] <= 16'b0000000000001010;
        weights2[998] <= 16'b0000000001001010;
        weights2[999] <= 16'b1111111101111100;
        weights2[1000] <= 16'b1111111111010111;
        weights2[1001] <= 16'b1111111101111011;
        weights2[1002] <= 16'b1111111111110010;
        weights2[1003] <= 16'b0000000000110101;
        weights2[1004] <= 16'b1111111111101101;
        weights2[1005] <= 16'b0000000000101000;
        weights2[1006] <= 16'b0000000000110011;
        weights2[1007] <= 16'b1111111100111100;
        weights2[1008] <= 16'b0000000000010010;
        weights2[1009] <= 16'b0000000000101010;
        weights2[1010] <= 16'b0000000000100110;
        weights2[1011] <= 16'b1111111111010110;
        weights2[1012] <= 16'b1111111110100000;
        weights2[1013] <= 16'b1111111101110010;
        weights2[1014] <= 16'b0000000000000000;
        weights2[1015] <= 16'b1111111111110110;
        weights2[1016] <= 16'b1111111110000011;
        weights2[1017] <= 16'b0000000000110110;
        weights2[1018] <= 16'b1111111111100010;
        weights2[1019] <= 16'b1111111101110001;
        weights2[1020] <= 16'b1111111101000010;
        weights2[1021] <= 16'b0000000000010111;
        weights2[1022] <= 16'b1111111111111000;
        weights2[1023] <= 16'b0000000000100110;
        weights2[1024] <= 16'b0000000000010010;
        weights2[1025] <= 16'b0000000001101100;
        weights2[1026] <= 16'b0000000001010010;
        weights2[1027] <= 16'b0000000000101111;
        weights2[1028] <= 16'b1111111101111010;
        weights2[1029] <= 16'b0000000000110000;
        weights2[1030] <= 16'b0000000000000000;
        weights2[1031] <= 16'b0000000000110101;
        weights2[1032] <= 16'b1111111111011110;
        weights2[1033] <= 16'b1111111110100000;
        weights2[1034] <= 16'b0000000000010011;
        weights2[1035] <= 16'b0000000000100110;
        weights2[1036] <= 16'b0000000001000110;
        weights2[1037] <= 16'b0000000010000000;
        weights2[1038] <= 16'b0000000001011011;
        weights2[1039] <= 16'b1111111110111011;
        weights2[1040] <= 16'b1111111111100110;
        weights2[1041] <= 16'b0000000000100110;
        weights2[1042] <= 16'b0000000000001111;
        weights2[1043] <= 16'b0000000000011011;
        weights2[1044] <= 16'b0000000001010001;
        weights2[1045] <= 16'b0000000001001010;
        weights2[1046] <= 16'b0000000000001100;
        weights2[1047] <= 16'b1111111111010000;
        weights2[1048] <= 16'b0000000000101011;
        weights2[1049] <= 16'b0000000000010110;
        weights2[1050] <= 16'b1111111110101011;
        weights2[1051] <= 16'b0000000001000101;
        weights2[1052] <= 16'b0000000001011111;
        weights2[1053] <= 16'b0000000000111000;
        weights2[1054] <= 16'b0000000001000111;
        weights2[1055] <= 16'b0000000001000110;
        weights2[1056] <= 16'b0000000000000101;
        weights2[1057] <= 16'b1111111101111101;
        weights2[1058] <= 16'b0000000000101000;
        weights2[1059] <= 16'b1111111101100101;
        weights2[1060] <= 16'b0000000000110111;
        weights2[1061] <= 16'b0000000001001111;
        weights2[1062] <= 16'b0000000000101001;
        weights2[1063] <= 16'b0000000000101001;
        weights2[1064] <= 16'b1111111110101111;
        weights2[1065] <= 16'b0000000000001101;
        weights2[1066] <= 16'b0000000000000100;
        weights2[1067] <= 16'b0000000000011101;
        weights2[1068] <= 16'b0000000000000111;
        weights2[1069] <= 16'b1111111111111111;
        weights2[1070] <= 16'b0000000000111010;
        weights2[1071] <= 16'b0000000001011000;
        weights2[1072] <= 16'b1111111111001101;
        weights2[1073] <= 16'b0000000000101001;
        weights2[1074] <= 16'b0000000001010101;
        weights2[1075] <= 16'b1111111111100001;
        weights2[1076] <= 16'b1111111111110000;
        weights2[1077] <= 16'b0000000000101000;
        weights2[1078] <= 16'b0000000000000000;
        weights2[1079] <= 16'b1111111110000110;
        weights2[1080] <= 16'b0000000001111001;
        weights2[1081] <= 16'b0000000000011011;
        weights2[1082] <= 16'b0000000000011001;
        weights2[1083] <= 16'b0000000000001011;
        weights2[1084] <= 16'b0000000000001101;
        weights2[1085] <= 16'b0000000000101000;
        weights2[1086] <= 16'b1111111110101110;
        weights2[1087] <= 16'b1111111110110011;
        weights2[1088] <= 16'b1111111110110110;
        weights2[1089] <= 16'b0000000000000100;
        weights2[1090] <= 16'b1111111111001011;
        weights2[1091] <= 16'b1111111111110100;
        weights2[1092] <= 16'b0000000001101111;
        weights2[1093] <= 16'b1111111111110100;
        weights2[1094] <= 16'b0000000000000000;
        weights2[1095] <= 16'b1111111110110110;
        weights2[1096] <= 16'b1111111101111100;
        weights2[1097] <= 16'b0000000000101110;
        weights2[1098] <= 16'b1111111111111010;
        weights2[1099] <= 16'b1111111110101110;
        weights2[1100] <= 16'b1111111111010010;
        weights2[1101] <= 16'b0000000000011011;
        weights2[1102] <= 16'b0000000000100000;
        weights2[1103] <= 16'b1111111100101001;
        weights2[1104] <= 16'b1111111111100110;
        weights2[1105] <= 16'b1111111101110110;
        weights2[1106] <= 16'b1111111101101110;
        weights2[1107] <= 16'b1111111110010100;
        weights2[1108] <= 16'b1111111111011001;
        weights2[1109] <= 16'b1111111101111110;
        weights2[1110] <= 16'b1111111110011110;
        weights2[1111] <= 16'b1111111101001111;
        weights2[1112] <= 16'b0000000000001010;
        weights2[1113] <= 16'b1111111111011011;
        weights2[1114] <= 16'b0000000000011110;
        weights2[1115] <= 16'b1111111110111000;
        weights2[1116] <= 16'b1111111111100111;
        weights2[1117] <= 16'b1111111111110111;
        weights2[1118] <= 16'b1111111110100111;
        weights2[1119] <= 16'b0000000000100000;
        weights2[1120] <= 16'b1111111111110011;
        weights2[1121] <= 16'b0000000000011100;
        weights2[1122] <= 16'b1111111111111001;
        weights2[1123] <= 16'b1111111111000000;
        weights2[1124] <= 16'b1111111111111100;
        weights2[1125] <= 16'b0000000000110100;
        weights2[1126] <= 16'b1111111111100001;
        weights2[1127] <= 16'b0000000000111000;
        weights2[1128] <= 16'b1111111111011001;
        weights2[1129] <= 16'b0000000000011000;
        weights2[1130] <= 16'b1111111110111101;
        weights2[1131] <= 16'b0000000000000101;
        weights2[1132] <= 16'b1111111111111100;
        weights2[1133] <= 16'b1111111111111110;
        weights2[1134] <= 16'b0000000000000000;
        weights2[1135] <= 16'b1111111111101101;
        weights2[1136] <= 16'b1111111101000000;
        weights2[1137] <= 16'b1111111110111010;
        weights2[1138] <= 16'b1111111111111010;
        weights2[1139] <= 16'b0000000000000100;
        weights2[1140] <= 16'b1111111111010000;
        weights2[1141] <= 16'b0000000000000111;
        weights2[1142] <= 16'b0000000000000000;
        weights2[1143] <= 16'b1111111111111000;
        weights2[1144] <= 16'b0000000000011000;
        weights2[1145] <= 16'b1111111111111100;
        weights2[1146] <= 16'b1111111111110101;
        weights2[1147] <= 16'b1111111111000101;
        weights2[1148] <= 16'b1111111111100010;
        weights2[1149] <= 16'b1111111111010011;
        weights2[1150] <= 16'b1111111110000000;
        weights2[1151] <= 16'b0000000000100000;
        weights2[1152] <= 16'b0000000001110100;
        weights2[1153] <= 16'b0000000001101101;
        weights2[1154] <= 16'b1111111111111010;
        weights2[1155] <= 16'b0000000000000011;
        weights2[1156] <= 16'b1111111111110110;
        weights2[1157] <= 16'b0000000000100111;
        weights2[1158] <= 16'b0000000000000000;
        weights2[1159] <= 16'b1111111110110001;
        weights2[1160] <= 16'b0000000000000101;
        weights2[1161] <= 16'b1111111111111100;
        weights2[1162] <= 16'b1111111111101100;
        weights2[1163] <= 16'b0000000000111110;
        weights2[1164] <= 16'b0000000001101011;
        weights2[1165] <= 16'b0000000001101110;
        weights2[1166] <= 16'b1111111111101011;
        weights2[1167] <= 16'b0000000000001001;
        weights2[1168] <= 16'b0000000001000101;
        weights2[1169] <= 16'b0000000000010101;
        weights2[1170] <= 16'b0000000000111110;
        weights2[1171] <= 16'b0000000000110001;
        weights2[1172] <= 16'b0000000000000011;
        weights2[1173] <= 16'b0000000001000110;
        weights2[1174] <= 16'b0000000001011101;
        weights2[1175] <= 16'b1111111111100001;
        weights2[1176] <= 16'b1111111111011110;
        weights2[1177] <= 16'b0000000000110000;
        weights2[1178] <= 16'b0000000000000011;
        weights2[1179] <= 16'b0000000001011011;
        weights2[1180] <= 16'b1111111111011010;
        weights2[1181] <= 16'b1111111111110001;
        weights2[1182] <= 16'b0000000001000011;
        weights2[1183] <= 16'b1111111111100110;
        weights2[1184] <= 16'b0000000001001010;
        weights2[1185] <= 16'b1111111111111101;
        weights2[1186] <= 16'b1111111111101110;
        weights2[1187] <= 16'b0000000000001110;
        weights2[1188] <= 16'b1111111101111011;
        weights2[1189] <= 16'b1111111110110111;
        weights2[1190] <= 16'b1111111111100110;
        weights2[1191] <= 16'b1111111111010000;
        weights2[1192] <= 16'b1111111111101001;
        weights2[1193] <= 16'b0000000000000101;
        weights2[1194] <= 16'b0000000000101001;
        weights2[1195] <= 16'b1111111111001011;
        weights2[1196] <= 16'b0000000001001001;
        weights2[1197] <= 16'b1111111111111101;
        weights2[1198] <= 16'b1111111111101101;
        weights2[1199] <= 16'b0000000010000101;
        weights2[1200] <= 16'b0000000000101010;
        weights2[1201] <= 16'b0000000001010110;
        weights2[1202] <= 16'b1111111111111010;
        weights2[1203] <= 16'b1111111111110111;
        weights2[1204] <= 16'b0000000010000011;
        weights2[1205] <= 16'b0000000000010101;
        weights2[1206] <= 16'b0000000000000000;
        weights2[1207] <= 16'b0000000000001111;
        weights2[1208] <= 16'b0000000001010000;
        weights2[1209] <= 16'b1111111111011110;
        weights2[1210] <= 16'b1111111110110111;
        weights2[1211] <= 16'b0000000000101110;
        weights2[1212] <= 16'b0000000001111101;
        weights2[1213] <= 16'b0000000000110001;
        weights2[1214] <= 16'b0000000000101101;
        weights2[1215] <= 16'b1111111111110000;
        weights2[1216] <= 16'b1111111111110011;
        weights2[1217] <= 16'b0000000000010100;
        weights2[1218] <= 16'b0000000000101110;
        weights2[1219] <= 16'b0000000010001001;
        weights2[1220] <= 16'b0000000000110101;
        weights2[1221] <= 16'b0000000000010011;
        weights2[1222] <= 16'b0000000000000000;
        weights2[1223] <= 16'b1111111111011000;
        weights2[1224] <= 16'b0000000001101001;
        weights2[1225] <= 16'b0000000000001001;
        weights2[1226] <= 16'b0000000000000010;
        weights2[1227] <= 16'b0000000000010011;
        weights2[1228] <= 16'b0000000000000011;
        weights2[1229] <= 16'b0000000000011010;
        weights2[1230] <= 16'b0000000000001001;
        weights2[1231] <= 16'b0000000000000010;
        weights2[1232] <= 16'b1111111111010100;
        weights2[1233] <= 16'b0000000000010101;
        weights2[1234] <= 16'b0000000000000010;
        weights2[1235] <= 16'b1111111111111011;
        weights2[1236] <= 16'b1111111110101011;
        weights2[1237] <= 16'b0000000000101110;
        weights2[1238] <= 16'b0000000000001111;
        weights2[1239] <= 16'b0000000001001110;
        weights2[1240] <= 16'b0000000010000101;
        weights2[1241] <= 16'b1111111110111110;
        weights2[1242] <= 16'b0000000000111010;
        weights2[1243] <= 16'b0000000000101001;
        weights2[1244] <= 16'b1111111101111101;
        weights2[1245] <= 16'b0000000000110011;
        weights2[1246] <= 16'b0000000000111010;
        weights2[1247] <= 16'b0000000000010000;
        weights2[1248] <= 16'b0000000000001000;
        weights2[1249] <= 16'b0000000001001000;
        weights2[1250] <= 16'b0000000001110110;
        weights2[1251] <= 16'b0000000001011101;
        weights2[1252] <= 16'b0000000000011010;
        weights2[1253] <= 16'b0000000000000111;
        weights2[1254] <= 16'b0000000000100101;
        weights2[1255] <= 16'b0000000000000100;
        weights2[1256] <= 16'b1111111111111101;
        weights2[1257] <= 16'b0000000000000000;
        weights2[1258] <= 16'b1111111111110000;
        weights2[1259] <= 16'b0000000010000101;
        weights2[1260] <= 16'b0000000000001000;
        weights2[1261] <= 16'b0000000000001111;
        weights2[1262] <= 16'b1111111101010011;
        weights2[1263] <= 16'b0000000000110010;
        weights2[1264] <= 16'b0000000000001100;
        weights2[1265] <= 16'b1111111111111100;
        weights2[1266] <= 16'b1111111110100101;
        weights2[1267] <= 16'b1111111111010011;
        weights2[1268] <= 16'b0000000000001010;
        weights2[1269] <= 16'b1111111111110110;
        weights2[1270] <= 16'b0000000000000000;
        weights2[1271] <= 16'b0000000000100111;
        weights2[1272] <= 16'b0000000000100110;
        weights2[1273] <= 16'b0000000001101101;
        weights2[1274] <= 16'b1111111111110011;
        weights2[1275] <= 16'b1111111110101111;
        weights2[1276] <= 16'b1111111110100110;
        weights2[1277] <= 16'b1111111111100000;
        weights2[1278] <= 16'b0000000000110000;
        weights2[1279] <= 16'b0000000000011011;
        weights2[1280] <= 16'b1111111111001000;
        weights2[1281] <= 16'b1111111111101111;
        weights2[1282] <= 16'b1111111111001011;
        weights2[1283] <= 16'b1111111101100011;
        weights2[1284] <= 16'b1111111111101011;
        weights2[1285] <= 16'b1111111110010111;
        weights2[1286] <= 16'b0000000000000000;
        weights2[1287] <= 16'b0000000000110110;
        weights2[1288] <= 16'b0000000000100110;
        weights2[1289] <= 16'b1111111111110011;
        weights2[1290] <= 16'b1111111110010001;
        weights2[1291] <= 16'b1111111110011110;
        weights2[1292] <= 16'b1111111111111011;
        weights2[1293] <= 16'b1111111111110011;
        weights2[1294] <= 16'b1111111110011001;
        weights2[1295] <= 16'b0000000000000010;
        weights2[1296] <= 16'b0000000000000000;
        weights2[1297] <= 16'b1111111110101110;
        weights2[1298] <= 16'b1111111110100001;
        weights2[1299] <= 16'b1111111110111011;
        weights2[1300] <= 16'b1111111111011110;
        weights2[1301] <= 16'b1111111110100001;
        weights2[1302] <= 16'b1111111110100000;
        weights2[1303] <= 16'b0000000000001111;
        weights2[1304] <= 16'b1111111111011011;
        weights2[1305] <= 16'b0000000000100101;
        weights2[1306] <= 16'b1111111111101100;
        weights2[1307] <= 16'b1111111111101111;
        weights2[1308] <= 16'b0000000001010101;
        weights2[1309] <= 16'b0000000001001011;
        weights2[1310] <= 16'b1111111110001110;
        weights2[1311] <= 16'b1111111101110010;
        weights2[1312] <= 16'b1111111111000000;
        weights2[1313] <= 16'b1111111111111000;
        weights2[1314] <= 16'b1111111100001011;
        weights2[1315] <= 16'b0000000000011010;
        weights2[1316] <= 16'b0000000001010000;
        weights2[1317] <= 16'b1111111110111010;
        weights2[1318] <= 16'b1111111110110010;
        weights2[1319] <= 16'b1111111111010010;
        weights2[1320] <= 16'b1111111111111000;
        weights2[1321] <= 16'b1111111111111111;
        weights2[1322] <= 16'b0000000000100110;
        weights2[1323] <= 16'b0000000000010111;
        weights2[1324] <= 16'b1111111110110100;
        weights2[1325] <= 16'b0000000001100001;
        weights2[1326] <= 16'b0000000001111001;
        weights2[1327] <= 16'b1111111111100110;
        weights2[1328] <= 16'b0000000000001100;
        weights2[1329] <= 16'b0000000000111000;
        weights2[1330] <= 16'b0000000001101111;
        weights2[1331] <= 16'b0000000000110100;
        weights2[1332] <= 16'b1111111111110001;
        weights2[1333] <= 16'b0000000000000011;
        weights2[1334] <= 16'b0000000000000000;
        weights2[1335] <= 16'b1111111111110001;
        weights2[1336] <= 16'b1111111111101011;
        weights2[1337] <= 16'b0000000000000101;
        weights2[1338] <= 16'b0000000000000001;
        weights2[1339] <= 16'b0000000000001010;
        weights2[1340] <= 16'b0000000000001100;
        weights2[1341] <= 16'b0000000000111010;
        weights2[1342] <= 16'b0000000000010001;
        weights2[1343] <= 16'b0000000000000011;
        weights2[1344] <= 16'b1111111100110100;
        weights2[1345] <= 16'b1111111111111011;
        weights2[1346] <= 16'b1111111110111111;
        weights2[1347] <= 16'b1111111111101011;
        weights2[1348] <= 16'b0000000000011100;
        weights2[1349] <= 16'b1111111110010111;
        weights2[1350] <= 16'b0000000000000000;
        weights2[1351] <= 16'b0000000000101011;
        weights2[1352] <= 16'b0000000000011110;
        weights2[1353] <= 16'b0000000000001100;
        weights2[1354] <= 16'b0000000000100111;
        weights2[1355] <= 16'b1111111110000100;
        weights2[1356] <= 16'b0000000000000110;
        weights2[1357] <= 16'b0000000000011100;
        weights2[1358] <= 16'b0000000000000001;
        weights2[1359] <= 16'b0000000000000101;
        weights2[1360] <= 16'b1111111111000100;
        weights2[1361] <= 16'b1111111111111000;
        weights2[1362] <= 16'b1111111100111111;
        weights2[1363] <= 16'b1111111110110011;
        weights2[1364] <= 16'b1111111110010111;
        weights2[1365] <= 16'b1111111110110011;
        weights2[1366] <= 16'b1111111100011111;
        weights2[1367] <= 16'b0000000000010101;
        weights2[1368] <= 16'b0000000000100010;
        weights2[1369] <= 16'b1111111111001110;
        weights2[1370] <= 16'b0000000000100110;
        weights2[1371] <= 16'b1111111111101001;
        weights2[1372] <= 16'b0000000010000111;
        weights2[1373] <= 16'b0000000000101001;
        weights2[1374] <= 16'b1111111101111000;
        weights2[1375] <= 16'b0000000000001101;
        weights2[1376] <= 16'b1111111110100100;
        weights2[1377] <= 16'b0000000000100000;
        weights2[1378] <= 16'b0000000000000001;
        weights2[1379] <= 16'b1111111111100010;
        weights2[1380] <= 16'b1111111110011101;
        weights2[1381] <= 16'b1111111111111010;
        weights2[1382] <= 16'b1111111111111010;
        weights2[1383] <= 16'b0000000000101110;
        weights2[1384] <= 16'b1111111111111010;
        weights2[1385] <= 16'b0000000000110101;
        weights2[1386] <= 16'b1111111111011111;
        weights2[1387] <= 16'b0000000000101110;
        weights2[1388] <= 16'b1111111110000110;
        weights2[1389] <= 16'b0000000000101011;
        weights2[1390] <= 16'b0000000010010001;
        weights2[1391] <= 16'b1111111111110001;
        weights2[1392] <= 16'b1111111111111001;
        weights2[1393] <= 16'b1111111111010100;
        weights2[1394] <= 16'b0000000001101001;
        weights2[1395] <= 16'b0000000000001011;
        weights2[1396] <= 16'b1111111110101100;
        weights2[1397] <= 16'b0000000000001110;
        weights2[1398] <= 16'b1111111111111111;
        weights2[1399] <= 16'b1111111111111101;
        weights2[1400] <= 16'b0000000000011000;
        weights2[1401] <= 16'b0000000000101010;
        weights2[1402] <= 16'b0000000000000101;
        weights2[1403] <= 16'b1111111110101101;
        weights2[1404] <= 16'b1111111111101101;
        weights2[1405] <= 16'b1111111111110100;
        weights2[1406] <= 16'b1111111111110000;
        weights2[1407] <= 16'b0000000000010011;
        weights2[1408] <= 16'b0000000000000100;
        weights2[1409] <= 16'b1111111110101110;
        weights2[1410] <= 16'b1111111110011011;
        weights2[1411] <= 16'b1111111111100000;
        weights2[1412] <= 16'b1111111110111001;
        weights2[1413] <= 16'b1111111111100011;
        weights2[1414] <= 16'b0000000000000000;
        weights2[1415] <= 16'b0000000000101010;
        weights2[1416] <= 16'b1111111111100110;
        weights2[1417] <= 16'b1111111111101010;
        weights2[1418] <= 16'b0000000000001110;
        weights2[1419] <= 16'b0000000000000000;
        weights2[1420] <= 16'b1111111111111011;
        weights2[1421] <= 16'b0000000000101010;
        weights2[1422] <= 16'b1111111101010111;
        weights2[1423] <= 16'b0000000001011101;
        weights2[1424] <= 16'b1111111111111000;
        weights2[1425] <= 16'b1111111110000100;
        weights2[1426] <= 16'b0000000000001010;
        weights2[1427] <= 16'b1111111111110100;
        weights2[1428] <= 16'b1111111111011011;
        weights2[1429] <= 16'b1111111111011011;
        weights2[1430] <= 16'b1111111111111111;
        weights2[1431] <= 16'b1111111110101000;
        weights2[1432] <= 16'b1111111111011011;
        weights2[1433] <= 16'b1111111111111101;
        weights2[1434] <= 16'b1111111111011000;
        weights2[1435] <= 16'b1111111110110100;
        weights2[1436] <= 16'b0000000001111111;
        weights2[1437] <= 16'b0000000000001110;
        weights2[1438] <= 16'b1111111111111000;
        weights2[1439] <= 16'b1111111110000110;
        weights2[1440] <= 16'b0000000000000111;
        weights2[1441] <= 16'b0000000000000100;
        weights2[1442] <= 16'b1111111111001101;
        weights2[1443] <= 16'b0000000010110110;
        weights2[1444] <= 16'b1111111111100001;
        weights2[1445] <= 16'b1111111101010011;
        weights2[1446] <= 16'b1111111111000001;
        weights2[1447] <= 16'b1111111111110010;
        weights2[1448] <= 16'b0000000000001111;
        weights2[1449] <= 16'b1111111111101111;
        weights2[1450] <= 16'b1111111111110011;
        weights2[1451] <= 16'b1111111111101010;
        weights2[1452] <= 16'b1111111111111111;
        weights2[1453] <= 16'b1111111111111100;
        weights2[1454] <= 16'b0000000000110001;
        weights2[1455] <= 16'b0000000000011010;
        weights2[1456] <= 16'b0000000010011110;
        weights2[1457] <= 16'b1111111111000011;
        weights2[1458] <= 16'b0000000000100000;
        weights2[1459] <= 16'b0000000000011000;
        weights2[1460] <= 16'b1111111111011000;
        weights2[1461] <= 16'b1111111111000011;
        weights2[1462] <= 16'b0000000000000000;
        weights2[1463] <= 16'b1111111111100001;
        weights2[1464] <= 16'b1111111111010100;
        weights2[1465] <= 16'b1111111111100110;
        weights2[1466] <= 16'b1111111111110101;
        weights2[1467] <= 16'b0000000000000101;
        weights2[1468] <= 16'b1111111111011111;
        weights2[1469] <= 16'b1111111111111001;
        weights2[1470] <= 16'b0000000001111100;
        weights2[1471] <= 16'b1111111110101111;
        weights2[1472] <= 16'b0000000000101011;
        weights2[1473] <= 16'b1111111111111001;
        weights2[1474] <= 16'b0000000000011010;
        weights2[1475] <= 16'b1111111110001010;
        weights2[1476] <= 16'b1111111110001111;
        weights2[1477] <= 16'b0000000001001100;
        weights2[1478] <= 16'b0000000000000000;
        weights2[1479] <= 16'b1111111111101010;
        weights2[1480] <= 16'b1111111111110101;
        weights2[1481] <= 16'b1111111111101100;
        weights2[1482] <= 16'b1111111111100100;
        weights2[1483] <= 16'b1111111111111011;
        weights2[1484] <= 16'b1111111111110110;
        weights2[1485] <= 16'b0000000000000000;
        weights2[1486] <= 16'b0000000000010100;
        weights2[1487] <= 16'b0000000000000011;
        weights2[1488] <= 16'b0000000000101110;
        weights2[1489] <= 16'b0000000000001100;
        weights2[1490] <= 16'b1111111111111001;
        weights2[1491] <= 16'b0000000000100110;
        weights2[1492] <= 16'b0000000000000111;
        weights2[1493] <= 16'b1111111111110001;
        weights2[1494] <= 16'b0000000000010011;
        weights2[1495] <= 16'b1111111111100010;
        weights2[1496] <= 16'b1111111110010101;
        weights2[1497] <= 16'b1111111110111111;
        weights2[1498] <= 16'b1111111101111011;
        weights2[1499] <= 16'b1111111111110001;
        weights2[1500] <= 16'b1111111111001111;
        weights2[1501] <= 16'b1111111110000011;
        weights2[1502] <= 16'b0000000001001001;
        weights2[1503] <= 16'b0000000000000110;
        weights2[1504] <= 16'b0000000001100111;
        weights2[1505] <= 16'b1111111101000110;
        weights2[1506] <= 16'b1111111111001100;
        weights2[1507] <= 16'b1111111100110101;
        weights2[1508] <= 16'b1111111111011110;
        weights2[1509] <= 16'b0000000000001000;
        weights2[1510] <= 16'b0000000000010100;
        weights2[1511] <= 16'b1111111111110111;
        weights2[1512] <= 16'b1111111111101111;
        weights2[1513] <= 16'b0000000000000010;
        weights2[1514] <= 16'b1111111111101011;
        weights2[1515] <= 16'b1111111101101110;
        weights2[1516] <= 16'b0000000001100110;
        weights2[1517] <= 16'b1111111110101010;
        weights2[1518] <= 16'b1111111111000101;
        weights2[1519] <= 16'b1111111111110001;
        weights2[1520] <= 16'b1111111111110101;
        weights2[1521] <= 16'b1111111111010011;
        weights2[1522] <= 16'b1111111110111001;
        weights2[1523] <= 16'b1111111111101000;
        weights2[1524] <= 16'b1111111111101010;
        weights2[1525] <= 16'b1111111111111111;
        weights2[1526] <= 16'b0000000000000000;
        weights2[1527] <= 16'b1111111111010010;
        weights2[1528] <= 16'b1111111111110111;
        weights2[1529] <= 16'b1111111110010000;
        weights2[1530] <= 16'b0000000000000000;
        weights2[1531] <= 16'b1111111111101101;
        weights2[1532] <= 16'b0000000000011100;
        weights2[1533] <= 16'b1111111110100101;
        weights2[1534] <= 16'b1111111110100110;
        weights2[1535] <= 16'b1111111111100101;
        weights2[1536] <= 16'b0000000000010100;
        weights2[1537] <= 16'b1111111111100111;
        weights2[1538] <= 16'b0000000001100001;
        weights2[1539] <= 16'b0000000001111001;
        weights2[1540] <= 16'b0000000000010001;
        weights2[1541] <= 16'b0000000000000111;
        weights2[1542] <= 16'b0000000000000000;
        weights2[1543] <= 16'b1111111110100001;
        weights2[1544] <= 16'b0000000000001101;
        weights2[1545] <= 16'b0000000000001111;
        weights2[1546] <= 16'b1111111100011011;
        weights2[1547] <= 16'b1111111111111101;
        weights2[1548] <= 16'b1111111111111000;
        weights2[1549] <= 16'b1111111110111001;
        weights2[1550] <= 16'b0000000000000101;
        weights2[1551] <= 16'b0000000000010001;
        weights2[1552] <= 16'b1111111111110111;
        weights2[1553] <= 16'b0000000000011110;
        weights2[1554] <= 16'b1111111111110000;
        weights2[1555] <= 16'b0000000000000100;
        weights2[1556] <= 16'b1111111111001000;
        weights2[1557] <= 16'b0000000000110010;
        weights2[1558] <= 16'b1111111111101110;
        weights2[1559] <= 16'b0000000000001000;
        weights2[1560] <= 16'b0000000001101011;
        weights2[1561] <= 16'b0000000000010110;
        weights2[1562] <= 16'b0000000000100110;
        weights2[1563] <= 16'b1111111111111101;
        weights2[1564] <= 16'b1111111110001101;
        weights2[1565] <= 16'b0000000000111101;
        weights2[1566] <= 16'b0000000000011111;
        weights2[1567] <= 16'b1111111111111000;
        weights2[1568] <= 16'b0000000000011111;
        weights2[1569] <= 16'b0000000000010101;
        weights2[1570] <= 16'b0000000001100110;
        weights2[1571] <= 16'b0000000001100111;
        weights2[1572] <= 16'b1111111110110101;
        weights2[1573] <= 16'b1111111111111000;
        weights2[1574] <= 16'b0000000000011110;
        weights2[1575] <= 16'b1111111110011100;
        weights2[1576] <= 16'b1111111111111011;
        weights2[1577] <= 16'b1111111111001000;
        weights2[1578] <= 16'b0000000000100111;
        weights2[1579] <= 16'b0000000010000001;
        weights2[1580] <= 16'b0000000000100001;
        weights2[1581] <= 16'b0000000001010000;
        weights2[1582] <= 16'b1111111110100000;
        weights2[1583] <= 16'b1111111111010111;
        weights2[1584] <= 16'b0000000000110111;
        weights2[1585] <= 16'b0000000001001100;
        weights2[1586] <= 16'b1111111111000101;
        weights2[1587] <= 16'b1111111111111011;
        weights2[1588] <= 16'b1111111111100110;
        weights2[1589] <= 16'b0000000000000011;
        weights2[1590] <= 16'b0000000000000000;
        weights2[1591] <= 16'b0000000001001001;
        weights2[1592] <= 16'b0000000000000000;
        weights2[1593] <= 16'b0000000001111111;
        weights2[1594] <= 16'b1111111110011110;
        weights2[1595] <= 16'b0000000000010100;
        weights2[1596] <= 16'b1111111111001001;
        weights2[1597] <= 16'b0000000000101101;
        weights2[1598] <= 16'b0000000001010011;
        weights2[1599] <= 16'b0000000000011110;
        weights2[1600] <= 16'b1111111110110000;
        weights2[1601] <= 16'b1111111111001111;
        weights2[1602] <= 16'b1111111111111111;
        weights2[1603] <= 16'b0000000000100110;
        weights2[1604] <= 16'b0000000000000100;
        weights2[1605] <= 16'b1111111111101101;
        weights2[1606] <= 16'b0000000000000000;
        weights2[1607] <= 16'b1111111111101010;
        weights2[1608] <= 16'b1111111111111110;
        weights2[1609] <= 16'b0000000000010010;
        weights2[1610] <= 16'b1111111111110110;
        weights2[1611] <= 16'b1111111101111111;
        weights2[1612] <= 16'b1111111111000011;
        weights2[1613] <= 16'b1111111111101000;
        weights2[1614] <= 16'b0000000000111100;
        weights2[1615] <= 16'b1111111111110101;
        weights2[1616] <= 16'b0000000000000110;
        weights2[1617] <= 16'b1111111110110100;
        weights2[1618] <= 16'b1111111110000010;
        weights2[1619] <= 16'b1111111110100010;
        weights2[1620] <= 16'b0000000000000100;
        weights2[1621] <= 16'b1111111111010010;
        weights2[1622] <= 16'b1111111101111100;
        weights2[1623] <= 16'b0000000000011100;
        weights2[1624] <= 16'b1111111111111111;
        weights2[1625] <= 16'b1111111110111100;
        weights2[1626] <= 16'b1111111111110110;
        weights2[1627] <= 16'b1111111110110001;
        weights2[1628] <= 16'b1111111110101111;
        weights2[1629] <= 16'b1111111111110010;
        weights2[1630] <= 16'b1111111110110101;
        weights2[1631] <= 16'b0000000000101100;
        weights2[1632] <= 16'b1111111111111000;
        weights2[1633] <= 16'b1111111111011011;
        weights2[1634] <= 16'b0000000000011110;
        weights2[1635] <= 16'b1111111110010111;
        weights2[1636] <= 16'b0000000000101000;
        weights2[1637] <= 16'b0000000000111011;
        weights2[1638] <= 16'b1111111111101111;
        weights2[1639] <= 16'b1111111101011110;
        weights2[1640] <= 16'b1111111111110011;
        weights2[1641] <= 16'b0000000000111010;
        weights2[1642] <= 16'b1111111110010111;
        weights2[1643] <= 16'b1111111111101001;
        weights2[1644] <= 16'b1111111111111001;
        weights2[1645] <= 16'b0000000000001011;
        weights2[1646] <= 16'b1111111110011000;
        weights2[1647] <= 16'b1111111110101010;
        weights2[1648] <= 16'b1111111111000110;
        weights2[1649] <= 16'b1111111111010111;
        weights2[1650] <= 16'b1111111110101001;
        weights2[1651] <= 16'b1111111111110010;
        weights2[1652] <= 16'b1111111110000011;
        weights2[1653] <= 16'b0000000000100101;
        weights2[1654] <= 16'b0000000000000000;
        weights2[1655] <= 16'b1111111111101001;
        weights2[1656] <= 16'b1111111111111100;
        weights2[1657] <= 16'b1111111111110011;
        weights2[1658] <= 16'b0000000000110001;
        weights2[1659] <= 16'b1111111110100101;
        weights2[1660] <= 16'b1111111111101001;
        weights2[1661] <= 16'b1111111110110110;
        weights2[1662] <= 16'b1111111110101011;
        weights2[1663] <= 16'b1111111111100010;
        weights2[1664] <= 16'b1111111111110010;
        weights2[1665] <= 16'b0000000000111001;
        weights2[1666] <= 16'b1111111111111111;
        weights2[1667] <= 16'b0000000001101111;
        weights2[1668] <= 16'b1111111111100000;
        weights2[1669] <= 16'b0000000000010011;
        weights2[1670] <= 16'b0000000000000000;
        weights2[1671] <= 16'b1111111111111001;
        weights2[1672] <= 16'b1111111111110111;
        weights2[1673] <= 16'b1111111111101100;
        weights2[1674] <= 16'b0000000000111111;
        weights2[1675] <= 16'b1111111111010001;
        weights2[1676] <= 16'b0000000000100101;
        weights2[1677] <= 16'b0000000000111000;
        weights2[1678] <= 16'b0000000000000111;
        weights2[1679] <= 16'b0000000000000011;
        weights2[1680] <= 16'b1111111111111100;
        weights2[1681] <= 16'b1111111111101000;
        weights2[1682] <= 16'b1111111111100100;
        weights2[1683] <= 16'b1111111111011011;
        weights2[1684] <= 16'b1111111110110101;
        weights2[1685] <= 16'b1111111111011000;
        weights2[1686] <= 16'b1111111111101101;
        weights2[1687] <= 16'b1111111111101001;
        weights2[1688] <= 16'b0000000001011101;
        weights2[1689] <= 16'b1111111110000001;
        weights2[1690] <= 16'b1111111111100011;
        weights2[1691] <= 16'b0000000000000010;
        weights2[1692] <= 16'b1111111111000100;
        weights2[1693] <= 16'b1111111111110100;
        weights2[1694] <= 16'b0000000000110010;
        weights2[1695] <= 16'b0000000000010001;
        weights2[1696] <= 16'b0000000000011110;
        weights2[1697] <= 16'b1111111111110100;
        weights2[1698] <= 16'b0000000001101110;
        weights2[1699] <= 16'b1111111111001001;
        weights2[1700] <= 16'b1111111111011000;
        weights2[1701] <= 16'b0000000000000100;
        weights2[1702] <= 16'b0000000000010111;
        weights2[1703] <= 16'b0000000000010011;
        weights2[1704] <= 16'b1111111111110110;
        weights2[1705] <= 16'b0000000000110011;
        weights2[1706] <= 16'b1111111110110001;
        weights2[1707] <= 16'b0000000000110010;
        weights2[1708] <= 16'b0000000000010111;
        weights2[1709] <= 16'b1111111111010000;
        weights2[1710] <= 16'b1111111101001011;
        weights2[1711] <= 16'b0000000000010111;
        weights2[1712] <= 16'b0000000000011011;
        weights2[1713] <= 16'b1111111110101101;
        weights2[1714] <= 16'b1111111100111110;
        weights2[1715] <= 16'b1111111111101100;
        weights2[1716] <= 16'b1111111111000000;
        weights2[1717] <= 16'b0000000000000000;
        weights2[1718] <= 16'b0000000000000000;
        weights2[1719] <= 16'b1111111111101110;
        weights2[1720] <= 16'b0000000001010100;
        weights2[1721] <= 16'b0000000000110010;
        weights2[1722] <= 16'b0000000001001011;
        weights2[1723] <= 16'b1111111110011001;
        weights2[1724] <= 16'b1111111111001011;
        weights2[1725] <= 16'b1111111101000110;
        weights2[1726] <= 16'b0000000000000101;
        weights2[1727] <= 16'b1111111111000000;
        weights2[1728] <= 16'b1111111111100110;
        weights2[1729] <= 16'b0000000001010010;
        weights2[1730] <= 16'b1111111111011000;
        weights2[1731] <= 16'b0000000000010011;
        weights2[1732] <= 16'b1111111110000001;
        weights2[1733] <= 16'b1111111111100101;
        weights2[1734] <= 16'b0000000000000000;
        weights2[1735] <= 16'b0000000000100111;
        weights2[1736] <= 16'b1111111111011110;
        weights2[1737] <= 16'b1111111111111011;
        weights2[1738] <= 16'b0000000000010011;
        weights2[1739] <= 16'b0000000001010100;
        weights2[1740] <= 16'b0000000000010101;
        weights2[1741] <= 16'b0000000001111001;
        weights2[1742] <= 16'b0000000000011110;
        weights2[1743] <= 16'b1111111111100110;
        weights2[1744] <= 16'b0000000000010001;
        weights2[1745] <= 16'b1111111111110111;
        weights2[1746] <= 16'b0000000000101100;
        weights2[1747] <= 16'b0000000001011101;
        weights2[1748] <= 16'b0000000001001101;
        weights2[1749] <= 16'b1111111111101000;
        weights2[1750] <= 16'b0000000000110010;
        weights2[1751] <= 16'b1111111110011000;
        weights2[1752] <= 16'b0000000000000111;
        weights2[1753] <= 16'b0000000000001010;
        weights2[1754] <= 16'b0000000000001101;
        weights2[1755] <= 16'b0000000001011010;
        weights2[1756] <= 16'b0000000001001111;
        weights2[1757] <= 16'b0000000000000011;
        weights2[1758] <= 16'b0000000000110100;
        weights2[1759] <= 16'b0000000000100011;
        weights2[1760] <= 16'b1111111111111100;
        weights2[1761] <= 16'b0000000000000001;
        weights2[1762] <= 16'b0000000000010011;
        weights2[1763] <= 16'b1111111101010000;
        weights2[1764] <= 16'b1111111111111111;
        weights2[1765] <= 16'b0000000000100100;
        weights2[1766] <= 16'b1111111111011101;
        weights2[1767] <= 16'b0000000010000110;
        weights2[1768] <= 16'b1111111111111110;
        weights2[1769] <= 16'b0000000000110111;
        weights2[1770] <= 16'b0000000000001000;
        weights2[1771] <= 16'b1111111111111101;
        weights2[1772] <= 16'b1111111111001010;
        weights2[1773] <= 16'b1111111111101100;
        weights2[1774] <= 16'b0000000000010111;
        weights2[1775] <= 16'b0000000010011101;
        weights2[1776] <= 16'b1111111111010111;
        weights2[1777] <= 16'b1111111111110110;
        weights2[1778] <= 16'b1111111111110111;
        weights2[1779] <= 16'b0000000000001101;
        weights2[1780] <= 16'b0000000000010101;
        weights2[1781] <= 16'b0000000001100001;
        weights2[1782] <= 16'b0000000000000000;
        weights2[1783] <= 16'b1111111110111100;
        weights2[1784] <= 16'b0000000010000010;
        weights2[1785] <= 16'b0000000000000101;
        weights2[1786] <= 16'b0000000000001010;
        weights2[1787] <= 16'b0000000000010100;
        weights2[1788] <= 16'b0000000000101010;
        weights2[1789] <= 16'b1111111111111010;
        weights2[1790] <= 16'b1111111110111111;
        weights2[1791] <= 16'b1111111111000110;
        weights2[1792] <= 16'b0000000000110101;
        weights2[1793] <= 16'b1111111111101110;
        weights2[1794] <= 16'b1111111111100111;
        weights2[1795] <= 16'b1111111111111011;
        weights2[1796] <= 16'b1111111111110010;
        weights2[1797] <= 16'b0000000000100100;
        weights2[1798] <= 16'b0000000000000000;
        weights2[1799] <= 16'b0000000000001101;
        weights2[1800] <= 16'b0000000000110101;
        weights2[1801] <= 16'b1111111111110110;
        weights2[1802] <= 16'b0000000000001000;
        weights2[1803] <= 16'b0000000000111111;
        weights2[1804] <= 16'b1111111111111011;
        weights2[1805] <= 16'b1111111111110000;
        weights2[1806] <= 16'b1111111111100100;
        weights2[1807] <= 16'b0000000000000101;
        weights2[1808] <= 16'b0000000000110000;
        weights2[1809] <= 16'b0000000001000001;
        weights2[1810] <= 16'b0000000001100111;
        weights2[1811] <= 16'b0000000010010101;
        weights2[1812] <= 16'b1111111110011100;
        weights2[1813] <= 16'b0000000000110111;
        weights2[1814] <= 16'b0000000010010010;
        weights2[1815] <= 16'b0000000001001010;
        weights2[1816] <= 16'b1111111111000111;
        weights2[1817] <= 16'b1111111101010010;
        weights2[1818] <= 16'b0000000000000001;
        weights2[1819] <= 16'b0000000000010001;
        weights2[1820] <= 16'b1111111111000101;
        weights2[1821] <= 16'b1111111101001110;
        weights2[1822] <= 16'b0000000001110101;
        weights2[1823] <= 16'b1111111111100001;
        weights2[1824] <= 16'b0000000000010000;
        weights2[1825] <= 16'b0000000000011101;
        weights2[1826] <= 16'b0000000000000101;
        weights2[1827] <= 16'b0000000000000000;
        weights2[1828] <= 16'b0000000000100111;
        weights2[1829] <= 16'b1111111111011100;
        weights2[1830] <= 16'b1111111111111101;
        weights2[1831] <= 16'b1111111110011110;
        weights2[1832] <= 16'b0000000000001011;
        weights2[1833] <= 16'b0000000000001111;
        weights2[1834] <= 16'b1111111111000011;
        weights2[1835] <= 16'b1111111111010111;
        weights2[1836] <= 16'b0000000000010000;
        weights2[1837] <= 16'b1111111111100010;
        weights2[1838] <= 16'b1111111110111001;
        weights2[1839] <= 16'b0000000000000010;
        weights2[1840] <= 16'b0000000000010000;
        weights2[1841] <= 16'b1111111110111110;
        weights2[1842] <= 16'b1111111101100000;
        weights2[1843] <= 16'b1111111111001101;
        weights2[1844] <= 16'b0000000000000101;
        weights2[1845] <= 16'b1111111111100010;
        weights2[1846] <= 16'b0000000000000000;
        weights2[1847] <= 16'b1111111111101001;
        weights2[1848] <= 16'b1111111111111100;
        weights2[1849] <= 16'b1111111110101000;
        weights2[1850] <= 16'b1111111111111100;
        weights2[1851] <= 16'b1111111101000010;
        weights2[1852] <= 16'b0000000000000111;
        weights2[1853] <= 16'b1111111110101011;
        weights2[1854] <= 16'b0000000000000100;
        weights2[1855] <= 16'b1111111110101011;
        weights2[1856] <= 16'b0000000001011111;
        weights2[1857] <= 16'b0000000000011101;
        weights2[1858] <= 16'b0000000001011000;
        weights2[1859] <= 16'b0000000000011011;
        weights2[1860] <= 16'b1111111111111111;
        weights2[1861] <= 16'b0000000001101101;
        weights2[1862] <= 16'b0000000000000000;
        weights2[1863] <= 16'b1111111111110101;
        weights2[1864] <= 16'b0000000000100011;
        weights2[1865] <= 16'b1111111111111011;
        weights2[1866] <= 16'b1111111111110010;
        weights2[1867] <= 16'b0000000000111010;
        weights2[1868] <= 16'b0000000000011010;
        weights2[1869] <= 16'b0000000000000100;
        weights2[1870] <= 16'b0000000000110110;
        weights2[1871] <= 16'b0000000000000000;
        weights2[1872] <= 16'b0000000000111000;
        weights2[1873] <= 16'b0000000010001110;
        weights2[1874] <= 16'b0000000000111110;
        weights2[1875] <= 16'b0000000001110011;
        weights2[1876] <= 16'b0000000000100100;
        weights2[1877] <= 16'b0000000010100100;
        weights2[1878] <= 16'b0000000001101010;
        weights2[1879] <= 16'b0000000000100100;
        weights2[1880] <= 16'b1111111111110100;
        weights2[1881] <= 16'b1111111110101101;
        weights2[1882] <= 16'b0000000000011010;
        weights2[1883] <= 16'b0000000001011000;
        weights2[1884] <= 16'b1111111111101001;
        weights2[1885] <= 16'b1111111110010000;
        weights2[1886] <= 16'b0000000010110100;
        weights2[1887] <= 16'b0000000000110011;
        weights2[1888] <= 16'b0000000000110010;
        weights2[1889] <= 16'b0000000000100110;
        weights2[1890] <= 16'b0000000000100010;
        weights2[1891] <= 16'b0000000000101010;
        weights2[1892] <= 16'b1111111111010011;
        weights2[1893] <= 16'b0000000000101100;
        weights2[1894] <= 16'b0000000000101110;
        weights2[1895] <= 16'b1111111111100100;
        weights2[1896] <= 16'b1111111111011011;
        weights2[1897] <= 16'b1111111111101111;
        weights2[1898] <= 16'b1111111111111000;
        weights2[1899] <= 16'b1111111111010110;
        weights2[1900] <= 16'b0000000000110111;
        weights2[1901] <= 16'b1111111101110100;
        weights2[1902] <= 16'b1111111111011011;
        weights2[1903] <= 16'b0000000000101101;
        weights2[1904] <= 16'b0000000000001010;
        weights2[1905] <= 16'b0000000000101001;
        weights2[1906] <= 16'b1111111110101111;
        weights2[1907] <= 16'b1111111111000000;
        weights2[1908] <= 16'b0000000000110000;
        weights2[1909] <= 16'b1111111111111111;
        weights2[1910] <= 16'b0000000000000000;
        weights2[1911] <= 16'b0000000000000010;
        weights2[1912] <= 16'b0000000000011010;
        weights2[1913] <= 16'b1111111111010001;
        weights2[1914] <= 16'b1111111111100011;
        weights2[1915] <= 16'b1111111110101111;
        weights2[1916] <= 16'b0000000000011101;
        weights2[1917] <= 16'b1111111111011000;
        weights2[1918] <= 16'b0000000000001010;
        weights2[1919] <= 16'b0000000000000001;
        weights2[1920] <= 16'b1111111111111001;
        weights2[1921] <= 16'b0000000010111100;
        weights2[1922] <= 16'b0000000001011010;
        weights2[1923] <= 16'b0000000000001101;
        weights2[1924] <= 16'b1111111111100011;
        weights2[1925] <= 16'b0000000000011111;
        weights2[1926] <= 16'b0000000000000000;
        weights2[1927] <= 16'b0000000001110001;
        weights2[1928] <= 16'b0000000000111010;
        weights2[1929] <= 16'b1111111111101101;
        weights2[1930] <= 16'b0000000000111011;
        weights2[1931] <= 16'b0000000000010100;
        weights2[1932] <= 16'b0000000010101101;
        weights2[1933] <= 16'b0000000010001001;
        weights2[1934] <= 16'b1111111111111010;
        weights2[1935] <= 16'b1111111111111010;
        weights2[1936] <= 16'b1111111111010001;
        weights2[1937] <= 16'b0000000001001110;
        weights2[1938] <= 16'b1111111111110110;
        weights2[1939] <= 16'b1111111111100011;
        weights2[1940] <= 16'b1111111110001100;
        weights2[1941] <= 16'b0000000001010011;
        weights2[1942] <= 16'b0000000000000001;
        weights2[1943] <= 16'b0000000000000111;
        weights2[1944] <= 16'b0000000000010110;
        weights2[1945] <= 16'b0000000000001011;
        weights2[1946] <= 16'b1111111111111110;
        weights2[1947] <= 16'b0000000000110101;
        weights2[1948] <= 16'b0000000010001001;
        weights2[1949] <= 16'b0000000001001000;
        weights2[1950] <= 16'b0000000001000010;
        weights2[1951] <= 16'b1111111111011110;
        weights2[1952] <= 16'b1111111111010111;
        weights2[1953] <= 16'b1111111111111001;
        weights2[1954] <= 16'b0000000000000010;
        weights2[1955] <= 16'b0000000001000001;
        weights2[1956] <= 16'b0000000001100101;
        weights2[1957] <= 16'b1111111111101101;
        weights2[1958] <= 16'b0000000000011101;
        weights2[1959] <= 16'b1111111111010010;
        weights2[1960] <= 16'b1111111111001001;
        weights2[1961] <= 16'b1111111111101000;
        weights2[1962] <= 16'b0000000000000101;
        weights2[1963] <= 16'b0000000000011001;
        weights2[1964] <= 16'b1111111111101010;
        weights2[1965] <= 16'b0000000000011111;
        weights2[1966] <= 16'b0000000010010010;
        weights2[1967] <= 16'b0000000001010010;
        weights2[1968] <= 16'b0000000000100101;
        weights2[1969] <= 16'b0000000000101011;
        weights2[1970] <= 16'b0000000010011110;
        weights2[1971] <= 16'b1111111111011000;
        weights2[1972] <= 16'b1111111111100100;
        weights2[1973] <= 16'b1111111111001101;
        weights2[1974] <= 16'b0000000000000000;
        weights2[1975] <= 16'b1111111111110000;
        weights2[1976] <= 16'b1111111111111100;
        weights2[1977] <= 16'b0000000000011110;
        weights2[1978] <= 16'b1111111111110001;
        weights2[1979] <= 16'b1111111111100111;
        weights2[1980] <= 16'b1111111111101110;
        weights2[1981] <= 16'b0000000000011010;
        weights2[1982] <= 16'b0000000001010100;
        weights2[1983] <= 16'b0000000000000101;
        weights2[1984] <= 16'b0000000000001001;
        weights2[1985] <= 16'b1111111101101111;
        weights2[1986] <= 16'b0000000000100110;
        weights2[1987] <= 16'b0000000000010011;
        weights2[1988] <= 16'b1111111110111101;
        weights2[1989] <= 16'b0000000000101110;
        weights2[1990] <= 16'b0000000000000000;
        weights2[1991] <= 16'b1111111111100110;
        weights2[1992] <= 16'b0000000000100111;
        weights2[1993] <= 16'b1111111110110100;
        weights2[1994] <= 16'b0000000000000110;
        weights2[1995] <= 16'b1111111101001001;
        weights2[1996] <= 16'b1111111111111111;
        weights2[1997] <= 16'b1111111110100000;
        weights2[1998] <= 16'b0000000000011111;
        weights2[1999] <= 16'b1111111111111001;
        weights2[2000] <= 16'b1111111110011111;
        weights2[2001] <= 16'b0000000000100001;
        weights2[2002] <= 16'b1111111110000101;
        weights2[2003] <= 16'b1111111111000100;
        weights2[2004] <= 16'b1111111111011100;
        weights2[2005] <= 16'b0000000000111101;
        weights2[2006] <= 16'b1111111110101100;
        weights2[2007] <= 16'b0000000000011001;
        weights2[2008] <= 16'b0000000000100100;
        weights2[2009] <= 16'b0000000000110101;
        weights2[2010] <= 16'b1111111110100101;
        weights2[2011] <= 16'b1111111110011010;
        weights2[2012] <= 16'b0000000000001001;
        weights2[2013] <= 16'b0000000000111001;
        weights2[2014] <= 16'b0000000000111100;
        weights2[2015] <= 16'b0000000000010010;
        weights2[2016] <= 16'b0000000000011111;
        weights2[2017] <= 16'b1111111111000101;
        weights2[2018] <= 16'b0000000000010110;
        weights2[2019] <= 16'b0000000000110101;
        weights2[2020] <= 16'b0000000000000100;
        weights2[2021] <= 16'b0000000000010100;
        weights2[2022] <= 16'b0000000000101101;
        weights2[2023] <= 16'b1111111101101100;
        weights2[2024] <= 16'b1111111101110011;
        weights2[2025] <= 16'b1111111101001110;
        weights2[2026] <= 16'b0000000000001001;
        weights2[2027] <= 16'b0000000000011111;
        weights2[2028] <= 16'b0000000000101110;
        weights2[2029] <= 16'b0000000000111001;
        weights2[2030] <= 16'b1111111111101100;
        weights2[2031] <= 16'b1111111101010111;
        weights2[2032] <= 16'b1111111111101110;
        weights2[2033] <= 16'b0000000000110110;
        weights2[2034] <= 16'b0000000000100100;
        weights2[2035] <= 16'b1111111111010001;
        weights2[2036] <= 16'b1111111111010100;
        weights2[2037] <= 16'b1111111110000111;
        weights2[2038] <= 16'b0000000000000000;
        weights2[2039] <= 16'b1111111110111010;
        weights2[2040] <= 16'b1111111110011101;
        weights2[2041] <= 16'b0000000000100101;
        weights2[2042] <= 16'b0000000000000111;
        weights2[2043] <= 16'b1111111110101100;
        weights2[2044] <= 16'b1111111110001000;
        weights2[2045] <= 16'b0000000000111001;
        weights2[2046] <= 16'b1111111111100111;
        weights2[2047] <= 16'b1111111111010000;
        biases2[0] <= 16'b0000000010000011;
        biases2[1] <= 16'b0000000001110011;
        biases2[2] <= 16'b0000000010001011;
        biases2[3] <= 16'b0000000011010100;
        biases2[4] <= 16'b0000000010101100;
        biases2[5] <= 16'b0000000000111101;
        biases2[6] <= 16'b0000000011111100;
        biases2[7] <= 16'b0000000011110111;
        biases2[8] <= 16'b0000000010110001;
        biases2[9] <= 16'b1111111110001000;
        biases2[10] <= 16'b0000000000100001;
        biases2[11] <= 16'b0000000100101101;
        biases2[12] <= 16'b1111111101101000;
        biases2[13] <= 16'b0000000110110010;
        biases2[14] <= 16'b0000000100000101;
        biases2[15] <= 16'b0000000010011100;
        biases2[16] <= 16'b0000000000010100;
        biases2[17] <= 16'b0000000100100011;
        biases2[18] <= 16'b1111111101111111;
        biases2[19] <= 16'b1111111110010101;
        biases2[20] <= 16'b0000000011101001;
        biases2[21] <= 16'b0000000010101111;
        biases2[22] <= 16'b0000000011010101;
        biases2[23] <= 16'b0000000100011011;
        biases2[24] <= 16'b1111111111010110;
        biases2[25] <= 16'b0000000101010010;
        biases2[26] <= 16'b0000000010000000;
        biases2[27] <= 16'b0000000000000111;
        biases2[28] <= 16'b0000000001011011;
        biases2[29] <= 16'b1111111100101010;
        biases2[30] <= 16'b1111111110011101;
        biases2[31] <= 16'b0000000001110000;
        weights3[0] <= 16'b0000000001111011;
        weights3[1] <= 16'b1111111110001010;
        weights3[2] <= 16'b0000000000111111;
        weights3[3] <= 16'b0000000010110101;
        weights3[4] <= 16'b1111111101101011;
        weights3[5] <= 16'b0000000000110001;
        weights3[6] <= 16'b0000000010011111;
        weights3[7] <= 16'b0000000000000000;
        weights3[8] <= 16'b1111111101101001;
        weights3[9] <= 16'b1111111101101000;
        weights3[10] <= 16'b1111111101111110;
        weights3[11] <= 16'b1111111111101110;
        weights3[12] <= 16'b0000000000010110;
        weights3[13] <= 16'b0000000000100100;
        weights3[14] <= 16'b0000000001100010;
        weights3[15] <= 16'b1111111111011101;
        weights3[16] <= 16'b1111111101001100;
        weights3[17] <= 16'b1111111110100000;
        weights3[18] <= 16'b0000000001001101;
        weights3[19] <= 16'b1111111110101111;
        weights3[20] <= 16'b0000000001000001;
        weights3[21] <= 16'b1111111101101101;
        weights3[22] <= 16'b0000000001000000;
        weights3[23] <= 16'b0000000000011101;
        weights3[24] <= 16'b0000000001000100;
        weights3[25] <= 16'b1111111110010100;
        weights3[26] <= 16'b1111111110100000;
        weights3[27] <= 16'b1111111110101011;
        weights3[28] <= 16'b1111111110101010;
        weights3[29] <= 16'b1111111110101010;
        weights3[30] <= 16'b1111111101111001;
        weights3[31] <= 16'b0000000000011010;
        weights3[32] <= 16'b1111111110000100;
        weights3[33] <= 16'b1111111110000010;
        weights3[34] <= 16'b0000000000100111;
        weights3[35] <= 16'b1111111110100111;
        weights3[36] <= 16'b0000000000110110;
        weights3[37] <= 16'b0000000000000110;
        weights3[38] <= 16'b1111111100000000;
        weights3[39] <= 16'b0000000001110000;
        weights3[40] <= 16'b1111111111100011;
        weights3[41] <= 16'b0000000000000011;
        weights3[42] <= 16'b1111111111011101;
        weights3[43] <= 16'b1111111110101101;
        weights3[44] <= 16'b0000000001001011;
        weights3[45] <= 16'b0000000001101011;
        weights3[46] <= 16'b1111111101101010;
        weights3[47] <= 16'b0000000010000111;
        weights3[48] <= 16'b0000000001001011;
        weights3[49] <= 16'b1111111100100011;
        weights3[50] <= 16'b0000000000000101;
        weights3[51] <= 16'b0000000000110001;
        weights3[52] <= 16'b0000000000011111;
        weights3[53] <= 16'b1111111101011101;
        weights3[54] <= 16'b1111111101111001;
        weights3[55] <= 16'b0000000000010100;
        weights3[56] <= 16'b0000000000110110;
        weights3[57] <= 16'b0000000001010010;
        weights3[58] <= 16'b0000000001000001;
        weights3[59] <= 16'b1111111101101010;
        weights3[60] <= 16'b0000000000001001;
        weights3[61] <= 16'b0000000001001101;
        weights3[62] <= 16'b0000000001011100;
        weights3[63] <= 16'b0000000011000111;
        weights3[64] <= 16'b0000000001001011;
        weights3[65] <= 16'b1111111110001110;
        weights3[66] <= 16'b0000000000101000;
        weights3[67] <= 16'b1111111101101011;
        weights3[68] <= 16'b1111111110011001;
        weights3[69] <= 16'b0000000000011101;
        weights3[70] <= 16'b1111111111011101;
        weights3[71] <= 16'b1111111111010010;
        weights3[72] <= 16'b1111111110101100;
        weights3[73] <= 16'b0000000000110010;
        weights3[74] <= 16'b0000000000110101;
        weights3[75] <= 16'b0000000001111000;
        weights3[76] <= 16'b0000000000001100;
        weights3[77] <= 16'b1111111101011010;
        weights3[78] <= 16'b1111111110111110;
        weights3[79] <= 16'b1111111101111110;
        weights3[80] <= 16'b1111111110100000;
        weights3[81] <= 16'b0000000000010111;
        weights3[82] <= 16'b0000000001000000;
        weights3[83] <= 16'b0000000000111000;
        weights3[84] <= 16'b1111111110001110;
        weights3[85] <= 16'b1111111110110010;
        weights3[86] <= 16'b1111111111111100;
        weights3[87] <= 16'b0000000000000001;
        weights3[88] <= 16'b0000000000110110;
        weights3[89] <= 16'b1111111101011101;
        weights3[90] <= 16'b1111111101100110;
        weights3[91] <= 16'b1111111111111010;
        weights3[92] <= 16'b0000000001001101;
        weights3[93] <= 16'b0000000001010110;
        weights3[94] <= 16'b0000000000000101;
        weights3[95] <= 16'b1111111110011001;
        weights3[96] <= 16'b1111111111000010;
        weights3[97] <= 16'b0000000001000101;
        weights3[98] <= 16'b0000000000110010;
        weights3[99] <= 16'b1111111101111100;
        weights3[100] <= 16'b1111111110110110;
        weights3[101] <= 16'b1111111110101100;
        weights3[102] <= 16'b1111111110111011;
        weights3[103] <= 16'b1111111110111111;
        weights3[104] <= 16'b0000000000110011;
        weights3[105] <= 16'b1111111110111101;
        weights3[106] <= 16'b0000000000110000;
        weights3[107] <= 16'b1111111111011001;
        weights3[108] <= 16'b1111111110110100;
        weights3[109] <= 16'b1111111101101001;
        weights3[110] <= 16'b1111111111011100;
        weights3[111] <= 16'b1111111101100011;
        weights3[112] <= 16'b0000000001000110;
        weights3[113] <= 16'b1111111110101010;
        weights3[114] <= 16'b0000000000111111;
        weights3[115] <= 16'b0000000000010011;
        weights3[116] <= 16'b1111111101101111;
        weights3[117] <= 16'b1111111110011111;
        weights3[118] <= 16'b0000000000110110;
        weights3[119] <= 16'b0000000001000100;
        weights3[120] <= 16'b1111111111001011;
        weights3[121] <= 16'b1111111110101001;
        weights3[122] <= 16'b0000000000111001;
        weights3[123] <= 16'b0000000000110011;
        weights3[124] <= 16'b0000000001001011;
        weights3[125] <= 16'b0000000001000011;
        weights3[126] <= 16'b0000000000100111;
        weights3[127] <= 16'b1111111110011101;
        weights3[128] <= 16'b1111111111011101;
        weights3[129] <= 16'b1111111110101010;
        weights3[130] <= 16'b1111111100011000;
        weights3[131] <= 16'b1111111111101100;
        weights3[132] <= 16'b0000000001010011;
        weights3[133] <= 16'b0000000001000001;
        weights3[134] <= 16'b0000000001100101;
        weights3[135] <= 16'b1111111110010100;
        weights3[136] <= 16'b1111111110000100;
        weights3[137] <= 16'b0000000000011110;
        weights3[138] <= 16'b1111111110100101;
        weights3[139] <= 16'b1111111111010110;
        weights3[140] <= 16'b0000000001000001;
        weights3[141] <= 16'b0000000000111000;
        weights3[142] <= 16'b1111111101111000;
        weights3[143] <= 16'b1111111111111101;
        weights3[144] <= 16'b0000000000011001;
        weights3[145] <= 16'b0000000001101110;
        weights3[146] <= 16'b1111111101110110;
        weights3[147] <= 16'b0000000000111010;
        weights3[148] <= 16'b1111111111010010;
        weights3[149] <= 16'b0000000001000001;
        weights3[150] <= 16'b1111111110001111;
        weights3[151] <= 16'b1111111110001011;
        weights3[152] <= 16'b0000000000111001;
        weights3[153] <= 16'b0000000001011011;
        weights3[154] <= 16'b0000000001001110;
        weights3[155] <= 16'b0000000000111000;
        weights3[156] <= 16'b1111111110000110;
        weights3[157] <= 16'b1111111110100111;
        weights3[158] <= 16'b1111111101011111;
        weights3[159] <= 16'b1111111101011101;
        weights3[160] <= 16'b1111111110111101;
        weights3[161] <= 16'b0000000001001010;
        weights3[162] <= 16'b1111111111111110;
        weights3[163] <= 16'b1111111110000100;
        weights3[164] <= 16'b1111111110100011;
        weights3[165] <= 16'b1111111110111010;
        weights3[166] <= 16'b1111111110110010;
        weights3[167] <= 16'b1111111111010110;
        weights3[168] <= 16'b0000000001010100;
        weights3[169] <= 16'b1111111111110111;
        weights3[170] <= 16'b0000000000101111;
        weights3[171] <= 16'b1111111110110110;
        weights3[172] <= 16'b0000000001000101;
        weights3[173] <= 16'b1111111101110110;
        weights3[174] <= 16'b0000000000111111;
        weights3[175] <= 16'b1111111111000110;
        weights3[176] <= 16'b0000000000111111;
        weights3[177] <= 16'b1111111110101111;
        weights3[178] <= 16'b0000000000101011;
        weights3[179] <= 16'b1111111111100001;
        weights3[180] <= 16'b0000000001010010;
        weights3[181] <= 16'b0000000001001001;
        weights3[182] <= 16'b0000000000110001;
        weights3[183] <= 16'b1111111101000100;
        weights3[184] <= 16'b1111111110101101;
        weights3[185] <= 16'b1111111110100000;
        weights3[186] <= 16'b1111111111001011;
        weights3[187] <= 16'b0000000000101111;
        weights3[188] <= 16'b1111111110101010;
        weights3[189] <= 16'b1111111110011000;
        weights3[190] <= 16'b0000000000110100;
        weights3[191] <= 16'b1111111110110111;
        weights3[192] <= 16'b0000000001011101;
        weights3[193] <= 16'b1111111111110000;
        weights3[194] <= 16'b1111111110011011;
        weights3[195] <= 16'b0000000001110011;
        weights3[196] <= 16'b1111111110001110;
        weights3[197] <= 16'b1111111100110001;
        weights3[198] <= 16'b0000000010000001;
        weights3[199] <= 16'b1111111110001011;
        weights3[200] <= 16'b0000000001001001;
        weights3[201] <= 16'b0000000000101100;
        weights3[202] <= 16'b1111111100100100;
        weights3[203] <= 16'b0000000001001001;
        weights3[204] <= 16'b0000000001000001;
        weights3[205] <= 16'b1111111111011100;
        weights3[206] <= 16'b1111111110111110;
        weights3[207] <= 16'b0000000010101000;
        weights3[208] <= 16'b1111111101111100;
        weights3[209] <= 16'b0000000000111101;
        weights3[210] <= 16'b1111111101001111;
        weights3[211] <= 16'b0000000000101110;
        weights3[212] <= 16'b0000000001100010;
        weights3[213] <= 16'b0000000001011111;
        weights3[214] <= 16'b0000000000101001;
        weights3[215] <= 16'b1111111100011010;
        weights3[216] <= 16'b0000000000110000;
        weights3[217] <= 16'b1111111110000110;
        weights3[218] <= 16'b1111111111101001;
        weights3[219] <= 16'b1111111101010101;
        weights3[220] <= 16'b1111111110001001;
        weights3[221] <= 16'b1111111111001101;
        weights3[222] <= 16'b0000000000101111;
        weights3[223] <= 16'b0000000000010001;
        weights3[224] <= 16'b1111111101110011;
        weights3[225] <= 16'b1111111101100001;
        weights3[226] <= 16'b0000000000110011;
        weights3[227] <= 16'b1111111110101111;
        weights3[228] <= 16'b0000000001100100;
        weights3[229] <= 16'b0000000001001111;
        weights3[230] <= 16'b1111111110000001;
        weights3[231] <= 16'b0000000010000010;
        weights3[232] <= 16'b1111111101111111;
        weights3[233] <= 16'b0000000000101100;
        weights3[234] <= 16'b0000000000101111;
        weights3[235] <= 16'b1111111111011100;
        weights3[236] <= 16'b0000000001000000;
        weights3[237] <= 16'b1111111110101011;
        weights3[238] <= 16'b0000000001010000;
        weights3[239] <= 16'b1111111100111100;
        weights3[240] <= 16'b0000000001010101;
        weights3[241] <= 16'b1111111111010111;
        weights3[242] <= 16'b0000000000111000;
        weights3[243] <= 16'b1111111110101111;
        weights3[244] <= 16'b1111111110001100;
        weights3[245] <= 16'b1111111111010000;
        weights3[246] <= 16'b1111111100111111;
        weights3[247] <= 16'b0000000001000110;
        weights3[248] <= 16'b1111111110101000;
        weights3[249] <= 16'b1111111111001000;
        weights3[250] <= 16'b1111111110001110;
        weights3[251] <= 16'b0000000001000010;
        weights3[252] <= 16'b0000000000110010;
        weights3[253] <= 16'b0000000001001111;
        weights3[254] <= 16'b1111111110001111;
        weights3[255] <= 16'b1111111110111111;
        weights3[256] <= 16'b1111111111101110;
        weights3[257] <= 16'b0000000000100110;
        weights3[258] <= 16'b0000000000101110;
        weights3[259] <= 16'b1111111101100001;
        weights3[260] <= 16'b1111111110011111;
        weights3[261] <= 16'b1111111110100000;
        weights3[262] <= 16'b1111111101111011;
        weights3[263] <= 16'b0000000010010011;
        weights3[264] <= 16'b0000000001000011;
        weights3[265] <= 16'b1111111110101001;
        weights3[266] <= 16'b1111111111111100;
        weights3[267] <= 16'b0000000001101101;
        weights3[268] <= 16'b1111111111010001;
        weights3[269] <= 16'b0000000001100000;
        weights3[270] <= 16'b0000000000111011;
        weights3[271] <= 16'b1111111111001011;
        weights3[272] <= 16'b1111111110111110;
        weights3[273] <= 16'b1111111101110000;
        weights3[274] <= 16'b1111111111000101;
        weights3[275] <= 16'b1111111111100011;
        weights3[276] <= 16'b0000000000111010;
        weights3[277] <= 16'b0000000000011101;
        weights3[278] <= 16'b0000000000010110;
        weights3[279] <= 16'b0000000000100110;
        weights3[280] <= 16'b1111111111001010;
        weights3[281] <= 16'b0000000001101000;
        weights3[282] <= 16'b0000000000010010;
        weights3[283] <= 16'b1111111111001110;
        weights3[284] <= 16'b0000000000110011;
        weights3[285] <= 16'b1111111111001011;
        weights3[286] <= 16'b1111111111001111;
        weights3[287] <= 16'b0000000000010110;
        weights3[288] <= 16'b1111111111101101;
        weights3[289] <= 16'b0000000000111111;
        weights3[290] <= 16'b1111111110010010;
        weights3[291] <= 16'b0000000000001110;
        weights3[292] <= 16'b0000000001010011;
        weights3[293] <= 16'b0000000001000001;
        weights3[294] <= 16'b0000000001101111;
        weights3[295] <= 16'b1111111111001111;
        weights3[296] <= 16'b1111111111001010;
        weights3[297] <= 16'b1111111111001000;
        weights3[298] <= 16'b0000000000100000;
        weights3[299] <= 16'b1111111111000110;
        weights3[300] <= 16'b1111111101110110;
        weights3[301] <= 16'b0000000000010011;
        weights3[302] <= 16'b0000000001001001;
        weights3[303] <= 16'b1111111110001010;
        weights3[304] <= 16'b0000000000111101;
        weights3[305] <= 16'b0000000001110010;
        weights3[306] <= 16'b0000000000000110;
        weights3[307] <= 16'b1111111101100110;
        weights3[308] <= 16'b1111111110111001;
        weights3[309] <= 16'b0000000000001010;
        weights3[310] <= 16'b1111111110000010;
        weights3[311] <= 16'b0000000001100010;
        weights3[312] <= 16'b1111111101110010;
        weights3[313] <= 16'b0000000001000110;
        weights3[314] <= 16'b0000000000011011;
        weights3[315] <= 16'b0000000000101011;
        weights3[316] <= 16'b1111111101011110;
        weights3[317] <= 16'b1111111111011111;
        weights3[318] <= 16'b1111111111011101;
        weights3[319] <= 16'b1111111101111110;
        biases3[0] <= 16'b0000000000000100;
        biases3[1] <= 16'b1111111011110110;
        biases3[2] <= 16'b0000000000011001;
        biases3[3] <= 16'b1111111111110100;
        biases3[4] <= 16'b0000000001000000;
        biases3[5] <= 16'b0000000000110111;
        biases3[6] <= 16'b1111111110001101;
        biases3[7] <= 16'b1111111101100110;
        biases3[8] <= 16'b0000000011001010;
        biases3[9] <= 16'b0000000010001111;
    end

endmodule
