module neural_tb ();
    reg clk;
    reg rst;
    reg start;
    reg [783:0] in_features;
    wire [3:0] prediction;
    wire done;

    // instantiate the unit under test
    NeuralNetwork dut (
        .clk(clk),
        .rst(rst),
        .start(start),
        .in_features(in_features),
        .prediction(prediction),
        .done(done)
    );

    // clock generation
    always begin
        #5 clk = 0;
        #5 clk = 1;
    end

    // reset generation
    initial begin
        rst = 1;
        start = 0;
        in_features = 0;
        #10 rst = 0;
        in_features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000011111100000000000000000000011000000000000000000000000001000000000000000000000000001100000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000000000000000000101111111000000000000000000010100000111000000000000000001110000000110000000000000000110000000001000000000000000011000000000100000000000000000100000000010000000000000000010000000001000000000000000000110000001000000000000000000001111111000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        #10 start = 1;
        #10 start = 0;
        #50;
        in_features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000110011000000000000000000000110000110000000000000000000010000001100000000000000000011000000110000000000000000001100000010000000000000000000010000001000000000000000000001100001100000000000000000000010000100000000000000000000000100100000000000000000000000001100000000000000000000000001001100000000000000000000001000001000000000000000000001000000010000000000000000000100000001000000000000000000100000000110000000000000000010000000011000000000000000001000000011000000000000000000111111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        #10 start = 1;
        #10 start = 0;
    end
endmodule